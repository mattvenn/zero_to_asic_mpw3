magic
tech sky130A
magscale 1 2
timestamp 1635348390
<< metal1 >>
rect 191742 703400 191748 703452
rect 191800 703440 191806 703452
rect 283834 703440 283840 703452
rect 191800 703412 283840 703440
rect 191800 703400 191806 703412
rect 283834 703400 283840 703412
rect 283892 703400 283898 703452
rect 282822 703332 282828 703384
rect 282880 703372 282886 703384
rect 348786 703372 348792 703384
rect 282880 703344 348792 703372
rect 282880 703332 282886 703344
rect 348786 703332 348792 703344
rect 348844 703332 348850 703384
rect 214558 703264 214564 703316
rect 214616 703304 214622 703316
rect 364978 703304 364984 703316
rect 214616 703276 364984 703304
rect 214616 703264 214622 703276
rect 364978 703264 364984 703276
rect 365036 703264 365042 703316
rect 240778 703196 240784 703248
rect 240836 703236 240842 703248
rect 332502 703236 332508 703248
rect 240836 703208 332508 703236
rect 240836 703196 240842 703208
rect 332502 703196 332508 703208
rect 332560 703196 332566 703248
rect 249058 703128 249064 703180
rect 249116 703168 249122 703180
rect 413646 703168 413652 703180
rect 249116 703140 413652 703168
rect 249116 703128 249122 703140
rect 413646 703128 413652 703140
rect 413704 703128 413710 703180
rect 273898 703060 273904 703112
rect 273956 703100 273962 703112
rect 462314 703100 462320 703112
rect 273956 703072 462320 703100
rect 273956 703060 273962 703072
rect 462314 703060 462320 703072
rect 462372 703060 462378 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 102042 702992 102048 703044
rect 102100 703032 102106 703044
rect 300118 703032 300124 703044
rect 102100 703004 300124 703032
rect 102100 702992 102106 703004
rect 300118 702992 300124 703004
rect 300176 702992 300182 703044
rect 271138 702924 271144 702976
rect 271196 702964 271202 702976
rect 478506 702964 478512 702976
rect 271196 702936 478512 702964
rect 271196 702924 271202 702936
rect 478506 702924 478512 702936
rect 478564 702924 478570 702976
rect 8110 702856 8116 702908
rect 8168 702896 8174 702908
rect 96614 702896 96620 702908
rect 8168 702868 96620 702896
rect 8168 702856 8174 702868
rect 96614 702856 96620 702868
rect 96672 702856 96678 702908
rect 213178 702856 213184 702908
rect 213236 702896 213242 702908
rect 429838 702896 429844 702908
rect 213236 702868 429844 702896
rect 213236 702856 213242 702868
rect 429838 702856 429844 702868
rect 429896 702856 429902 702908
rect 24302 702788 24308 702840
rect 24360 702828 24366 702840
rect 86218 702828 86224 702840
rect 24360 702800 86224 702828
rect 24360 702788 24366 702800
rect 86218 702788 86224 702800
rect 86276 702788 86282 702840
rect 177298 702788 177304 702840
rect 177356 702828 177362 702840
rect 397454 702828 397460 702840
rect 177356 702800 397460 702828
rect 177356 702788 177362 702800
rect 397454 702788 397460 702800
rect 397512 702788 397518 702840
rect 69658 702720 69664 702772
rect 69716 702760 69722 702772
rect 154114 702760 154120 702772
rect 69716 702732 154120 702760
rect 69716 702720 69722 702732
rect 154114 702720 154120 702732
rect 154172 702720 154178 702772
rect 280798 702720 280804 702772
rect 280856 702760 280862 702772
rect 543458 702760 543464 702772
rect 280856 702732 543464 702760
rect 280856 702720 280862 702732
rect 543458 702720 543464 702732
rect 543516 702720 543522 702772
rect 90358 702652 90364 702704
rect 90416 702692 90422 702704
rect 235166 702692 235172 702704
rect 90416 702664 235172 702692
rect 90416 702652 90422 702664
rect 235166 702652 235172 702664
rect 235224 702652 235230 702704
rect 258718 702652 258724 702704
rect 258776 702692 258782 702704
rect 559650 702692 559656 702704
rect 258776 702664 559656 702692
rect 258776 702652 258782 702664
rect 559650 702652 559656 702664
rect 559708 702652 559714 702704
rect 84102 702584 84108 702636
rect 84160 702624 84166 702636
rect 202782 702624 202788 702636
rect 84160 702596 202788 702624
rect 84160 702584 84166 702596
rect 202782 702584 202788 702596
rect 202840 702584 202846 702636
rect 215938 702584 215944 702636
rect 215996 702624 216002 702636
rect 527082 702624 527088 702636
rect 215996 702596 527088 702624
rect 215996 702584 216002 702596
rect 527082 702584 527088 702596
rect 527140 702584 527146 702636
rect 67634 702516 67640 702568
rect 67692 702556 67698 702568
rect 170306 702556 170312 702568
rect 67692 702528 170312 702556
rect 67692 702516 67698 702528
rect 170306 702516 170312 702528
rect 170364 702516 170370 702568
rect 184842 702516 184848 702568
rect 184900 702556 184906 702568
rect 580902 702556 580908 702568
rect 184900 702528 580908 702556
rect 184900 702516 184906 702528
rect 580902 702516 580908 702528
rect 580960 702516 580966 702568
rect 79962 702448 79968 702500
rect 80020 702488 80026 702500
rect 494790 702488 494796 702500
rect 80020 702460 494796 702488
rect 80020 702448 80026 702460
rect 494790 702448 494796 702460
rect 494848 702448 494854 702500
rect 71682 700272 71688 700324
rect 71740 700312 71746 700324
rect 105446 700312 105452 700324
rect 71740 700284 105452 700312
rect 71740 700272 71746 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 220078 700272 220084 700324
rect 220136 700312 220142 700324
rect 267642 700312 267648 700324
rect 220136 700284 267648 700312
rect 220136 700272 220142 700284
rect 267642 700272 267648 700284
rect 267700 700272 267706 700324
rect 218974 698912 218980 698964
rect 219032 698952 219038 698964
rect 241514 698952 241520 698964
rect 219032 698924 241520 698952
rect 219032 698912 219038 698924
rect 241514 698912 241520 698924
rect 241572 698912 241578 698964
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 11698 683176 11704 683188
rect 3476 683148 11704 683176
rect 3476 683136 3482 683148
rect 11698 683136 11704 683148
rect 11756 683136 11762 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 14458 670732 14464 670744
rect 3568 670704 14464 670732
rect 3568 670692 3574 670704
rect 14458 670692 14464 670704
rect 14516 670692 14522 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 74534 656928 74540 656940
rect 3476 656900 74540 656928
rect 3476 656888 3482 656900
rect 74534 656888 74540 656900
rect 74592 656888 74598 656940
rect 3510 618604 3516 618656
rect 3568 618644 3574 618656
rect 7558 618644 7564 618656
rect 3568 618616 7564 618644
rect 3568 618604 3574 618616
rect 7558 618604 7564 618616
rect 7616 618604 7622 618656
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 93118 605860 93124 605872
rect 3568 605832 93124 605860
rect 3568 605820 3574 605832
rect 93118 605820 93124 605832
rect 93176 605820 93182 605872
rect 81434 592628 81440 592680
rect 81492 592668 81498 592680
rect 84102 592668 84108 592680
rect 81492 592640 84108 592668
rect 81492 592628 81498 592640
rect 84102 592628 84108 592640
rect 84160 592668 84166 592680
rect 143534 592668 143540 592680
rect 84160 592640 143540 592668
rect 84160 592628 84166 592640
rect 143534 592628 143540 592640
rect 143592 592628 143598 592680
rect 79318 589840 79324 589892
rect 79376 589880 79382 589892
rect 79962 589880 79968 589892
rect 79376 589852 79968 589880
rect 79376 589840 79382 589852
rect 79962 589840 79968 589852
rect 80020 589840 80026 589892
rect 79962 589296 79968 589348
rect 80020 589336 80026 589348
rect 124214 589336 124220 589348
rect 80020 589308 124220 589336
rect 80020 589296 80026 589308
rect 124214 589296 124220 589308
rect 124272 589296 124278 589348
rect 67542 588548 67548 588600
rect 67600 588588 67606 588600
rect 71682 588588 71688 588600
rect 67600 588560 71688 588588
rect 67600 588548 67606 588560
rect 71682 588548 71688 588560
rect 71740 588588 71746 588600
rect 128354 588588 128360 588600
rect 71740 588560 128360 588588
rect 71740 588548 71746 588560
rect 128354 588548 128360 588560
rect 128412 588548 128418 588600
rect 40034 587120 40040 587172
rect 40092 587160 40098 587172
rect 96706 587160 96712 587172
rect 40092 587132 96712 587160
rect 40092 587120 40098 587132
rect 96706 587120 96712 587132
rect 96764 587120 96770 587172
rect 82722 586508 82728 586560
rect 82780 586548 82786 586560
rect 123478 586548 123484 586560
rect 82780 586520 123484 586548
rect 82780 586508 82786 586520
rect 123478 586508 123484 586520
rect 123536 586508 123542 586560
rect 78122 585760 78128 585812
rect 78180 585800 78186 585812
rect 88334 585800 88340 585812
rect 78180 585772 88340 585800
rect 78180 585760 78186 585772
rect 88334 585760 88340 585772
rect 88392 585800 88398 585812
rect 112438 585800 112444 585812
rect 88392 585772 112444 585800
rect 88392 585760 88398 585772
rect 112438 585760 112444 585772
rect 112496 585760 112502 585812
rect 121730 585760 121736 585812
rect 121788 585800 121794 585812
rect 582742 585800 582748 585812
rect 121788 585772 582748 585800
rect 121788 585760 121794 585772
rect 582742 585760 582748 585772
rect 582800 585760 582806 585812
rect 52362 585148 52368 585200
rect 52420 585188 52426 585200
rect 84286 585188 84292 585200
rect 52420 585160 84292 585188
rect 52420 585148 52426 585160
rect 84286 585148 84292 585160
rect 84344 585148 84350 585200
rect 87506 585148 87512 585200
rect 87564 585188 87570 585200
rect 121454 585188 121460 585200
rect 87564 585160 121460 585188
rect 87564 585148 87570 585160
rect 121454 585148 121460 585160
rect 121512 585188 121518 585200
rect 121730 585188 121736 585200
rect 121512 585160 121736 585188
rect 121512 585148 121518 585160
rect 121730 585148 121736 585160
rect 121788 585148 121794 585200
rect 93118 584400 93124 584452
rect 93176 584440 93182 584452
rect 97258 584440 97264 584452
rect 93176 584412 97264 584440
rect 93176 584400 93182 584412
rect 97258 584400 97264 584412
rect 97316 584400 97322 584452
rect 76282 583720 76288 583772
rect 76340 583760 76346 583772
rect 108298 583760 108304 583772
rect 76340 583732 108304 583760
rect 76340 583720 76346 583732
rect 108298 583720 108304 583732
rect 108356 583720 108362 583772
rect 77202 582768 77208 582820
rect 77260 582808 77266 582820
rect 79318 582808 79324 582820
rect 77260 582780 79324 582808
rect 77260 582768 77266 582780
rect 79318 582768 79324 582780
rect 79376 582768 79382 582820
rect 86218 582496 86224 582548
rect 86276 582536 86282 582548
rect 106918 582536 106924 582548
rect 86276 582508 106924 582536
rect 86276 582496 86282 582508
rect 106918 582496 106924 582508
rect 106976 582496 106982 582548
rect 79042 582428 79048 582480
rect 79100 582468 79106 582480
rect 86862 582468 86868 582480
rect 79100 582440 86868 582468
rect 79100 582428 79106 582440
rect 86862 582428 86868 582440
rect 86920 582428 86926 582480
rect 50982 582360 50988 582412
rect 51040 582400 51046 582412
rect 69934 582400 69940 582412
rect 51040 582372 69940 582400
rect 51040 582360 51046 582372
rect 69934 582360 69940 582372
rect 69992 582360 69998 582412
rect 73522 582360 73528 582412
rect 73580 582400 73586 582412
rect 95878 582400 95884 582412
rect 73580 582372 95884 582400
rect 73580 582360 73586 582372
rect 95878 582360 95884 582372
rect 95936 582360 95942 582412
rect 62022 581068 62028 581120
rect 62080 581108 62086 581120
rect 90542 581108 90548 581120
rect 62080 581080 90548 581108
rect 62080 581068 62086 581080
rect 90542 581068 90548 581080
rect 90600 581068 90606 581120
rect 60642 581000 60648 581052
rect 60700 581040 60706 581052
rect 69014 581040 69020 581052
rect 60700 581012 69020 581040
rect 60700 581000 60706 581012
rect 69014 581000 69020 581012
rect 69072 581000 69078 581052
rect 80238 581040 80244 581052
rect 69676 581012 80244 581040
rect 3142 580932 3148 580984
rect 3200 580972 3206 580984
rect 69676 580972 69704 581012
rect 80238 581000 80244 581012
rect 80296 581000 80302 581052
rect 90266 581000 90272 581052
rect 90324 581040 90330 581052
rect 104250 581040 104256 581052
rect 90324 581012 104256 581040
rect 90324 581000 90330 581012
rect 104250 581000 104256 581012
rect 104308 581000 104314 581052
rect 3200 580944 69704 580972
rect 3200 580932 3206 580944
rect 86862 580660 86868 580712
rect 86920 580660 86926 580712
rect 93762 580660 93768 580712
rect 93820 580700 93826 580712
rect 93820 580672 103514 580700
rect 93820 580660 93826 580672
rect 86880 580632 86908 580660
rect 86880 580604 93854 580632
rect 93826 580292 93854 580604
rect 102778 580292 102784 580304
rect 93826 580264 102784 580292
rect 102778 580252 102784 580264
rect 102836 580252 102842 580304
rect 103486 579680 103514 580672
rect 141418 579680 141424 579692
rect 103486 579652 141424 579680
rect 141418 579640 141424 579652
rect 141476 579640 141482 579692
rect 97166 578212 97172 578264
rect 97224 578252 97230 578264
rect 134518 578252 134524 578264
rect 97224 578224 134524 578252
rect 97224 578212 97230 578224
rect 134518 578212 134524 578224
rect 134576 578212 134582 578264
rect 97994 576852 98000 576904
rect 98052 576892 98058 576904
rect 132586 576892 132592 576904
rect 98052 576864 132592 576892
rect 98052 576852 98058 576864
rect 132586 576852 132592 576864
rect 132644 576852 132650 576904
rect 3418 576784 3424 576836
rect 3476 576824 3482 576836
rect 67726 576824 67732 576836
rect 3476 576796 67732 576824
rect 3476 576784 3482 576796
rect 67726 576784 67732 576796
rect 67784 576784 67790 576836
rect 97902 576716 97908 576768
rect 97960 576756 97966 576768
rect 102042 576756 102048 576768
rect 97960 576728 102048 576756
rect 97960 576716 97966 576728
rect 102042 576716 102048 576728
rect 102100 576716 102106 576768
rect 102042 576104 102048 576156
rect 102100 576144 102106 576156
rect 125594 576144 125600 576156
rect 102100 576116 125600 576144
rect 102100 576104 102106 576116
rect 125594 576104 125600 576116
rect 125652 576104 125658 576156
rect 94682 573316 94688 573368
rect 94740 573356 94746 573368
rect 126974 573356 126980 573368
rect 94740 573328 126980 573356
rect 94740 573316 94746 573328
rect 126974 573316 126980 573328
rect 127032 573316 127038 573368
rect 96982 572704 96988 572756
rect 97040 572744 97046 572756
rect 100846 572744 100852 572756
rect 97040 572716 100852 572744
rect 97040 572704 97046 572716
rect 100846 572704 100852 572716
rect 100904 572704 100910 572756
rect 53650 571344 53656 571396
rect 53708 571384 53714 571396
rect 66806 571384 66812 571396
rect 53708 571356 66812 571384
rect 53708 571344 53714 571356
rect 66806 571344 66812 571356
rect 66864 571344 66870 571396
rect 97534 571344 97540 571396
rect 97592 571384 97598 571396
rect 99374 571384 99380 571396
rect 97592 571356 99380 571384
rect 97592 571344 97598 571356
rect 99374 571344 99380 571356
rect 99432 571344 99438 571396
rect 97258 570664 97264 570716
rect 97316 570704 97322 570716
rect 98730 570704 98736 570716
rect 97316 570676 98736 570704
rect 97316 570664 97322 570676
rect 98730 570664 98736 570676
rect 98788 570664 98794 570716
rect 55030 570596 55036 570648
rect 55088 570636 55094 570648
rect 66714 570636 66720 570648
rect 55088 570608 66720 570636
rect 55088 570596 55094 570608
rect 66714 570596 66720 570608
rect 66772 570596 66778 570648
rect 59262 569984 59268 570036
rect 59320 570024 59326 570036
rect 66898 570024 66904 570036
rect 59320 569996 66904 570024
rect 59320 569984 59326 569996
rect 66898 569984 66904 569996
rect 66956 569984 66962 570036
rect 97902 569916 97908 569968
rect 97960 569956 97966 569968
rect 109678 569956 109684 569968
rect 97960 569928 109684 569956
rect 97960 569916 97966 569928
rect 109678 569916 109684 569928
rect 109736 569916 109742 569968
rect 64690 568556 64696 568608
rect 64748 568596 64754 568608
rect 66530 568596 66536 568608
rect 64748 568568 66536 568596
rect 64748 568556 64754 568568
rect 66530 568556 66536 568568
rect 66588 568556 66594 568608
rect 95878 567808 95884 567860
rect 95936 567848 95942 567860
rect 111058 567848 111064 567860
rect 95936 567820 111064 567848
rect 95936 567808 95942 567820
rect 111058 567808 111064 567820
rect 111116 567808 111122 567860
rect 57698 565836 57704 565888
rect 57756 565876 57762 565888
rect 67634 565876 67640 565888
rect 57756 565848 67640 565876
rect 57756 565836 57762 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 56502 564408 56508 564460
rect 56560 564448 56566 564460
rect 66898 564448 66904 564460
rect 56560 564420 66904 564448
rect 56560 564408 56566 564420
rect 66898 564408 66904 564420
rect 66956 564408 66962 564460
rect 52270 563048 52276 563100
rect 52328 563088 52334 563100
rect 66898 563088 66904 563100
rect 52328 563060 66904 563088
rect 52328 563048 52334 563060
rect 66898 563048 66904 563060
rect 66956 563048 66962 563100
rect 96798 561688 96804 561740
rect 96856 561728 96862 561740
rect 113174 561728 113180 561740
rect 96856 561700 113180 561728
rect 96856 561688 96862 561700
rect 113174 561688 113180 561700
rect 113232 561688 113238 561740
rect 48130 560260 48136 560312
rect 48188 560300 48194 560312
rect 66806 560300 66812 560312
rect 48188 560272 66812 560300
rect 48188 560260 48194 560272
rect 66806 560260 66812 560272
rect 66864 560260 66870 560312
rect 96798 560260 96804 560312
rect 96856 560300 96862 560312
rect 117314 560300 117320 560312
rect 96856 560272 117320 560300
rect 96856 560260 96862 560272
rect 117314 560260 117320 560272
rect 117372 560260 117378 560312
rect 97074 558968 97080 559020
rect 97132 559008 97138 559020
rect 100018 559008 100024 559020
rect 97132 558980 100024 559008
rect 97132 558968 97138 558980
rect 100018 558968 100024 558980
rect 100076 558968 100082 559020
rect 57882 558900 57888 558952
rect 57940 558940 57946 558952
rect 66806 558940 66812 558952
rect 57940 558912 66812 558940
rect 57940 558900 57946 558912
rect 66806 558900 66812 558912
rect 66864 558900 66870 558952
rect 97902 558152 97908 558204
rect 97960 558192 97966 558204
rect 122834 558192 122840 558204
rect 97960 558164 122840 558192
rect 97960 558152 97966 558164
rect 122834 558152 122840 558164
rect 122892 558152 122898 558204
rect 61930 557540 61936 557592
rect 61988 557580 61994 557592
rect 66806 557580 66812 557592
rect 61988 557552 66812 557580
rect 61988 557540 61994 557552
rect 66806 557540 66812 557552
rect 66864 557540 66870 557592
rect 96614 556928 96620 556980
rect 96672 556968 96678 556980
rect 97074 556968 97080 556980
rect 96672 556940 97080 556968
rect 96672 556928 96678 556940
rect 97074 556928 97080 556940
rect 97132 556928 97138 556980
rect 96706 554752 96712 554804
rect 96764 554792 96770 554804
rect 128998 554792 129004 554804
rect 96764 554764 129004 554792
rect 96764 554752 96770 554764
rect 128998 554752 129004 554764
rect 129056 554752 129062 554804
rect 2774 553800 2780 553852
rect 2832 553840 2838 553852
rect 4798 553840 4804 553852
rect 2832 553812 4804 553840
rect 2832 553800 2838 553812
rect 4798 553800 4804 553812
rect 4856 553800 4862 553852
rect 63310 553392 63316 553444
rect 63368 553432 63374 553444
rect 66898 553432 66904 553444
rect 63368 553404 66904 553432
rect 63368 553392 63374 553404
rect 66898 553392 66904 553404
rect 66956 553392 66962 553444
rect 96982 552032 96988 552084
rect 97040 552072 97046 552084
rect 112530 552072 112536 552084
rect 97040 552044 112536 552072
rect 97040 552032 97046 552044
rect 112530 552032 112536 552044
rect 112588 552032 112594 552084
rect 96614 551828 96620 551880
rect 96672 551868 96678 551880
rect 96890 551868 96896 551880
rect 96672 551840 96896 551868
rect 96672 551828 96678 551840
rect 96890 551828 96896 551840
rect 96948 551828 96954 551880
rect 97442 549312 97448 549364
rect 97500 549352 97506 549364
rect 100754 549352 100760 549364
rect 97500 549324 100760 549352
rect 97500 549312 97506 549324
rect 100754 549312 100760 549324
rect 100812 549312 100818 549364
rect 53742 549244 53748 549296
rect 53800 549284 53806 549296
rect 66714 549284 66720 549296
rect 53800 549256 66720 549284
rect 53800 549244 53806 549256
rect 66714 549244 66720 549256
rect 66772 549244 66778 549296
rect 55122 546456 55128 546508
rect 55180 546496 55186 546508
rect 66806 546496 66812 546508
rect 55180 546468 66812 546496
rect 55180 546456 55186 546468
rect 66806 546456 66812 546468
rect 66864 546456 66870 546508
rect 59170 545096 59176 545148
rect 59228 545136 59234 545148
rect 66806 545136 66812 545148
rect 59228 545108 66812 545136
rect 59228 545096 59234 545108
rect 66806 545096 66812 545108
rect 66864 545096 66870 545148
rect 97074 543736 97080 543788
rect 97132 543776 97138 543788
rect 108390 543776 108396 543788
rect 97132 543748 108396 543776
rect 97132 543736 97138 543748
rect 108390 543736 108396 543748
rect 108448 543736 108454 543788
rect 11698 543668 11704 543720
rect 11756 543708 11762 543720
rect 67634 543708 67640 543720
rect 11756 543680 67640 543708
rect 11756 543668 11762 543680
rect 67634 543668 67640 543680
rect 67692 543708 67698 543720
rect 68370 543708 68376 543720
rect 67692 543680 68376 543708
rect 67692 543668 67698 543680
rect 68370 543668 68376 543680
rect 68428 543668 68434 543720
rect 97074 542376 97080 542428
rect 97132 542416 97138 542428
rect 125686 542416 125692 542428
rect 97132 542388 125692 542416
rect 97132 542376 97138 542388
rect 125686 542376 125692 542388
rect 125744 542376 125750 542428
rect 14458 541628 14464 541680
rect 14516 541668 14522 541680
rect 42794 541668 42800 541680
rect 14516 541640 42800 541668
rect 14516 541628 14522 541640
rect 42794 541628 42800 541640
rect 42852 541628 42858 541680
rect 42794 540948 42800 541000
rect 42852 540988 42858 541000
rect 43990 540988 43996 541000
rect 42852 540960 43996 540988
rect 42852 540948 42858 540960
rect 43990 540948 43996 540960
rect 44048 540988 44054 541000
rect 66622 540988 66628 541000
rect 44048 540960 66628 540988
rect 44048 540948 44054 540960
rect 66622 540948 66628 540960
rect 66680 540948 66686 541000
rect 96614 540948 96620 541000
rect 96672 540988 96678 541000
rect 130378 540988 130384 541000
rect 96672 540960 130384 540988
rect 96672 540948 96678 540960
rect 130378 540948 130384 540960
rect 130436 540948 130442 541000
rect 3418 540200 3424 540252
rect 3476 540240 3482 540252
rect 3476 540212 64874 540240
rect 3476 540200 3482 540212
rect 64846 539832 64874 540212
rect 69382 539832 69388 539844
rect 64846 539804 69388 539832
rect 69382 539792 69388 539804
rect 69440 539792 69446 539844
rect 91002 539792 91008 539844
rect 91060 539832 91066 539844
rect 96798 539832 96804 539844
rect 91060 539804 96804 539832
rect 91060 539792 91066 539804
rect 96798 539792 96804 539804
rect 96856 539792 96862 539844
rect 70302 539656 70308 539708
rect 70360 539696 70366 539708
rect 76558 539696 76564 539708
rect 70360 539668 76564 539696
rect 70360 539656 70366 539668
rect 76558 539656 76564 539668
rect 76616 539656 76622 539708
rect 86586 539588 86592 539640
rect 86644 539628 86650 539640
rect 94314 539628 94320 539640
rect 86644 539600 94320 539628
rect 86644 539588 86650 539600
rect 94314 539588 94320 539600
rect 94372 539588 94378 539640
rect 67266 539044 67272 539096
rect 67324 539084 67330 539096
rect 71866 539084 71872 539096
rect 67324 539056 71872 539084
rect 67324 539044 67330 539056
rect 71866 539044 71872 539056
rect 71924 539044 71930 539096
rect 11698 538228 11704 538280
rect 11756 538268 11762 538280
rect 93946 538268 93952 538280
rect 11756 538240 93952 538268
rect 11756 538228 11762 538240
rect 93946 538228 93952 538240
rect 94004 538228 94010 538280
rect 4798 538160 4804 538212
rect 4856 538200 4862 538212
rect 70670 538200 70676 538212
rect 4856 538172 70676 538200
rect 4856 538160 4862 538172
rect 70670 538160 70676 538172
rect 70728 538160 70734 538212
rect 70670 536800 70676 536852
rect 70728 536840 70734 536852
rect 71038 536840 71044 536852
rect 70728 536812 71044 536840
rect 70728 536800 70734 536812
rect 71038 536800 71044 536812
rect 71096 536800 71102 536852
rect 7558 536732 7564 536784
rect 7616 536772 7622 536784
rect 73522 536772 73528 536784
rect 7616 536744 73528 536772
rect 7616 536732 7622 536744
rect 73522 536732 73528 536744
rect 73580 536732 73586 536784
rect 68922 536120 68928 536172
rect 68980 536160 68986 536172
rect 80698 536160 80704 536172
rect 68980 536132 80704 536160
rect 68980 536120 68986 536132
rect 80698 536120 80704 536132
rect 80756 536120 80762 536172
rect 82814 536120 82820 536172
rect 82872 536160 82878 536172
rect 87598 536160 87604 536172
rect 82872 536132 87604 536160
rect 82872 536120 82878 536132
rect 87598 536120 87604 536132
rect 87656 536120 87662 536172
rect 93394 536120 93400 536172
rect 93452 536160 93458 536172
rect 98638 536160 98644 536172
rect 93452 536132 98644 536160
rect 93452 536120 93458 536132
rect 98638 536120 98644 536132
rect 98696 536120 98702 536172
rect 73522 536052 73528 536104
rect 73580 536092 73586 536104
rect 77938 536092 77944 536104
rect 73580 536064 77944 536092
rect 73580 536052 73586 536064
rect 77938 536052 77944 536064
rect 77996 536052 78002 536104
rect 80054 536052 80060 536104
rect 80112 536092 80118 536104
rect 93118 536092 93124 536104
rect 80112 536064 93124 536092
rect 80112 536052 80118 536064
rect 93118 536052 93124 536064
rect 93176 536052 93182 536104
rect 88978 535440 88984 535492
rect 89036 535480 89042 535492
rect 91094 535480 91100 535492
rect 89036 535452 91100 535480
rect 89036 535440 89042 535452
rect 91094 535440 91100 535452
rect 91152 535440 91158 535492
rect 67818 534692 67824 534744
rect 67876 534732 67882 534744
rect 83458 534732 83464 534744
rect 67876 534704 83464 534732
rect 67876 534692 67882 534704
rect 83458 534692 83464 534704
rect 83516 534692 83522 534744
rect 48222 533332 48228 533384
rect 48280 533372 48286 533384
rect 76742 533372 76748 533384
rect 48280 533344 76748 533372
rect 48280 533332 48286 533344
rect 76742 533332 76748 533344
rect 76800 533332 76806 533384
rect 78306 533332 78312 533384
rect 78364 533372 78370 533384
rect 111150 533372 111156 533384
rect 78364 533344 111156 533372
rect 78364 533332 78370 533344
rect 111150 533332 111156 533344
rect 111208 533332 111214 533384
rect 64782 531972 64788 532024
rect 64840 532012 64846 532024
rect 96890 532012 96896 532024
rect 64840 531984 96896 532012
rect 64840 531972 64846 531984
rect 96890 531972 96896 531984
rect 96948 531972 96954 532024
rect 67358 530612 67364 530664
rect 67416 530652 67422 530664
rect 147674 530652 147680 530664
rect 67416 530624 147680 530652
rect 67416 530612 67422 530624
rect 147674 530612 147680 530624
rect 147732 530612 147738 530664
rect 3510 530544 3516 530596
rect 3568 530584 3574 530596
rect 97994 530584 98000 530596
rect 3568 530556 98000 530584
rect 3568 530544 3574 530556
rect 97994 530544 98000 530556
rect 98052 530544 98058 530596
rect 50890 529184 50896 529236
rect 50948 529224 50954 529236
rect 84194 529224 84200 529236
rect 50948 529196 84200 529224
rect 50948 529184 50954 529196
rect 84194 529184 84200 529196
rect 84252 529184 84258 529236
rect 64690 527824 64696 527876
rect 64748 527864 64754 527876
rect 115934 527864 115940 527876
rect 64748 527836 115940 527864
rect 64748 527824 64754 527836
rect 115934 527824 115940 527836
rect 115992 527824 115998 527876
rect 3418 526396 3424 526448
rect 3476 526436 3482 526448
rect 94498 526436 94504 526448
rect 3476 526408 94504 526436
rect 3476 526396 3482 526408
rect 94498 526396 94504 526408
rect 94556 526396 94562 526448
rect 95142 525784 95148 525836
rect 95200 525824 95206 525836
rect 95418 525824 95424 525836
rect 95200 525796 95424 525824
rect 95200 525784 95206 525796
rect 95418 525784 95424 525796
rect 95476 525784 95482 525836
rect 71774 525036 71780 525088
rect 71832 525076 71838 525088
rect 136726 525076 136732 525088
rect 71832 525048 136732 525076
rect 71832 525036 71838 525048
rect 136726 525036 136732 525048
rect 136784 525036 136790 525088
rect 85666 522384 85672 522436
rect 85724 522424 85730 522436
rect 105538 522424 105544 522436
rect 85724 522396 105544 522424
rect 85724 522384 85730 522396
rect 105538 522384 105544 522396
rect 105596 522384 105602 522436
rect 61930 522248 61936 522300
rect 61988 522288 61994 522300
rect 85666 522288 85672 522300
rect 61988 522260 85672 522288
rect 61988 522248 61994 522260
rect 85666 522248 85672 522260
rect 85724 522248 85730 522300
rect 59078 518168 59084 518220
rect 59136 518208 59142 518220
rect 100846 518208 100852 518220
rect 59136 518180 100852 518208
rect 59136 518168 59142 518180
rect 100846 518168 100852 518180
rect 100904 518168 100910 518220
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 21358 514808 21364 514820
rect 3568 514780 21364 514808
rect 3568 514768 3574 514780
rect 21358 514768 21364 514780
rect 21416 514768 21422 514820
rect 71038 497428 71044 497480
rect 71096 497468 71102 497480
rect 120718 497468 120724 497480
rect 71096 497440 120724 497468
rect 71096 497428 71102 497440
rect 120718 497428 120724 497440
rect 120776 497428 120782 497480
rect 85574 494708 85580 494760
rect 85632 494748 85638 494760
rect 118786 494748 118792 494760
rect 85632 494720 118792 494748
rect 85632 494708 85638 494720
rect 118786 494708 118792 494720
rect 118844 494708 118850 494760
rect 73154 493280 73160 493332
rect 73212 493320 73218 493332
rect 133874 493320 133880 493332
rect 73212 493292 133880 493320
rect 73212 493280 73218 493292
rect 133874 493280 133880 493292
rect 133932 493280 133938 493332
rect 65978 490560 65984 490612
rect 66036 490600 66042 490612
rect 92566 490600 92572 490612
rect 66036 490572 92572 490600
rect 66036 490560 66042 490572
rect 92566 490560 92572 490572
rect 92624 490560 92630 490612
rect 77938 487772 77944 487824
rect 77996 487812 78002 487824
rect 102870 487812 102876 487824
rect 77996 487784 102876 487812
rect 77996 487772 78002 487784
rect 102870 487772 102876 487784
rect 102928 487772 102934 487824
rect 80698 486412 80704 486464
rect 80756 486452 80762 486464
rect 99466 486452 99472 486464
rect 80756 486424 99472 486452
rect 80756 486412 80762 486424
rect 99466 486412 99472 486424
rect 99524 486412 99530 486464
rect 188982 484372 188988 484424
rect 189040 484412 189046 484424
rect 580166 484412 580172 484424
rect 189040 484384 580172 484412
rect 189040 484372 189046 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 67818 484304 67824 484356
rect 67876 484344 67882 484356
rect 69014 484344 69020 484356
rect 67876 484316 69020 484344
rect 67876 484304 67882 484316
rect 69014 484304 69020 484316
rect 69072 484304 69078 484356
rect 106918 483624 106924 483676
rect 106976 483664 106982 483676
rect 131114 483664 131120 483676
rect 106976 483636 131120 483664
rect 106976 483624 106982 483636
rect 131114 483624 131120 483636
rect 131172 483624 131178 483676
rect 77294 482264 77300 482316
rect 77352 482304 77358 482316
rect 88978 482304 88984 482316
rect 77352 482276 88984 482304
rect 77352 482264 77358 482276
rect 88978 482264 88984 482276
rect 89036 482264 89042 482316
rect 258166 481584 258172 481636
rect 258224 481624 258230 481636
rect 258718 481624 258724 481636
rect 258224 481596 258724 481624
rect 258224 481584 258230 481596
rect 258718 481584 258724 481596
rect 258776 481584 258782 481636
rect 93118 480904 93124 480956
rect 93176 480944 93182 480956
rect 121546 480944 121552 480956
rect 93176 480916 121552 480944
rect 93176 480904 93182 480916
rect 121546 480904 121552 480916
rect 121604 480904 121610 480956
rect 122742 480224 122748 480276
rect 122800 480264 122806 480276
rect 258166 480264 258172 480276
rect 122800 480236 258172 480264
rect 122800 480224 122806 480236
rect 258166 480224 258172 480236
rect 258224 480224 258230 480276
rect 110414 478864 110420 478916
rect 110472 478904 110478 478916
rect 111058 478904 111064 478916
rect 110472 478876 111064 478904
rect 110472 478864 110478 478876
rect 111058 478864 111064 478876
rect 111116 478904 111122 478916
rect 251818 478904 251824 478916
rect 111116 478876 251824 478904
rect 111116 478864 111122 478876
rect 251818 478864 251824 478876
rect 251876 478864 251882 478916
rect 98730 478116 98736 478168
rect 98788 478156 98794 478168
rect 124306 478156 124312 478168
rect 98788 478128 124312 478156
rect 98788 478116 98794 478128
rect 124306 478116 124312 478128
rect 124364 478116 124370 478168
rect 48130 477504 48136 477556
rect 48188 477544 48194 477556
rect 202138 477544 202144 477556
rect 48188 477516 202144 477544
rect 48188 477504 48194 477516
rect 202138 477504 202144 477516
rect 202196 477504 202202 477556
rect 85574 476756 85580 476808
rect 85632 476796 85638 476808
rect 95234 476796 95240 476808
rect 85632 476768 95240 476796
rect 85632 476756 85638 476768
rect 95234 476756 95240 476768
rect 95292 476756 95298 476808
rect 8202 476076 8208 476128
rect 8260 476116 8266 476128
rect 11698 476116 11704 476128
rect 8260 476088 11704 476116
rect 8260 476076 8266 476088
rect 11698 476076 11704 476088
rect 11756 476076 11762 476128
rect 109770 476076 109776 476128
rect 109828 476116 109834 476128
rect 249058 476116 249064 476128
rect 109828 476088 249064 476116
rect 109828 476076 109834 476088
rect 249058 476076 249064 476088
rect 249116 476076 249122 476128
rect 59170 476008 59176 476060
rect 59228 476048 59234 476060
rect 122742 476048 122748 476060
rect 59228 476020 122748 476048
rect 59228 476008 59234 476020
rect 122742 476008 122748 476020
rect 122800 476048 122806 476060
rect 123018 476048 123024 476060
rect 122800 476020 123024 476048
rect 122800 476008 122806 476020
rect 123018 476008 123024 476020
rect 123076 476008 123082 476060
rect 3418 475192 3424 475244
rect 3476 475232 3482 475244
rect 7558 475232 7564 475244
rect 3476 475204 7564 475232
rect 3476 475192 3482 475204
rect 7558 475192 7564 475204
rect 7616 475232 7622 475244
rect 8202 475232 8208 475244
rect 7616 475204 8208 475232
rect 7616 475192 7622 475204
rect 8202 475192 8208 475204
rect 8260 475192 8266 475244
rect 104250 474716 104256 474768
rect 104308 474756 104314 474768
rect 238018 474756 238024 474768
rect 104308 474728 238024 474756
rect 104308 474716 104314 474728
rect 238018 474716 238024 474728
rect 238076 474716 238082 474768
rect 90910 473356 90916 473408
rect 90968 473396 90974 473408
rect 226978 473396 226984 473408
rect 90968 473368 226984 473396
rect 90968 473356 90974 473368
rect 226978 473356 226984 473368
rect 227036 473356 227042 473408
rect 94498 473288 94504 473340
rect 94556 473328 94562 473340
rect 95050 473328 95056 473340
rect 94556 473300 95056 473328
rect 94556 473288 94562 473300
rect 95050 473288 95056 473300
rect 95108 473288 95114 473340
rect 202874 472064 202880 472116
rect 202932 472104 202938 472116
rect 295334 472104 295340 472116
rect 202932 472076 295340 472104
rect 202932 472064 202938 472076
rect 295334 472064 295340 472076
rect 295392 472064 295398 472116
rect 95050 471996 95056 472048
rect 95108 472036 95114 472048
rect 231854 472036 231860 472048
rect 95108 472008 231860 472036
rect 95108 471996 95114 472008
rect 231854 471996 231860 472008
rect 231912 471996 231918 472048
rect 240134 471928 240140 471980
rect 240192 471968 240198 471980
rect 240778 471968 240784 471980
rect 240192 471940 240784 471968
rect 240192 471928 240198 471940
rect 240778 471928 240784 471940
rect 240836 471928 240842 471980
rect 102134 471248 102140 471300
rect 102192 471288 102198 471300
rect 102778 471288 102784 471300
rect 102192 471260 102784 471288
rect 102192 471248 102198 471260
rect 102778 471248 102784 471260
rect 102836 471288 102842 471300
rect 240134 471288 240140 471300
rect 102836 471260 240140 471288
rect 102836 471248 102842 471260
rect 240134 471248 240140 471260
rect 240192 471248 240198 471300
rect 155770 470568 155776 470620
rect 155828 470608 155834 470620
rect 251174 470608 251180 470620
rect 155828 470580 251180 470608
rect 155828 470568 155834 470580
rect 251174 470568 251180 470580
rect 251232 470568 251238 470620
rect 70302 469820 70308 469872
rect 70360 469860 70366 469872
rect 91186 469860 91192 469872
rect 70360 469832 91192 469860
rect 70360 469820 70366 469832
rect 91186 469820 91192 469832
rect 91244 469820 91250 469872
rect 105538 469820 105544 469872
rect 105596 469860 105602 469872
rect 241514 469860 241520 469872
rect 105596 469832 241520 469860
rect 105596 469820 105602 469832
rect 241514 469820 241520 469832
rect 241572 469820 241578 469872
rect 241514 469276 241520 469328
rect 241572 469316 241578 469328
rect 242158 469316 242164 469328
rect 241572 469288 242164 469316
rect 241572 469276 241578 469288
rect 242158 469276 242164 469288
rect 242216 469276 242222 469328
rect 85482 469208 85488 469260
rect 85540 469248 85546 469260
rect 86218 469248 86224 469260
rect 85540 469220 86224 469248
rect 85540 469208 85546 469220
rect 86218 469208 86224 469220
rect 86276 469208 86282 469260
rect 104894 469208 104900 469260
rect 104952 469248 104958 469260
rect 105538 469248 105544 469260
rect 104952 469220 105544 469248
rect 104952 469208 104958 469220
rect 105538 469208 105544 469220
rect 105596 469208 105602 469260
rect 123478 469208 123484 469260
rect 123536 469248 123542 469260
rect 255406 469248 255412 469260
rect 123536 469220 255412 469248
rect 123536 469208 123542 469220
rect 255406 469208 255412 469220
rect 255464 469208 255470 469260
rect 111150 468460 111156 468512
rect 111208 468500 111214 468512
rect 117774 468500 117780 468512
rect 111208 468472 117780 468500
rect 111208 468460 111214 468472
rect 117774 468460 117780 468472
rect 117832 468460 117838 468512
rect 227806 467956 227812 467968
rect 103486 467928 227812 467956
rect 93854 467848 93860 467900
rect 93912 467888 93918 467900
rect 95142 467888 95148 467900
rect 93912 467860 95148 467888
rect 93912 467848 93918 467860
rect 95142 467848 95148 467860
rect 95200 467888 95206 467900
rect 103486 467888 103514 467928
rect 227806 467916 227812 467928
rect 227864 467916 227870 467968
rect 95200 467860 103514 467888
rect 95200 467848 95206 467860
rect 117406 467848 117412 467900
rect 117464 467888 117470 467900
rect 117774 467888 117780 467900
rect 117464 467860 117780 467888
rect 117464 467848 117470 467860
rect 117774 467848 117780 467860
rect 117832 467888 117838 467900
rect 258258 467888 258264 467900
rect 117832 467860 258264 467888
rect 117832 467848 117838 467860
rect 258258 467848 258264 467860
rect 258316 467848 258322 467900
rect 164142 466488 164148 466540
rect 164200 466528 164206 466540
rect 242894 466528 242900 466540
rect 164200 466500 242900 466528
rect 164200 466488 164206 466500
rect 242894 466488 242900 466500
rect 242952 466488 242958 466540
rect 112530 466420 112536 466472
rect 112588 466460 112594 466472
rect 142062 466460 142068 466472
rect 112588 466432 142068 466460
rect 112588 466420 112594 466432
rect 142062 466420 142068 466432
rect 142120 466460 142126 466472
rect 252554 466460 252560 466472
rect 142120 466432 252560 466460
rect 142120 466420 142126 466432
rect 252554 466420 252560 466432
rect 252612 466420 252618 466472
rect 170490 465128 170496 465180
rect 170548 465168 170554 465180
rect 259546 465168 259552 465180
rect 170548 465140 259552 465168
rect 170548 465128 170554 465140
rect 259546 465128 259552 465140
rect 259604 465128 259610 465180
rect 142798 465060 142804 465112
rect 142856 465100 142862 465112
rect 245654 465100 245660 465112
rect 142856 465072 245660 465100
rect 142856 465060 142862 465072
rect 245654 465060 245660 465072
rect 245712 465060 245718 465112
rect 119338 463768 119344 463820
rect 119396 463808 119402 463820
rect 255314 463808 255320 463820
rect 119396 463780 255320 463808
rect 119396 463768 119402 463780
rect 255314 463768 255320 463780
rect 255372 463768 255378 463820
rect 115198 463700 115204 463752
rect 115256 463740 115262 463752
rect 262214 463740 262220 463752
rect 115256 463712 262220 463740
rect 115256 463700 115262 463712
rect 262214 463700 262220 463712
rect 262272 463700 262278 463752
rect 212626 463632 212632 463684
rect 212684 463672 212690 463684
rect 213178 463672 213184 463684
rect 212684 463644 213184 463672
rect 212684 463632 212690 463644
rect 213178 463632 213184 463644
rect 213236 463632 213242 463684
rect 67634 463020 67640 463072
rect 67692 463060 67698 463072
rect 81342 463060 81348 463072
rect 67692 463032 81348 463060
rect 67692 463020 67698 463032
rect 81342 463020 81348 463032
rect 81400 463020 81406 463072
rect 80054 462952 80060 463004
rect 80112 462992 80118 463004
rect 113266 462992 113272 463004
rect 80112 462964 113272 462992
rect 80112 462952 80118 462964
rect 113266 462952 113272 462964
rect 113324 462952 113330 463004
rect 184198 462408 184204 462460
rect 184256 462448 184262 462460
rect 212626 462448 212632 462460
rect 184256 462420 212632 462448
rect 184256 462408 184262 462420
rect 212626 462408 212632 462420
rect 212684 462408 212690 462460
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 11698 462380 11704 462392
rect 3292 462352 11704 462380
rect 3292 462340 3298 462352
rect 11698 462340 11704 462352
rect 11756 462340 11762 462392
rect 64782 462340 64788 462392
rect 64840 462380 64846 462392
rect 186958 462380 186964 462392
rect 64840 462352 186964 462380
rect 64840 462340 64846 462352
rect 186958 462340 186964 462352
rect 187016 462340 187022 462392
rect 187050 462340 187056 462392
rect 187108 462380 187114 462392
rect 260834 462380 260840 462392
rect 187108 462352 260840 462380
rect 187108 462340 187114 462352
rect 260834 462340 260840 462352
rect 260892 462340 260898 462392
rect 215386 462272 215392 462324
rect 215444 462312 215450 462324
rect 215938 462312 215944 462324
rect 215444 462284 215944 462312
rect 215444 462272 215450 462284
rect 215938 462272 215944 462284
rect 215996 462272 216002 462324
rect 78674 461592 78680 461644
rect 78732 461632 78738 461644
rect 91738 461632 91744 461644
rect 78732 461604 91744 461632
rect 78732 461592 78738 461604
rect 91738 461592 91744 461604
rect 91796 461592 91802 461644
rect 286318 461592 286324 461644
rect 286376 461632 286382 461644
rect 583294 461632 583300 461644
rect 286376 461604 583300 461632
rect 286376 461592 286382 461604
rect 583294 461592 583300 461604
rect 583352 461592 583358 461644
rect 201494 461320 201500 461372
rect 201552 461360 201558 461372
rect 202138 461360 202144 461372
rect 201552 461332 202144 461360
rect 201552 461320 201558 461332
rect 202138 461320 202144 461332
rect 202196 461320 202202 461372
rect 182818 460980 182824 461032
rect 182876 461020 182882 461032
rect 215386 461020 215392 461032
rect 182876 460992 215392 461020
rect 182876 460980 182882 460992
rect 215386 460980 215392 460992
rect 215444 460980 215450 461032
rect 62022 460912 62028 460964
rect 62080 460952 62086 460964
rect 185578 460952 185584 460964
rect 62080 460924 185584 460952
rect 62080 460912 62086 460924
rect 185578 460912 185584 460924
rect 185636 460912 185642 460964
rect 202138 460912 202144 460964
rect 202196 460952 202202 460964
rect 286318 460952 286324 460964
rect 202196 460924 286324 460952
rect 202196 460912 202202 460924
rect 286318 460912 286324 460924
rect 286376 460912 286382 460964
rect 87598 460844 87604 460896
rect 87656 460884 87662 460896
rect 109034 460884 109040 460896
rect 87656 460856 109040 460884
rect 87656 460844 87662 460856
rect 109034 460844 109040 460856
rect 109092 460844 109098 460896
rect 109034 460164 109040 460216
rect 109092 460204 109098 460216
rect 109770 460204 109776 460216
rect 109092 460176 109776 460204
rect 109092 460164 109098 460176
rect 109770 460164 109776 460176
rect 109828 460164 109834 460216
rect 141418 459620 141424 459672
rect 141476 459660 141482 459672
rect 256786 459660 256792 459672
rect 141476 459632 256792 459660
rect 141476 459620 141482 459632
rect 256786 459620 256792 459632
rect 256844 459620 256850 459672
rect 81342 459552 81348 459604
rect 81400 459592 81406 459604
rect 208394 459592 208400 459604
rect 81400 459564 208400 459592
rect 81400 459552 81406 459564
rect 208394 459552 208400 459564
rect 208452 459552 208458 459604
rect 226978 459552 226984 459604
rect 227036 459592 227042 459604
rect 227622 459592 227628 459604
rect 227036 459564 227628 459592
rect 227036 459552 227042 459564
rect 227622 459552 227628 459564
rect 227680 459592 227686 459604
rect 258350 459592 258356 459604
rect 227680 459564 258356 459592
rect 227680 459552 227686 459564
rect 258350 459552 258356 459564
rect 258408 459552 258414 459604
rect 77202 458804 77208 458856
rect 77260 458844 77266 458856
rect 90358 458844 90364 458856
rect 77260 458816 90364 458844
rect 77260 458804 77266 458816
rect 90358 458804 90364 458816
rect 90416 458804 90422 458856
rect 95234 458260 95240 458312
rect 95292 458300 95298 458312
rect 195790 458300 195796 458312
rect 95292 458272 195796 458300
rect 95292 458260 95298 458272
rect 195790 458260 195796 458272
rect 195848 458300 195854 458312
rect 227714 458300 227720 458312
rect 195848 458272 227720 458300
rect 195848 458260 195854 458272
rect 227714 458260 227720 458272
rect 227772 458260 227778 458312
rect 237374 458260 237380 458312
rect 237432 458300 237438 458312
rect 291194 458300 291200 458312
rect 237432 458272 291200 458300
rect 237432 458260 237438 458272
rect 291194 458260 291200 458272
rect 291252 458260 291258 458312
rect 111702 458192 111708 458244
rect 111760 458232 111766 458244
rect 259454 458232 259460 458244
rect 111760 458204 259460 458232
rect 111760 458192 111766 458204
rect 259454 458192 259460 458204
rect 259512 458192 259518 458244
rect 193398 456832 193404 456884
rect 193456 456872 193462 456884
rect 218974 456872 218980 456884
rect 193456 456844 218980 456872
rect 193456 456832 193462 456844
rect 218974 456832 218980 456844
rect 219032 456832 219038 456884
rect 78674 456764 78680 456816
rect 78732 456804 78738 456816
rect 173618 456804 173624 456816
rect 78732 456776 173624 456804
rect 78732 456764 78738 456776
rect 173618 456764 173624 456776
rect 173676 456804 173682 456816
rect 173802 456804 173808 456816
rect 173676 456776 173808 456804
rect 173676 456764 173682 456776
rect 173802 456764 173808 456776
rect 173860 456764 173866 456816
rect 179322 456764 179328 456816
rect 179380 456804 179386 456816
rect 204530 456804 204536 456816
rect 179380 456776 204536 456804
rect 179380 456764 179386 456776
rect 204530 456764 204536 456776
rect 204588 456764 204594 456816
rect 230474 456764 230480 456816
rect 230532 456804 230538 456816
rect 287146 456804 287152 456816
rect 230532 456776 287152 456804
rect 230532 456764 230538 456776
rect 287146 456764 287152 456776
rect 287204 456804 287210 456816
rect 580166 456804 580172 456816
rect 287204 456776 580172 456804
rect 287204 456764 287210 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 251174 456084 251180 456136
rect 251232 456124 251238 456136
rect 252094 456124 252100 456136
rect 251232 456096 252100 456124
rect 251232 456084 251238 456096
rect 252094 456084 252100 456096
rect 252152 456084 252158 456136
rect 238018 456016 238024 456068
rect 238076 456056 238082 456068
rect 241514 456056 241520 456068
rect 238076 456028 241520 456056
rect 238076 456016 238082 456028
rect 241514 456016 241520 456028
rect 241572 456016 241578 456068
rect 72418 455472 72424 455524
rect 72476 455512 72482 455524
rect 160094 455512 160100 455524
rect 72476 455484 160100 455512
rect 72476 455472 72482 455484
rect 160094 455472 160100 455484
rect 160152 455512 160158 455524
rect 197354 455512 197360 455524
rect 160152 455484 197360 455512
rect 160152 455472 160158 455484
rect 197354 455472 197360 455484
rect 197412 455472 197418 455524
rect 225506 455472 225512 455524
rect 225564 455512 225570 455524
rect 261478 455512 261484 455524
rect 225564 455484 261484 455512
rect 225564 455472 225570 455484
rect 261478 455472 261484 455484
rect 261536 455472 261542 455524
rect 97994 455404 98000 455456
rect 98052 455444 98058 455456
rect 233234 455444 233240 455456
rect 98052 455416 233240 455444
rect 98052 455404 98058 455416
rect 233234 455404 233240 455416
rect 233292 455404 233298 455456
rect 82814 455336 82820 455388
rect 82872 455376 82878 455388
rect 111702 455376 111708 455388
rect 82872 455348 111708 455376
rect 82872 455336 82878 455348
rect 111702 455336 111708 455348
rect 111760 455376 111766 455388
rect 112714 455376 112720 455388
rect 111760 455348 112720 455376
rect 111760 455336 111766 455348
rect 112714 455336 112720 455348
rect 112772 455336 112778 455388
rect 191190 454112 191196 454164
rect 191248 454152 191254 454164
rect 218146 454152 218152 454164
rect 191248 454124 218152 454152
rect 191248 454112 191254 454124
rect 218146 454112 218152 454124
rect 218204 454112 218210 454164
rect 76558 454044 76564 454096
rect 76616 454084 76622 454096
rect 159450 454084 159456 454096
rect 76616 454056 159456 454084
rect 76616 454044 76622 454056
rect 159450 454044 159456 454056
rect 159508 454084 159514 454096
rect 200114 454084 200120 454096
rect 159508 454056 200120 454084
rect 159508 454044 159514 454056
rect 200114 454044 200120 454056
rect 200172 454044 200178 454096
rect 222562 454044 222568 454096
rect 222620 454084 222626 454096
rect 266998 454084 267004 454096
rect 222620 454056 267004 454084
rect 222620 454044 222626 454056
rect 266998 454044 267004 454056
rect 267056 454044 267062 454096
rect 227622 453976 227628 454028
rect 227680 454016 227686 454028
rect 228726 454016 228732 454028
rect 227680 453988 228732 454016
rect 227680 453976 227686 453988
rect 228726 453976 228732 453988
rect 228784 453976 228790 454028
rect 212718 453364 212724 453416
rect 212776 453404 212782 453416
rect 215478 453404 215484 453416
rect 212776 453376 215484 453404
rect 212776 453364 212782 453376
rect 215478 453364 215484 453376
rect 215536 453364 215542 453416
rect 195974 453296 195980 453348
rect 196032 453336 196038 453348
rect 212442 453336 212448 453348
rect 196032 453308 212448 453336
rect 196032 453296 196038 453308
rect 212442 453296 212448 453308
rect 212500 453296 212506 453348
rect 193306 452752 193312 452804
rect 193364 452792 193370 452804
rect 213638 452792 213644 452804
rect 193364 452764 213644 452792
rect 193364 452752 193370 452764
rect 213638 452752 213644 452764
rect 213696 452752 213702 452804
rect 251818 452752 251824 452804
rect 251876 452792 251882 452804
rect 268378 452792 268384 452804
rect 251876 452764 268384 452792
rect 251876 452752 251882 452764
rect 268378 452752 268384 452764
rect 268436 452752 268442 452804
rect 222102 452684 222108 452736
rect 222160 452724 222166 452736
rect 251450 452724 251456 452736
rect 222160 452696 251456 452724
rect 222160 452684 222166 452696
rect 251450 452684 251456 452696
rect 251508 452684 251514 452736
rect 60458 452616 60464 452668
rect 60516 452656 60522 452668
rect 170398 452656 170404 452668
rect 60516 452628 170404 452656
rect 60516 452616 60522 452628
rect 170398 452616 170404 452628
rect 170456 452616 170462 452668
rect 192478 452616 192484 452668
rect 192536 452656 192542 452668
rect 196526 452656 196532 452668
rect 192536 452628 196532 452656
rect 192536 452616 192542 452628
rect 196526 452616 196532 452628
rect 196584 452616 196590 452668
rect 211246 452616 211252 452668
rect 211304 452656 211310 452668
rect 226886 452656 226892 452668
rect 211304 452628 226892 452656
rect 211304 452616 211310 452628
rect 226886 452616 226892 452628
rect 226944 452616 226950 452668
rect 227714 452616 227720 452668
rect 227772 452656 227778 452668
rect 229646 452656 229652 452668
rect 227772 452628 229652 452656
rect 227772 452616 227778 452628
rect 229646 452616 229652 452628
rect 229704 452616 229710 452668
rect 237374 452616 237380 452668
rect 237432 452656 237438 452668
rect 274634 452656 274640 452668
rect 237432 452628 274640 452656
rect 237432 452616 237438 452628
rect 274634 452616 274640 452628
rect 274692 452616 274698 452668
rect 82722 451936 82728 451988
rect 82780 451976 82786 451988
rect 122834 451976 122840 451988
rect 82780 451948 122840 451976
rect 82780 451936 82786 451948
rect 122834 451936 122840 451948
rect 122892 451976 122898 451988
rect 124122 451976 124128 451988
rect 122892 451948 124128 451976
rect 122892 451936 122898 451948
rect 124122 451936 124128 451948
rect 124180 451936 124186 451988
rect 87598 451868 87604 451920
rect 87656 451908 87662 451920
rect 187602 451908 187608 451920
rect 87656 451880 187608 451908
rect 87656 451868 87662 451880
rect 187602 451868 187608 451880
rect 187660 451908 187666 451920
rect 188338 451908 188344 451920
rect 187660 451880 188344 451908
rect 187660 451868 187666 451880
rect 188338 451868 188344 451880
rect 188396 451868 188402 451920
rect 240226 451392 240232 451444
rect 240284 451432 240290 451444
rect 240284 451404 248414 451432
rect 240284 451392 240290 451404
rect 189810 451324 189816 451376
rect 189868 451364 189874 451376
rect 241054 451364 241060 451376
rect 189868 451336 241060 451364
rect 189868 451324 189874 451336
rect 241054 451324 241060 451336
rect 241112 451324 241118 451376
rect 248386 451364 248414 451404
rect 256694 451364 256700 451376
rect 248386 451336 256700 451364
rect 256694 451324 256700 451336
rect 256752 451324 256758 451376
rect 191834 451256 191840 451308
rect 191892 451296 191898 451308
rect 199286 451296 199292 451308
rect 191892 451268 199292 451296
rect 191892 451256 191898 451268
rect 199286 451256 199292 451268
rect 199344 451256 199350 451308
rect 210418 451256 210424 451308
rect 210476 451296 210482 451308
rect 583294 451296 583300 451308
rect 210476 451268 583300 451296
rect 210476 451256 210482 451268
rect 583294 451256 583300 451268
rect 583352 451256 583358 451308
rect 101398 450508 101404 450560
rect 101456 450548 101462 450560
rect 117958 450548 117964 450560
rect 101456 450520 117964 450548
rect 101456 450508 101462 450520
rect 117958 450508 117964 450520
rect 118016 450508 118022 450560
rect 192570 450508 192576 450560
rect 192628 450548 192634 450560
rect 211246 450548 211252 450560
rect 192628 450520 211252 450548
rect 192628 450508 192634 450520
rect 211246 450508 211252 450520
rect 211304 450508 211310 450560
rect 231854 449964 231860 450016
rect 231912 450004 231918 450016
rect 232866 450004 232872 450016
rect 231912 449976 232872 450004
rect 231912 449964 231918 449976
rect 232866 449964 232872 449976
rect 232924 450004 232930 450016
rect 267734 450004 267740 450016
rect 232924 449976 267740 450004
rect 232924 449964 232930 449976
rect 267734 449964 267740 449976
rect 267792 449964 267798 450016
rect 59262 449896 59268 449948
rect 59320 449936 59326 449948
rect 151078 449936 151084 449948
rect 59320 449908 151084 449936
rect 59320 449896 59326 449908
rect 151078 449896 151084 449908
rect 151136 449896 151142 449948
rect 178678 449896 178684 449948
rect 178736 449936 178742 449948
rect 240226 449936 240232 449948
rect 178736 449908 240232 449936
rect 178736 449896 178742 449908
rect 240226 449896 240232 449908
rect 240284 449896 240290 449948
rect 242434 449896 242440 449948
rect 242492 449936 242498 449948
rect 254578 449936 254584 449948
rect 242492 449908 254584 449936
rect 242492 449896 242498 449908
rect 254578 449896 254584 449908
rect 254636 449896 254642 449948
rect 73798 449828 73804 449880
rect 73856 449868 73862 449880
rect 200942 449868 200948 449880
rect 73856 449840 200948 449868
rect 73856 449828 73862 449840
rect 200942 449828 200948 449840
rect 201000 449828 201006 449880
rect 3234 449760 3240 449812
rect 3292 449800 3298 449812
rect 100754 449800 100760 449812
rect 3292 449772 100760 449800
rect 3292 449760 3298 449772
rect 100754 449760 100760 449772
rect 100812 449760 100818 449812
rect 251450 449692 251456 449744
rect 251508 449732 251514 449744
rect 251508 449704 251680 449732
rect 251508 449692 251514 449704
rect 173802 449148 173808 449200
rect 173860 449188 173866 449200
rect 193398 449188 193404 449200
rect 173860 449160 193404 449188
rect 173860 449148 173866 449160
rect 193398 449148 193404 449160
rect 193456 449148 193462 449200
rect 251652 449188 251680 449704
rect 255498 449216 255504 449268
rect 255556 449256 255562 449268
rect 271230 449256 271236 449268
rect 255556 449228 271236 449256
rect 255556 449216 255562 449228
rect 271230 449216 271236 449228
rect 271288 449216 271294 449268
rect 269114 449188 269120 449200
rect 251652 449160 269120 449188
rect 269114 449148 269120 449160
rect 269172 449148 269178 449200
rect 64690 448536 64696 448588
rect 64748 448576 64754 448588
rect 74534 448576 74540 448588
rect 64748 448548 74540 448576
rect 64748 448536 64754 448548
rect 74534 448536 74540 448548
rect 74592 448576 74598 448588
rect 75822 448576 75828 448588
rect 74592 448548 75828 448576
rect 74592 448536 74598 448548
rect 75822 448536 75828 448548
rect 75880 448536 75886 448588
rect 53650 447856 53656 447908
rect 53708 447896 53714 447908
rect 106918 447896 106924 447908
rect 53708 447868 106924 447896
rect 53708 447856 53714 447868
rect 106918 447856 106924 447868
rect 106976 447856 106982 447908
rect 112438 447856 112444 447908
rect 112496 447896 112502 447908
rect 122926 447896 122932 447908
rect 112496 447868 122932 447896
rect 112496 447856 112502 447868
rect 122926 447856 122932 447868
rect 122984 447856 122990 447908
rect 169018 447856 169024 447908
rect 169076 447896 169082 447908
rect 191650 447896 191656 447908
rect 169076 447868 191656 447896
rect 169076 447856 169082 447868
rect 191650 447856 191656 447868
rect 191708 447856 191714 447908
rect 75822 447788 75828 447840
rect 75880 447828 75886 447840
rect 181438 447828 181444 447840
rect 75880 447800 181444 447828
rect 75880 447788 75886 447800
rect 181438 447788 181444 447800
rect 181496 447788 181502 447840
rect 255406 447788 255412 447840
rect 255464 447828 255470 447840
rect 287054 447828 287060 447840
rect 255464 447800 287060 447828
rect 255464 447788 255470 447800
rect 287054 447788 287060 447800
rect 287112 447788 287118 447840
rect 188430 447108 188436 447160
rect 188488 447148 188494 447160
rect 191006 447148 191012 447160
rect 188488 447120 191012 447148
rect 188488 447108 188494 447120
rect 191006 447108 191012 447120
rect 191064 447108 191070 447160
rect 176562 446360 176568 446412
rect 176620 446400 176626 446412
rect 191834 446400 191840 446412
rect 176620 446372 191840 446400
rect 176620 446360 176626 446372
rect 191834 446360 191840 446372
rect 191892 446360 191898 446412
rect 59170 445816 59176 445868
rect 59228 445856 59234 445868
rect 152458 445856 152464 445868
rect 59228 445828 152464 445856
rect 59228 445816 59234 445828
rect 152458 445816 152464 445828
rect 152516 445816 152522 445868
rect 71130 445748 71136 445800
rect 71188 445788 71194 445800
rect 191650 445788 191656 445800
rect 71188 445760 191656 445788
rect 71188 445748 71194 445760
rect 191650 445748 191656 445760
rect 191708 445748 191714 445800
rect 186314 445680 186320 445732
rect 186372 445720 186378 445732
rect 187602 445720 187608 445732
rect 186372 445692 187608 445720
rect 186372 445680 186378 445692
rect 187602 445680 187608 445692
rect 187660 445720 187666 445732
rect 191190 445720 191196 445732
rect 187660 445692 191196 445720
rect 187660 445680 187666 445692
rect 191190 445680 191196 445692
rect 191248 445680 191254 445732
rect 52270 445000 52276 445052
rect 52328 445040 52334 445052
rect 60550 445040 60556 445052
rect 52328 445012 60556 445040
rect 52328 445000 52334 445012
rect 60550 445000 60556 445012
rect 60608 445000 60614 445052
rect 88242 445000 88248 445052
rect 88300 445040 88306 445052
rect 91002 445040 91008 445052
rect 88300 445012 91008 445040
rect 88300 445000 88306 445012
rect 91002 445000 91008 445012
rect 91060 445040 91066 445052
rect 186314 445040 186320 445052
rect 91060 445012 186320 445040
rect 91060 445000 91066 445012
rect 186314 445000 186320 445012
rect 186372 445000 186378 445052
rect 60550 444388 60556 444440
rect 60608 444428 60614 444440
rect 88518 444428 88524 444440
rect 60608 444400 88524 444428
rect 60608 444388 60614 444400
rect 88518 444388 88524 444400
rect 88576 444388 88582 444440
rect 255406 444388 255412 444440
rect 255464 444428 255470 444440
rect 263778 444428 263784 444440
rect 255464 444400 263784 444428
rect 255464 444388 255470 444400
rect 263778 444388 263784 444400
rect 263836 444388 263842 444440
rect 111886 444320 111892 444372
rect 111944 444360 111950 444372
rect 112530 444360 112536 444372
rect 111944 444332 112536 444360
rect 111944 444320 111950 444332
rect 112530 444320 112536 444332
rect 112588 444320 112594 444372
rect 107654 443776 107660 443828
rect 107712 443816 107718 443828
rect 108390 443816 108396 443828
rect 107712 443788 108396 443816
rect 107712 443776 107718 443788
rect 108390 443776 108396 443788
rect 108448 443816 108454 443828
rect 108448 443788 113174 443816
rect 108448 443776 108454 443788
rect 113146 443680 113174 443788
rect 142798 443680 142804 443692
rect 113146 443652 142804 443680
rect 142798 443640 142804 443652
rect 142856 443640 142862 443692
rect 65978 443504 65984 443556
rect 66036 443544 66042 443556
rect 70486 443544 70492 443556
rect 66036 443516 70492 443544
rect 66036 443504 66042 443516
rect 70486 443504 70492 443516
rect 70544 443504 70550 443556
rect 255406 443368 255412 443420
rect 255464 443408 255470 443420
rect 259454 443408 259460 443420
rect 255464 443380 259460 443408
rect 255464 443368 255470 443380
rect 259454 443368 259460 443380
rect 259512 443368 259518 443420
rect 3418 442960 3424 443012
rect 3476 443000 3482 443012
rect 111886 443000 111892 443012
rect 3476 442972 111892 443000
rect 3476 442960 3482 442972
rect 111886 442960 111892 442972
rect 111944 442960 111950 443012
rect 117314 442892 117320 442944
rect 117372 442932 117378 442944
rect 117774 442932 117780 442944
rect 117372 442904 117780 442932
rect 117372 442892 117378 442904
rect 117774 442892 117780 442904
rect 117832 442932 117838 442944
rect 192478 442932 192484 442944
rect 117832 442904 192484 442932
rect 117832 442892 117838 442904
rect 192478 442892 192484 442904
rect 192536 442892 192542 442944
rect 70394 442212 70400 442264
rect 70452 442252 70458 442264
rect 117774 442252 117780 442264
rect 70452 442224 117780 442252
rect 70452 442212 70458 442224
rect 117774 442212 117780 442224
rect 117832 442212 117838 442264
rect 125686 442076 125692 442128
rect 125744 442116 125750 442128
rect 126238 442116 126244 442128
rect 125744 442088 126244 442116
rect 125744 442076 125750 442088
rect 126238 442076 126244 442088
rect 126296 442076 126302 442128
rect 255406 442008 255412 442060
rect 255464 442048 255470 442060
rect 258166 442048 258172 442060
rect 255464 442020 258172 442048
rect 255464 442008 255470 442020
rect 258166 442008 258172 442020
rect 258224 442048 258230 442060
rect 258718 442048 258724 442060
rect 258224 442020 258724 442048
rect 258224 442008 258230 442020
rect 258718 442008 258724 442020
rect 258776 442008 258782 442060
rect 63218 441600 63224 441652
rect 63276 441640 63282 441652
rect 125686 441640 125692 441652
rect 63276 441612 125692 441640
rect 63276 441600 63282 441612
rect 125686 441600 125692 441612
rect 125744 441600 125750 441652
rect 67082 440852 67088 440904
rect 67140 440892 67146 440904
rect 122834 440892 122840 440904
rect 67140 440864 122840 440892
rect 67140 440852 67146 440864
rect 122834 440852 122840 440864
rect 122892 440852 122898 440904
rect 67358 440240 67364 440292
rect 67416 440280 67422 440292
rect 166350 440280 166356 440292
rect 67416 440252 166356 440280
rect 67416 440240 67422 440252
rect 166350 440240 166356 440252
rect 166408 440240 166414 440292
rect 176654 440240 176660 440292
rect 176712 440280 176718 440292
rect 191374 440280 191380 440292
rect 176712 440252 191380 440280
rect 176712 440240 176718 440252
rect 191374 440240 191380 440252
rect 191432 440240 191438 440292
rect 185762 439492 185768 439544
rect 185820 439532 185826 439544
rect 193306 439532 193312 439544
rect 185820 439504 193312 439532
rect 185820 439492 185826 439504
rect 193306 439492 193312 439504
rect 193364 439492 193370 439544
rect 255314 439492 255320 439544
rect 255372 439532 255378 439544
rect 288526 439532 288532 439544
rect 255372 439504 288532 439532
rect 255372 439492 255378 439504
rect 288526 439492 288532 439504
rect 288584 439532 288590 439544
rect 583018 439532 583024 439544
rect 288584 439504 583024 439532
rect 288584 439492 288590 439504
rect 583018 439492 583024 439504
rect 583076 439492 583082 439544
rect 44082 438948 44088 439000
rect 44140 438988 44146 439000
rect 69658 438988 69664 439000
rect 44140 438960 69664 438988
rect 44140 438948 44146 438960
rect 69658 438948 69664 438960
rect 69716 438948 69722 439000
rect 83458 438948 83464 439000
rect 83516 438988 83522 439000
rect 83734 438988 83740 439000
rect 83516 438960 83740 438988
rect 83516 438948 83522 438960
rect 83734 438948 83740 438960
rect 83792 438988 83798 439000
rect 185762 438988 185768 439000
rect 83792 438960 185768 438988
rect 83792 438948 83798 438960
rect 185762 438948 185768 438960
rect 185820 438988 185826 439000
rect 186130 438988 186136 439000
rect 185820 438960 186136 438988
rect 185820 438948 185826 438960
rect 186130 438948 186136 438960
rect 186188 438948 186194 439000
rect 68278 438880 68284 438932
rect 68336 438920 68342 438932
rect 191374 438920 191380 438932
rect 68336 438892 191380 438920
rect 68336 438880 68342 438892
rect 191374 438880 191380 438892
rect 191432 438880 191438 438932
rect 65978 438132 65984 438184
rect 66036 438172 66042 438184
rect 191558 438172 191564 438184
rect 66036 438144 191564 438172
rect 66036 438132 66042 438144
rect 191558 438132 191564 438144
rect 191616 438132 191622 438184
rect 255406 438132 255412 438184
rect 255464 438172 255470 438184
rect 258258 438172 258264 438184
rect 255464 438144 258264 438172
rect 255464 438132 255470 438144
rect 258258 438132 258264 438144
rect 258316 438172 258322 438184
rect 266354 438172 266360 438184
rect 258316 438144 266360 438172
rect 258316 438132 258322 438144
rect 266354 438132 266360 438144
rect 266412 438132 266418 438184
rect 95050 437588 95056 437640
rect 95108 437628 95114 437640
rect 96982 437628 96988 437640
rect 95108 437600 96988 437628
rect 95108 437588 95114 437600
rect 96982 437588 96988 437600
rect 97040 437588 97046 437640
rect 48130 437452 48136 437504
rect 48188 437492 48194 437504
rect 50982 437492 50988 437504
rect 48188 437464 50988 437492
rect 48188 437452 48194 437464
rect 50982 437452 50988 437464
rect 51040 437492 51046 437504
rect 74810 437492 74816 437504
rect 51040 437464 74816 437492
rect 51040 437452 51046 437464
rect 74810 437452 74816 437464
rect 74868 437452 74874 437504
rect 71682 437384 71688 437436
rect 71740 437424 71746 437436
rect 72418 437424 72424 437436
rect 71740 437396 72424 437424
rect 71740 437384 71746 437396
rect 72418 437384 72424 437396
rect 72476 437384 72482 437436
rect 82814 437384 82820 437436
rect 82872 437424 82878 437436
rect 83918 437424 83924 437436
rect 82872 437396 83924 437424
rect 82872 437384 82878 437396
rect 83918 437384 83924 437396
rect 83976 437424 83982 437436
rect 87598 437424 87604 437436
rect 83976 437396 87604 437424
rect 83976 437384 83982 437396
rect 87598 437384 87604 437396
rect 87656 437384 87662 437436
rect 90910 437384 90916 437436
rect 90968 437424 90974 437436
rect 94222 437424 94228 437436
rect 90968 437396 94228 437424
rect 90968 437384 90974 437396
rect 94222 437384 94228 437396
rect 94280 437384 94286 437436
rect 102870 437384 102876 437436
rect 102928 437424 102934 437436
rect 178678 437424 178684 437436
rect 102928 437396 178684 437424
rect 102928 437384 102934 437396
rect 178678 437384 178684 437396
rect 178736 437384 178742 437436
rect 263410 437384 263416 437436
rect 263468 437424 263474 437436
rect 582466 437424 582472 437436
rect 263468 437396 582472 437424
rect 263468 437384 263474 437396
rect 582466 437384 582472 437396
rect 582524 437384 582530 437436
rect 80974 437316 80980 437368
rect 81032 437356 81038 437368
rect 86218 437356 86224 437368
rect 81032 437328 86224 437356
rect 81032 437316 81038 437328
rect 86218 437316 86224 437328
rect 86276 437316 86282 437368
rect 68922 437112 68928 437164
rect 68980 437152 68986 437164
rect 69750 437152 69756 437164
rect 68980 437124 69756 437152
rect 68980 437112 68986 437124
rect 69750 437112 69756 437124
rect 69808 437112 69814 437164
rect 91738 436704 91744 436756
rect 91796 436744 91802 436756
rect 104434 436744 104440 436756
rect 91796 436716 104440 436744
rect 91796 436704 91802 436716
rect 104434 436704 104440 436716
rect 104492 436704 104498 436756
rect 136634 436704 136640 436756
rect 136692 436744 136698 436756
rect 189810 436744 189816 436756
rect 136692 436716 189816 436744
rect 136692 436704 136698 436716
rect 189810 436704 189816 436716
rect 189868 436704 189874 436756
rect 255406 436704 255412 436756
rect 255464 436744 255470 436756
rect 262306 436744 262312 436756
rect 255464 436716 262312 436744
rect 255464 436704 255470 436716
rect 262306 436704 262312 436716
rect 262364 436704 262370 436756
rect 120718 436500 120724 436552
rect 120776 436540 120782 436552
rect 122098 436540 122104 436552
rect 120776 436512 122104 436540
rect 120776 436500 120782 436512
rect 122098 436500 122104 436512
rect 122156 436500 122162 436552
rect 74074 436432 74080 436484
rect 74132 436472 74138 436484
rect 76558 436472 76564 436484
rect 74132 436444 76564 436472
rect 74132 436432 74138 436444
rect 76558 436432 76564 436444
rect 76616 436432 76622 436484
rect 87322 436296 87328 436348
rect 87380 436336 87386 436348
rect 88242 436336 88248 436348
rect 87380 436308 88248 436336
rect 87380 436296 87386 436308
rect 88242 436296 88248 436308
rect 88300 436296 88306 436348
rect 52178 436092 52184 436144
rect 52236 436132 52242 436144
rect 68922 436132 68928 436144
rect 52236 436104 68928 436132
rect 52236 436092 52242 436104
rect 68922 436092 68928 436104
rect 68980 436092 68986 436144
rect 69658 436092 69664 436144
rect 69716 436132 69722 436144
rect 71038 436132 71044 436144
rect 69716 436104 71044 436132
rect 69716 436092 69722 436104
rect 71038 436092 71044 436104
rect 71096 436092 71102 436144
rect 75822 436092 75828 436144
rect 75880 436132 75886 436144
rect 80422 436132 80428 436144
rect 75880 436104 80428 436132
rect 75880 436092 75886 436104
rect 80422 436092 80428 436104
rect 80480 436092 80486 436144
rect 108298 436092 108304 436144
rect 108356 436132 108362 436144
rect 120718 436132 120724 436144
rect 108356 436104 120724 436132
rect 108356 436092 108362 436104
rect 120718 436092 120724 436104
rect 120776 436092 120782 436144
rect 186958 436024 186964 436076
rect 187016 436064 187022 436076
rect 191558 436064 191564 436076
rect 187016 436036 191564 436064
rect 187016 436024 187022 436036
rect 191558 436024 191564 436036
rect 191616 436024 191622 436076
rect 103882 435412 103888 435464
rect 103940 435452 103946 435464
rect 104434 435452 104440 435464
rect 103940 435424 104440 435452
rect 103940 435412 103946 435424
rect 104434 435412 104440 435424
rect 104492 435452 104498 435464
rect 136634 435452 136640 435464
rect 104492 435424 136640 435452
rect 104492 435412 104498 435424
rect 136634 435412 136640 435424
rect 136692 435412 136698 435464
rect 67266 435344 67272 435396
rect 67324 435384 67330 435396
rect 176654 435384 176660 435396
rect 67324 435356 176660 435384
rect 67324 435344 67330 435356
rect 176654 435344 176660 435356
rect 176712 435344 176718 435396
rect 255406 435344 255412 435396
rect 255464 435384 255470 435396
rect 259638 435384 259644 435396
rect 255464 435356 259644 435384
rect 255464 435344 255470 435356
rect 259638 435344 259644 435356
rect 259696 435384 259702 435396
rect 271874 435384 271880 435396
rect 259696 435356 271880 435384
rect 259696 435344 259702 435356
rect 271874 435344 271880 435356
rect 271932 435344 271938 435396
rect 15838 434732 15844 434784
rect 15896 434772 15902 434784
rect 70578 434772 70584 434784
rect 15896 434744 70584 434772
rect 15896 434732 15902 434744
rect 70578 434732 70584 434744
rect 70636 434732 70642 434784
rect 115750 434664 115756 434716
rect 115808 434704 115814 434716
rect 180150 434704 180156 434716
rect 115808 434676 180156 434704
rect 115808 434664 115814 434676
rect 180150 434664 180156 434676
rect 180208 434664 180214 434716
rect 255406 434664 255412 434716
rect 255464 434704 255470 434716
rect 262214 434704 262220 434716
rect 255464 434676 262220 434704
rect 255464 434664 255470 434676
rect 262214 434664 262220 434676
rect 262272 434704 262278 434716
rect 263686 434704 263692 434716
rect 262272 434676 263692 434704
rect 262272 434664 262278 434676
rect 263686 434664 263692 434676
rect 263744 434664 263750 434716
rect 57606 434052 57612 434104
rect 57664 434092 57670 434104
rect 60642 434092 60648 434104
rect 57664 434064 60648 434092
rect 57664 434052 57670 434064
rect 60642 434052 60648 434064
rect 60700 434092 60706 434104
rect 66806 434092 66812 434104
rect 60700 434064 66812 434092
rect 60700 434052 60706 434064
rect 66806 434052 66812 434064
rect 66864 434052 66870 434104
rect 104158 433984 104164 434036
rect 104216 434024 104222 434036
rect 115290 434024 115296 434036
rect 104216 433996 115296 434024
rect 104216 433984 104222 433996
rect 115290 433984 115296 433996
rect 115348 433984 115354 434036
rect 180702 433984 180708 434036
rect 180760 434024 180766 434036
rect 191098 434024 191104 434036
rect 180760 433996 191104 434024
rect 180760 433984 180766 433996
rect 191098 433984 191104 433996
rect 191156 433984 191162 434036
rect 68370 433644 68376 433696
rect 68428 433684 68434 433696
rect 71130 433684 71136 433696
rect 68428 433656 71136 433684
rect 68428 433644 68434 433656
rect 71130 433644 71136 433656
rect 71188 433644 71194 433696
rect 112346 433644 112352 433696
rect 112404 433684 112410 433696
rect 114002 433684 114008 433696
rect 112404 433656 114008 433684
rect 112404 433644 112410 433656
rect 114002 433644 114008 433656
rect 114060 433644 114066 433696
rect 68646 433236 68652 433288
rect 68704 433276 68710 433288
rect 188430 433276 188436 433288
rect 68704 433248 188436 433276
rect 68704 433236 68710 433248
rect 188430 433236 188436 433248
rect 188488 433236 188494 433288
rect 115842 433168 115848 433220
rect 115900 433208 115906 433220
rect 123478 433208 123484 433220
rect 115900 433180 123484 433208
rect 115900 433168 115906 433180
rect 123478 433168 123484 433180
rect 123536 433168 123542 433220
rect 185578 433168 185584 433220
rect 185636 433208 185642 433220
rect 190638 433208 190644 433220
rect 185636 433180 190644 433208
rect 185636 433168 185642 433180
rect 190638 433168 190644 433180
rect 190696 433168 190702 433220
rect 64598 431944 64604 431996
rect 64656 431984 64662 431996
rect 67542 431984 67548 431996
rect 64656 431956 67548 431984
rect 64656 431944 64662 431956
rect 67542 431944 67548 431956
rect 67600 431944 67606 431996
rect 255406 431944 255412 431996
rect 255464 431984 255470 431996
rect 262214 431984 262220 431996
rect 255464 431956 262220 431984
rect 255464 431944 255470 431956
rect 262214 431944 262220 431956
rect 262272 431944 262278 431996
rect 115842 431196 115848 431248
rect 115900 431236 115906 431248
rect 118694 431236 118700 431248
rect 115900 431208 118700 431236
rect 115900 431196 115906 431208
rect 118694 431196 118700 431208
rect 118752 431196 118758 431248
rect 152458 431196 152464 431248
rect 152516 431236 152522 431248
rect 191190 431236 191196 431248
rect 152516 431208 191196 431236
rect 152516 431196 152522 431208
rect 191190 431196 191196 431208
rect 191248 431196 191254 431248
rect 170398 430516 170404 430568
rect 170456 430556 170462 430568
rect 191098 430556 191104 430568
rect 170456 430528 191104 430556
rect 170456 430516 170462 430528
rect 191098 430516 191104 430528
rect 191156 430516 191162 430568
rect 114002 429836 114008 429888
rect 114060 429876 114066 429888
rect 143626 429876 143632 429888
rect 114060 429848 143632 429876
rect 114060 429836 114066 429848
rect 143626 429836 143632 429848
rect 143684 429836 143690 429888
rect 255498 429496 255504 429548
rect 255556 429536 255562 429548
rect 259546 429536 259552 429548
rect 255556 429508 259552 429536
rect 255556 429496 255562 429508
rect 259546 429496 259552 429508
rect 259604 429496 259610 429548
rect 181438 429088 181444 429140
rect 181496 429128 181502 429140
rect 191742 429128 191748 429140
rect 181496 429100 191748 429128
rect 181496 429088 181502 429100
rect 191742 429088 191748 429100
rect 191800 429088 191806 429140
rect 115842 428408 115848 428460
rect 115900 428448 115906 428460
rect 122834 428448 122840 428460
rect 115900 428420 122840 428448
rect 115900 428408 115906 428420
rect 122834 428408 122840 428420
rect 122892 428448 122898 428460
rect 123018 428448 123024 428460
rect 122892 428420 123024 428448
rect 122892 428408 122898 428420
rect 123018 428408 123024 428420
rect 123076 428408 123082 428460
rect 255406 428408 255412 428460
rect 255464 428448 255470 428460
rect 270586 428448 270592 428460
rect 255464 428420 270592 428448
rect 255464 428408 255470 428420
rect 270586 428408 270592 428420
rect 270644 428408 270650 428460
rect 67542 428340 67548 428392
rect 67600 428380 67606 428392
rect 68278 428380 68284 428392
rect 67600 428352 68284 428380
rect 67600 428340 67606 428352
rect 68278 428340 68284 428352
rect 68336 428340 68342 428392
rect 255406 427796 255412 427848
rect 255464 427836 255470 427848
rect 288434 427836 288440 427848
rect 255464 427808 288440 427836
rect 255464 427796 255470 427808
rect 288434 427796 288440 427808
rect 288492 427796 288498 427848
rect 255498 427728 255504 427780
rect 255556 427768 255562 427780
rect 260834 427768 260840 427780
rect 255556 427740 260840 427768
rect 255556 427728 255562 427740
rect 260834 427728 260840 427740
rect 260892 427768 260898 427780
rect 262122 427768 262128 427780
rect 260892 427740 262128 427768
rect 260892 427728 260898 427740
rect 262122 427728 262128 427740
rect 262180 427728 262186 427780
rect 116578 427048 116584 427100
rect 116636 427088 116642 427100
rect 162118 427088 162124 427100
rect 116636 427060 162124 427088
rect 116636 427048 116642 427060
rect 162118 427048 162124 427060
rect 162176 427048 162182 427100
rect 262122 427048 262128 427100
rect 262180 427088 262186 427100
rect 285674 427088 285680 427100
rect 262180 427060 285680 427088
rect 262180 427048 262186 427060
rect 285674 427048 285680 427060
rect 285732 427048 285738 427100
rect 63402 426436 63408 426488
rect 63460 426476 63466 426488
rect 66990 426476 66996 426488
rect 63460 426448 66996 426476
rect 63460 426436 63466 426448
rect 66990 426436 66996 426448
rect 67048 426436 67054 426488
rect 190638 426476 190644 426488
rect 171106 426448 190644 426476
rect 151078 426368 151084 426420
rect 151136 426408 151142 426420
rect 170398 426408 170404 426420
rect 151136 426380 170404 426408
rect 151136 426368 151142 426380
rect 170398 426368 170404 426380
rect 170456 426408 170462 426420
rect 171106 426408 171134 426448
rect 190638 426436 190644 426448
rect 190696 426436 190702 426488
rect 285674 426436 285680 426488
rect 285732 426476 285738 426488
rect 582650 426476 582656 426488
rect 285732 426448 582656 426476
rect 285732 426436 285738 426448
rect 582650 426436 582656 426448
rect 582708 426436 582714 426488
rect 170456 426380 171134 426408
rect 170456 426368 170462 426380
rect 115382 426232 115388 426284
rect 115440 426272 115446 426284
rect 119338 426272 119344 426284
rect 115440 426244 119344 426272
rect 115440 426232 115446 426244
rect 119338 426232 119344 426244
rect 119396 426232 119402 426284
rect 57790 425688 57796 425740
rect 57848 425728 57854 425740
rect 67266 425728 67272 425740
rect 57848 425700 67272 425728
rect 57848 425688 57854 425700
rect 67266 425688 67272 425700
rect 67324 425688 67330 425740
rect 126330 425688 126336 425740
rect 126388 425728 126394 425740
rect 141418 425728 141424 425740
rect 126388 425700 141424 425728
rect 126388 425688 126394 425700
rect 141418 425688 141424 425700
rect 141476 425688 141482 425740
rect 174538 425688 174544 425740
rect 174596 425728 174602 425740
rect 191742 425728 191748 425740
rect 174596 425700 191748 425728
rect 174596 425688 174602 425700
rect 191742 425688 191748 425700
rect 191800 425688 191806 425740
rect 255866 425688 255872 425740
rect 255924 425728 255930 425740
rect 256786 425728 256792 425740
rect 255924 425700 256792 425728
rect 255924 425688 255930 425700
rect 256786 425688 256792 425700
rect 256844 425728 256850 425740
rect 269206 425728 269212 425740
rect 256844 425700 269212 425728
rect 256844 425688 256850 425700
rect 269206 425688 269212 425700
rect 269264 425688 269270 425740
rect 115014 425008 115020 425060
rect 115072 425048 115078 425060
rect 117498 425048 117504 425060
rect 115072 425020 117504 425048
rect 115072 425008 115078 425020
rect 117498 425008 117504 425020
rect 117556 425008 117562 425060
rect 115382 424940 115388 424992
rect 115440 424980 115446 424992
rect 117406 424980 117412 424992
rect 115440 424952 117412 424980
rect 115440 424940 115446 424952
rect 117406 424940 117412 424952
rect 117464 424940 117470 424992
rect 54938 423648 54944 423700
rect 54996 423688 55002 423700
rect 66622 423688 66628 423700
rect 54996 423660 66628 423688
rect 54996 423648 55002 423660
rect 66622 423648 66628 423660
rect 66680 423648 66686 423700
rect 115014 423512 115020 423564
rect 115072 423552 115078 423564
rect 120810 423552 120816 423564
rect 115072 423524 120816 423552
rect 115072 423512 115078 423524
rect 120810 423512 120816 423524
rect 120868 423512 120874 423564
rect 49602 422900 49608 422952
rect 49660 422940 49666 422952
rect 64782 422940 64788 422952
rect 49660 422912 64788 422940
rect 49660 422900 49666 422912
rect 64782 422900 64788 422912
rect 64840 422940 64846 422952
rect 66806 422940 66812 422952
rect 64840 422912 66812 422940
rect 64840 422900 64846 422912
rect 66806 422900 66812 422912
rect 66864 422900 66870 422952
rect 126238 422900 126244 422952
rect 126296 422940 126302 422952
rect 166258 422940 166264 422952
rect 126296 422912 166264 422940
rect 126296 422900 126302 422912
rect 166258 422900 166264 422912
rect 166316 422900 166322 422952
rect 166258 422288 166264 422340
rect 166316 422328 166322 422340
rect 190638 422328 190644 422340
rect 166316 422300 190644 422328
rect 166316 422288 166322 422300
rect 190638 422288 190644 422300
rect 190696 422288 190702 422340
rect 255498 422288 255504 422340
rect 255556 422328 255562 422340
rect 276106 422328 276112 422340
rect 255556 422300 276112 422328
rect 255556 422288 255562 422300
rect 276106 422288 276112 422300
rect 276164 422288 276170 422340
rect 62022 422220 62028 422272
rect 62080 422260 62086 422272
rect 66622 422260 66628 422272
rect 62080 422232 66628 422260
rect 62080 422220 62086 422232
rect 66622 422220 66628 422232
rect 66680 422220 66686 422272
rect 52270 421540 52276 421592
rect 52328 421580 52334 421592
rect 62022 421580 62028 421592
rect 52328 421552 62028 421580
rect 52328 421540 52334 421552
rect 62022 421540 62028 421552
rect 62080 421540 62086 421592
rect 255958 421540 255964 421592
rect 256016 421580 256022 421592
rect 262858 421580 262864 421592
rect 256016 421552 262864 421580
rect 256016 421540 256022 421552
rect 262858 421540 262864 421552
rect 262916 421540 262922 421592
rect 115290 420928 115296 420980
rect 115348 420968 115354 420980
rect 188430 420968 188436 420980
rect 115348 420940 188436 420968
rect 115348 420928 115354 420940
rect 188430 420928 188436 420940
rect 188488 420928 188494 420980
rect 255498 420928 255504 420980
rect 255556 420968 255562 420980
rect 283006 420968 283012 420980
rect 255556 420940 283012 420968
rect 255556 420928 255562 420940
rect 283006 420928 283012 420940
rect 283064 420928 283070 420980
rect 60458 420860 60464 420912
rect 60516 420900 60522 420912
rect 66806 420900 66812 420912
rect 60516 420872 66812 420900
rect 60516 420860 60522 420872
rect 66806 420860 66812 420872
rect 66864 420860 66870 420912
rect 64782 420248 64788 420300
rect 64840 420288 64846 420300
rect 67082 420288 67088 420300
rect 64840 420260 67088 420288
rect 64840 420248 64846 420260
rect 67082 420248 67088 420260
rect 67140 420248 67146 420300
rect 115750 419500 115756 419552
rect 115808 419540 115814 419552
rect 129826 419540 129832 419552
rect 115808 419512 129832 419540
rect 115808 419500 115814 419512
rect 129826 419500 129832 419512
rect 129884 419500 129890 419552
rect 171870 419500 171876 419552
rect 171928 419540 171934 419552
rect 191742 419540 191748 419552
rect 171928 419512 191748 419540
rect 171928 419500 171934 419512
rect 191742 419500 191748 419512
rect 191800 419500 191806 419552
rect 255498 419500 255504 419552
rect 255556 419540 255562 419552
rect 260834 419540 260840 419552
rect 255556 419512 260840 419540
rect 255556 419500 255562 419512
rect 260834 419500 260840 419512
rect 260892 419500 260898 419552
rect 59262 418752 59268 418804
rect 59320 418792 59326 418804
rect 67634 418792 67640 418804
rect 59320 418764 67640 418792
rect 59320 418752 59326 418764
rect 67634 418752 67640 418764
rect 67692 418752 67698 418804
rect 123478 418752 123484 418804
rect 123536 418792 123542 418804
rect 136726 418792 136732 418804
rect 123536 418764 136732 418792
rect 123536 418752 123542 418764
rect 136726 418752 136732 418764
rect 136784 418792 136790 418804
rect 187050 418792 187056 418804
rect 136784 418764 187056 418792
rect 136784 418752 136790 418764
rect 187050 418752 187056 418764
rect 187108 418752 187114 418804
rect 289722 418752 289728 418804
rect 289780 418792 289786 418804
rect 583110 418792 583116 418804
rect 289780 418764 583116 418792
rect 289780 418752 289786 418764
rect 583110 418752 583116 418764
rect 583168 418752 583174 418804
rect 59170 418276 59176 418328
rect 59228 418316 59234 418328
rect 66806 418316 66812 418328
rect 59228 418288 66812 418316
rect 59228 418276 59234 418288
rect 66806 418276 66812 418288
rect 66864 418276 66870 418328
rect 178678 418140 178684 418192
rect 178736 418180 178742 418192
rect 191742 418180 191748 418192
rect 178736 418152 191748 418180
rect 178736 418140 178742 418152
rect 191742 418140 191748 418152
rect 191800 418140 191806 418192
rect 255406 418140 255412 418192
rect 255464 418180 255470 418192
rect 288618 418180 288624 418192
rect 255464 418152 288624 418180
rect 255464 418140 255470 418152
rect 288618 418140 288624 418152
rect 288676 418180 288682 418192
rect 289722 418180 289728 418192
rect 288676 418152 289728 418180
rect 288676 418140 288682 418152
rect 289722 418140 289728 418152
rect 289780 418140 289786 418192
rect 64690 418072 64696 418124
rect 64748 418112 64754 418124
rect 67082 418112 67088 418124
rect 64748 418084 67088 418112
rect 64748 418072 64754 418084
rect 67082 418072 67088 418084
rect 67140 418072 67146 418124
rect 112714 418072 112720 418124
rect 112772 418112 112778 418124
rect 170490 418112 170496 418124
rect 112772 418084 170496 418112
rect 112772 418072 112778 418084
rect 170490 418072 170496 418084
rect 170548 418072 170554 418124
rect 265250 417460 265256 417512
rect 265308 417500 265314 417512
rect 271138 417500 271144 417512
rect 265308 417472 271144 417500
rect 265308 417460 265314 417472
rect 271138 417460 271144 417472
rect 271196 417460 271202 417512
rect 162118 417392 162124 417444
rect 162176 417432 162182 417444
rect 162762 417432 162768 417444
rect 162176 417404 162768 417432
rect 162176 417392 162182 417404
rect 162762 417392 162768 417404
rect 162820 417432 162826 417444
rect 191742 417432 191748 417444
rect 162820 417404 191748 417432
rect 162820 417392 162826 417404
rect 191742 417392 191748 417404
rect 191800 417392 191806 417444
rect 270402 417392 270408 417444
rect 270460 417432 270466 417444
rect 583202 417432 583208 417444
rect 270460 417404 583208 417432
rect 270460 417392 270466 417404
rect 583202 417392 583208 417404
rect 583260 417392 583266 417444
rect 113910 417052 113916 417104
rect 113968 417092 113974 417104
rect 117958 417092 117964 417104
rect 113968 417064 117964 417092
rect 113968 417052 113974 417064
rect 117958 417052 117964 417064
rect 118016 417052 118022 417104
rect 255406 416848 255412 416900
rect 255464 416888 255470 416900
rect 265066 416888 265072 416900
rect 255464 416860 265072 416888
rect 255464 416848 255470 416860
rect 265066 416848 265072 416860
rect 265124 416888 265130 416900
rect 265250 416888 265256 416900
rect 265124 416860 265256 416888
rect 265124 416848 265130 416860
rect 265250 416848 265256 416860
rect 265308 416848 265314 416900
rect 255498 416780 255504 416832
rect 255556 416820 255562 416832
rect 269298 416820 269304 416832
rect 255556 416792 269304 416820
rect 255556 416780 255562 416792
rect 269298 416780 269304 416792
rect 269356 416820 269362 416832
rect 270402 416820 270408 416832
rect 269356 416792 270408 416820
rect 269356 416780 269362 416792
rect 270402 416780 270408 416792
rect 270460 416780 270466 416832
rect 63310 416712 63316 416764
rect 63368 416752 63374 416764
rect 66254 416752 66260 416764
rect 63368 416724 66260 416752
rect 63368 416712 63374 416724
rect 66254 416712 66260 416724
rect 66312 416712 66318 416764
rect 116118 416100 116124 416152
rect 116176 416140 116182 416152
rect 126330 416140 126336 416152
rect 116176 416112 126336 416140
rect 116176 416100 116182 416112
rect 126330 416100 126336 416112
rect 126388 416100 126394 416152
rect 116578 416032 116584 416084
rect 116636 416072 116642 416084
rect 142154 416072 142160 416084
rect 116636 416044 142160 416072
rect 116636 416032 116642 416044
rect 142154 416032 142160 416044
rect 142212 416072 142218 416084
rect 173158 416072 173164 416084
rect 142212 416044 173164 416072
rect 142212 416032 142218 416044
rect 173158 416032 173164 416044
rect 173216 416032 173222 416084
rect 187694 415896 187700 415948
rect 187752 415936 187758 415948
rect 188982 415936 188988 415948
rect 187752 415908 188988 415936
rect 187752 415896 187758 415908
rect 188982 415896 188988 415908
rect 189040 415936 189046 415948
rect 190638 415936 190644 415948
rect 189040 415908 190644 415936
rect 189040 415896 189046 415908
rect 190638 415896 190644 415908
rect 190696 415896 190702 415948
rect 63218 415012 63224 415064
rect 63276 415052 63282 415064
rect 66898 415052 66904 415064
rect 63276 415024 66904 415052
rect 63276 415012 63282 415024
rect 66898 415012 66904 415024
rect 66956 415012 66962 415064
rect 115842 414672 115848 414724
rect 115900 414712 115906 414724
rect 125686 414712 125692 414724
rect 115900 414684 125692 414712
rect 115900 414672 115906 414684
rect 125686 414672 125692 414684
rect 125744 414672 125750 414724
rect 53650 413992 53656 414044
rect 53708 414032 53714 414044
rect 66806 414032 66812 414044
rect 53708 414004 66812 414032
rect 53708 413992 53714 414004
rect 66806 413992 66812 414004
rect 66864 413992 66870 414044
rect 142154 413992 142160 414044
rect 142212 414032 142218 414044
rect 191742 414032 191748 414044
rect 142212 414004 191748 414032
rect 142212 413992 142218 414004
rect 191742 413992 191748 414004
rect 191800 413992 191806 414044
rect 255406 413516 255412 413568
rect 255464 413556 255470 413568
rect 258166 413556 258172 413568
rect 255464 413528 258172 413556
rect 255464 413516 255470 413528
rect 258166 413516 258172 413528
rect 258224 413516 258230 413568
rect 113174 412972 113180 413024
rect 113232 413012 113238 413024
rect 117314 413012 117320 413024
rect 113232 412984 117320 413012
rect 113232 412972 113238 412984
rect 117314 412972 117320 412984
rect 117372 412972 117378 413024
rect 46842 412632 46848 412684
rect 46900 412672 46906 412684
rect 66254 412672 66260 412684
rect 46900 412644 66260 412672
rect 46900 412632 46906 412644
rect 66254 412632 66260 412644
rect 66312 412632 66318 412684
rect 121638 412632 121644 412684
rect 121696 412672 121702 412684
rect 148318 412672 148324 412684
rect 121696 412644 148324 412672
rect 121696 412632 121702 412644
rect 148318 412632 148324 412644
rect 148376 412632 148382 412684
rect 115842 412564 115848 412616
rect 115900 412604 115906 412616
rect 123478 412604 123484 412616
rect 115900 412576 123484 412604
rect 115900 412564 115906 412576
rect 123478 412564 123484 412576
rect 123536 412564 123542 412616
rect 166350 411884 166356 411936
rect 166408 411924 166414 411936
rect 166902 411924 166908 411936
rect 166408 411896 166908 411924
rect 166408 411884 166414 411896
rect 166902 411884 166908 411896
rect 166960 411924 166966 411936
rect 191742 411924 191748 411936
rect 166960 411896 191748 411924
rect 166960 411884 166966 411896
rect 191742 411884 191748 411896
rect 191800 411884 191806 411936
rect 39942 411272 39948 411324
rect 40000 411312 40006 411324
rect 66254 411312 66260 411324
rect 40000 411284 66260 411312
rect 40000 411272 40006 411284
rect 66254 411272 66260 411284
rect 66312 411272 66318 411324
rect 50798 411204 50804 411256
rect 50856 411244 50862 411256
rect 57698 411244 57704 411256
rect 50856 411216 57704 411244
rect 50856 411204 50862 411216
rect 57698 411204 57704 411216
rect 57756 411244 57762 411256
rect 66622 411244 66628 411256
rect 57756 411216 66628 411244
rect 57756 411204 57762 411216
rect 66622 411204 66628 411216
rect 66680 411204 66686 411256
rect 114738 410592 114744 410644
rect 114796 410632 114802 410644
rect 116578 410632 116584 410644
rect 114796 410604 116584 410632
rect 114796 410592 114802 410604
rect 116578 410592 116584 410604
rect 116636 410592 116642 410644
rect 118694 410524 118700 410576
rect 118752 410564 118758 410576
rect 131114 410564 131120 410576
rect 118752 410536 131120 410564
rect 118752 410524 118758 410536
rect 131114 410524 131120 410536
rect 131172 410564 131178 410576
rect 180150 410564 180156 410576
rect 131172 410536 180156 410564
rect 131172 410524 131178 410536
rect 180150 410524 180156 410536
rect 180208 410524 180214 410576
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 7650 409884 7656 409896
rect 3200 409856 7656 409884
rect 3200 409844 3206 409856
rect 7650 409844 7656 409856
rect 7708 409844 7714 409896
rect 188890 409844 188896 409896
rect 188948 409884 188954 409896
rect 191006 409884 191012 409896
rect 188948 409856 191012 409884
rect 188948 409844 188954 409856
rect 191006 409844 191012 409856
rect 191064 409844 191070 409896
rect 255406 409844 255412 409896
rect 255464 409884 255470 409896
rect 266446 409884 266452 409896
rect 255464 409856 266452 409884
rect 255464 409844 255470 409856
rect 266446 409844 266452 409856
rect 266504 409844 266510 409896
rect 125502 409096 125508 409148
rect 125560 409136 125566 409148
rect 143534 409136 143540 409148
rect 125560 409108 143540 409136
rect 125560 409096 125566 409108
rect 143534 409096 143540 409108
rect 143592 409136 143598 409148
rect 187142 409136 187148 409148
rect 143592 409108 187148 409136
rect 143592 409096 143598 409108
rect 187142 409096 187148 409108
rect 187200 409096 187206 409148
rect 62758 408524 62764 408536
rect 62224 408496 62764 408524
rect 59078 408416 59084 408468
rect 59136 408456 59142 408468
rect 62224 408456 62252 408496
rect 62758 408484 62764 408496
rect 62816 408524 62822 408536
rect 66806 408524 66812 408536
rect 62816 408496 66812 408524
rect 62816 408484 62822 408496
rect 66806 408484 66812 408496
rect 66864 408484 66870 408536
rect 115842 408484 115848 408536
rect 115900 408524 115906 408536
rect 152458 408524 152464 408536
rect 115900 408496 152464 408524
rect 115900 408484 115906 408496
rect 152458 408484 152464 408496
rect 152516 408484 152522 408536
rect 186222 408484 186228 408536
rect 186280 408524 186286 408536
rect 191006 408524 191012 408536
rect 186280 408496 191012 408524
rect 186280 408484 186286 408496
rect 191006 408484 191012 408496
rect 191064 408484 191070 408536
rect 255406 408484 255412 408536
rect 255464 408524 255470 408536
rect 273346 408524 273352 408536
rect 255464 408496 273352 408524
rect 255464 408484 255470 408496
rect 273346 408484 273352 408496
rect 273404 408484 273410 408536
rect 59136 408428 62252 408456
rect 59136 408416 59142 408428
rect 130378 408416 130384 408468
rect 130436 408456 130442 408468
rect 142154 408456 142160 408468
rect 130436 408428 142160 408456
rect 130436 408416 130442 408428
rect 142154 408416 142160 408428
rect 142212 408416 142218 408468
rect 115382 408348 115388 408400
rect 115440 408388 115446 408400
rect 121638 408388 121644 408400
rect 115440 408360 121644 408388
rect 115440 408348 115446 408360
rect 121638 408348 121644 408360
rect 121696 408348 121702 408400
rect 48130 407124 48136 407176
rect 48188 407164 48194 407176
rect 66898 407164 66904 407176
rect 48188 407136 66904 407164
rect 48188 407124 48194 407136
rect 66898 407124 66904 407136
rect 66956 407124 66962 407176
rect 53834 407056 53840 407108
rect 53892 407096 53898 407108
rect 55030 407096 55036 407108
rect 53892 407068 55036 407096
rect 53892 407056 53898 407068
rect 55030 407056 55036 407068
rect 55088 407096 55094 407108
rect 66806 407096 66812 407108
rect 55088 407068 66812 407096
rect 55088 407056 55094 407068
rect 66806 407056 66812 407068
rect 66864 407056 66870 407108
rect 254578 407056 254584 407108
rect 254636 407096 254642 407108
rect 259546 407096 259552 407108
rect 254636 407068 259552 407096
rect 254636 407056 254642 407068
rect 259546 407056 259552 407068
rect 259604 407056 259610 407108
rect 41230 406376 41236 406428
rect 41288 406416 41294 406428
rect 53834 406416 53840 406428
rect 41288 406388 53840 406416
rect 41288 406376 41294 406388
rect 53834 406376 53840 406388
rect 53892 406376 53898 406428
rect 255406 406240 255412 406292
rect 255464 406280 255470 406292
rect 259638 406280 259644 406292
rect 255464 406252 259644 406280
rect 255464 406240 255470 406252
rect 259638 406240 259644 406252
rect 259696 406240 259702 406292
rect 159358 405696 159364 405748
rect 159416 405736 159422 405748
rect 191742 405736 191748 405748
rect 159416 405708 191748 405736
rect 159416 405696 159422 405708
rect 191742 405696 191748 405708
rect 191800 405696 191806 405748
rect 115842 405628 115848 405680
rect 115900 405668 115906 405680
rect 125502 405668 125508 405680
rect 115900 405640 125508 405668
rect 115900 405628 115906 405640
rect 125502 405628 125508 405640
rect 125560 405628 125566 405680
rect 115750 405560 115756 405612
rect 115808 405600 115814 405612
rect 118694 405600 118700 405612
rect 115808 405572 118700 405600
rect 115808 405560 115814 405572
rect 118694 405560 118700 405572
rect 118752 405560 118758 405612
rect 64690 404336 64696 404388
rect 64748 404376 64754 404388
rect 66806 404376 66812 404388
rect 64748 404348 66812 404376
rect 64748 404336 64754 404348
rect 66806 404336 66812 404348
rect 66864 404336 66870 404388
rect 162118 404336 162124 404388
rect 162176 404376 162182 404388
rect 191742 404376 191748 404388
rect 162176 404348 191748 404376
rect 162176 404336 162182 404348
rect 191742 404336 191748 404348
rect 191800 404336 191806 404388
rect 147674 403724 147680 403776
rect 147732 403764 147738 403776
rect 148410 403764 148416 403776
rect 147732 403736 148416 403764
rect 147732 403724 147738 403736
rect 148410 403724 148416 403736
rect 148468 403724 148474 403776
rect 117222 403044 117228 403096
rect 117280 403084 117286 403096
rect 147674 403084 147680 403096
rect 117280 403056 147680 403084
rect 117280 403044 117286 403056
rect 147674 403044 147680 403056
rect 147732 403044 147738 403096
rect 55030 402976 55036 403028
rect 55088 403016 55094 403028
rect 66806 403016 66812 403028
rect 55088 402988 66812 403016
rect 55088 402976 55094 402988
rect 66806 402976 66812 402988
rect 66864 402976 66870 403028
rect 115842 402976 115848 403028
rect 115900 403016 115906 403028
rect 155218 403016 155224 403028
rect 115900 402988 155224 403016
rect 115900 402976 115906 402988
rect 155218 402976 155224 402988
rect 155276 402976 155282 403028
rect 156598 402976 156604 403028
rect 156656 403016 156662 403028
rect 191742 403016 191748 403028
rect 156656 402988 191748 403016
rect 156656 402976 156662 402988
rect 191742 402976 191748 402988
rect 191800 402976 191806 403028
rect 113450 402364 113456 402416
rect 113508 402404 113514 402416
rect 118786 402404 118792 402416
rect 113508 402376 118792 402404
rect 113508 402364 113514 402376
rect 118786 402364 118792 402376
rect 118844 402364 118850 402416
rect 64598 401616 64604 401668
rect 64656 401656 64662 401668
rect 66254 401656 66260 401668
rect 64656 401628 66260 401656
rect 64656 401616 64662 401628
rect 66254 401616 66260 401628
rect 66312 401616 66318 401668
rect 114738 401072 114744 401124
rect 114796 401112 114802 401124
rect 117222 401112 117228 401124
rect 114796 401084 117228 401112
rect 114796 401072 114802 401084
rect 117222 401072 117228 401084
rect 117280 401072 117286 401124
rect 121638 400868 121644 400920
rect 121696 400908 121702 400920
rect 128354 400908 128360 400920
rect 121696 400880 128360 400908
rect 121696 400868 121702 400880
rect 128354 400868 128360 400880
rect 128412 400868 128418 400920
rect 60642 400188 60648 400240
rect 60700 400228 60706 400240
rect 66714 400228 66720 400240
rect 60700 400200 66720 400228
rect 60700 400188 60706 400200
rect 66714 400188 66720 400200
rect 66772 400188 66778 400240
rect 115566 400188 115572 400240
rect 115624 400228 115630 400240
rect 119338 400228 119344 400240
rect 115624 400200 119344 400228
rect 115624 400188 115630 400200
rect 119338 400188 119344 400200
rect 119396 400188 119402 400240
rect 255406 400188 255412 400240
rect 255464 400228 255470 400240
rect 277486 400228 277492 400240
rect 255464 400200 277492 400228
rect 255464 400188 255470 400200
rect 277486 400188 277492 400200
rect 277544 400188 277550 400240
rect 255406 399440 255412 399492
rect 255464 399480 255470 399492
rect 258258 399480 258264 399492
rect 255464 399452 258264 399480
rect 255464 399440 255470 399452
rect 258258 399440 258264 399452
rect 258316 399480 258322 399492
rect 582834 399480 582840 399492
rect 258316 399452 582840 399480
rect 258316 399440 258322 399452
rect 582834 399440 582840 399452
rect 582892 399440 582898 399492
rect 192662 398936 192668 398948
rect 180766 398908 192668 398936
rect 115842 398828 115848 398880
rect 115900 398868 115906 398880
rect 180766 398868 180794 398908
rect 192662 398896 192668 398908
rect 192720 398896 192726 398948
rect 115900 398840 180794 398868
rect 115900 398828 115906 398840
rect 184290 398828 184296 398880
rect 184348 398868 184354 398880
rect 191742 398868 191748 398880
rect 184348 398840 191748 398868
rect 184348 398828 184354 398840
rect 191742 398828 191748 398840
rect 191800 398828 191806 398880
rect 4798 397468 4804 397520
rect 4856 397508 4862 397520
rect 63310 397508 63316 397520
rect 4856 397480 63316 397508
rect 4856 397468 4862 397480
rect 63310 397468 63316 397480
rect 63368 397508 63374 397520
rect 67174 397508 67180 397520
rect 63368 397480 67180 397508
rect 63368 397468 63374 397480
rect 67174 397468 67180 397480
rect 67232 397468 67238 397520
rect 115382 397468 115388 397520
rect 115440 397508 115446 397520
rect 118602 397508 118608 397520
rect 115440 397480 118608 397508
rect 115440 397468 115446 397480
rect 118602 397468 118608 397480
rect 118660 397508 118666 397520
rect 121638 397508 121644 397520
rect 118660 397480 121644 397508
rect 118660 397468 118666 397480
rect 121638 397468 121644 397480
rect 121696 397468 121702 397520
rect 159542 397468 159548 397520
rect 159600 397508 159606 397520
rect 190822 397508 190828 397520
rect 159600 397480 190828 397508
rect 159600 397468 159606 397480
rect 190822 397468 190828 397480
rect 190880 397468 190886 397520
rect 115290 397128 115296 397180
rect 115348 397168 115354 397180
rect 119430 397168 119436 397180
rect 115348 397140 119436 397168
rect 115348 397128 115354 397140
rect 119430 397128 119436 397140
rect 119488 397128 119494 397180
rect 53374 396720 53380 396772
rect 53432 396760 53438 396772
rect 66806 396760 66812 396772
rect 53432 396732 66812 396760
rect 53432 396720 53438 396732
rect 66806 396720 66812 396732
rect 66864 396720 66870 396772
rect 160738 396720 160744 396772
rect 160796 396760 160802 396772
rect 184842 396760 184848 396772
rect 160796 396732 184848 396760
rect 160796 396720 160802 396732
rect 184842 396720 184848 396732
rect 184900 396760 184906 396772
rect 191742 396760 191748 396772
rect 184900 396732 191748 396760
rect 184900 396720 184906 396732
rect 191742 396720 191748 396732
rect 191800 396720 191806 396772
rect 50890 395972 50896 396024
rect 50948 396012 50954 396024
rect 67174 396012 67180 396024
rect 50948 395984 67180 396012
rect 50948 395972 50954 395984
rect 67174 395972 67180 395984
rect 67232 395972 67238 396024
rect 271230 395292 271236 395344
rect 271288 395332 271294 395344
rect 287238 395332 287244 395344
rect 271288 395304 287244 395332
rect 271288 395292 271294 395304
rect 287238 395292 287244 395304
rect 287296 395292 287302 395344
rect 157978 394748 157984 394800
rect 158036 394788 158042 394800
rect 190822 394788 190828 394800
rect 158036 394760 190828 394788
rect 158036 394748 158042 394760
rect 190822 394748 190828 394760
rect 190880 394748 190886 394800
rect 115842 394680 115848 394732
rect 115900 394720 115906 394732
rect 189810 394720 189816 394732
rect 115900 394692 189816 394720
rect 115900 394680 115906 394692
rect 189810 394680 189816 394692
rect 189868 394680 189874 394732
rect 61838 393388 61844 393440
rect 61896 393428 61902 393440
rect 67634 393428 67640 393440
rect 61896 393400 67640 393428
rect 61896 393388 61902 393400
rect 67634 393388 67640 393400
rect 67692 393388 67698 393440
rect 131758 393388 131764 393440
rect 131816 393428 131822 393440
rect 132586 393428 132592 393440
rect 131816 393400 132592 393428
rect 131816 393388 131822 393400
rect 132586 393388 132592 393400
rect 132644 393388 132650 393440
rect 115750 393320 115756 393372
rect 115808 393360 115814 393372
rect 151170 393360 151176 393372
rect 115808 393332 151176 393360
rect 115808 393320 115814 393332
rect 151170 393320 151176 393332
rect 151228 393320 151234 393372
rect 188522 393320 188528 393372
rect 188580 393360 188586 393372
rect 190822 393360 190828 393372
rect 188580 393332 190828 393360
rect 188580 393320 188586 393332
rect 190822 393320 190828 393332
rect 190880 393320 190886 393372
rect 256878 393320 256884 393372
rect 256936 393360 256942 393372
rect 271966 393360 271972 393372
rect 256936 393332 271972 393360
rect 256936 393320 256942 393332
rect 271966 393320 271972 393332
rect 272024 393320 272030 393372
rect 67358 393252 67364 393304
rect 67416 393292 67422 393304
rect 67634 393292 67640 393304
rect 67416 393264 67640 393292
rect 67416 393252 67422 393264
rect 67634 393252 67640 393264
rect 67692 393252 67698 393304
rect 115566 392028 115572 392080
rect 115624 392068 115630 392080
rect 116026 392068 116032 392080
rect 115624 392040 116032 392068
rect 115624 392028 115630 392040
rect 116026 392028 116032 392040
rect 116084 392068 116090 392080
rect 131758 392068 131764 392080
rect 116084 392040 131764 392068
rect 116084 392028 116090 392040
rect 131758 392028 131764 392040
rect 131816 392028 131822 392080
rect 184382 392028 184388 392080
rect 184440 392068 184446 392080
rect 191558 392068 191564 392080
rect 184440 392040 191564 392068
rect 184440 392028 184446 392040
rect 191558 392028 191564 392040
rect 191616 392028 191622 392080
rect 56410 391960 56416 392012
rect 56468 392000 56474 392012
rect 66806 392000 66812 392012
rect 56468 391972 66812 392000
rect 56468 391960 56474 391972
rect 66806 391960 66812 391972
rect 66864 391960 66870 392012
rect 115750 391960 115756 392012
rect 115808 392000 115814 392012
rect 193398 392000 193404 392012
rect 115808 391972 193404 392000
rect 115808 391960 115814 391972
rect 193398 391960 193404 391972
rect 193456 391960 193462 392012
rect 266998 391212 267004 391264
rect 267056 391252 267062 391264
rect 273438 391252 273444 391264
rect 267056 391224 273444 391252
rect 267056 391212 267062 391224
rect 273438 391212 273444 391224
rect 273496 391212 273502 391264
rect 114830 390736 114836 390788
rect 114888 390776 114894 390788
rect 116578 390776 116584 390788
rect 114888 390748 116584 390776
rect 114888 390736 114894 390748
rect 116578 390736 116584 390748
rect 116636 390736 116642 390788
rect 111978 390640 111984 390652
rect 68664 390612 111984 390640
rect 68664 390584 68692 390612
rect 111978 390600 111984 390612
rect 112036 390600 112042 390652
rect 117222 390600 117228 390652
rect 117280 390640 117286 390652
rect 196894 390640 196900 390652
rect 117280 390612 196900 390640
rect 117280 390600 117286 390612
rect 67726 390532 67732 390584
rect 67784 390572 67790 390584
rect 68646 390572 68652 390584
rect 67784 390544 68652 390572
rect 67784 390532 67790 390544
rect 68646 390532 68652 390544
rect 68704 390532 68710 390584
rect 73706 390532 73712 390584
rect 73764 390572 73770 390584
rect 178034 390572 178040 390584
rect 73764 390544 178040 390572
rect 73764 390532 73770 390544
rect 178034 390532 178040 390544
rect 178092 390532 178098 390584
rect 196084 390312 196112 390612
rect 196894 390600 196900 390612
rect 196952 390600 196958 390652
rect 196066 390260 196072 390312
rect 196124 390260 196130 390312
rect 247678 389784 247684 389836
rect 247736 389824 247742 389836
rect 254026 389824 254032 389836
rect 247736 389796 254032 389824
rect 247736 389784 247742 389796
rect 254026 389784 254032 389796
rect 254084 389784 254090 389836
rect 109402 389240 109408 389292
rect 109460 389280 109466 389292
rect 165614 389280 165620 389292
rect 109460 389252 165620 389280
rect 109460 389240 109466 389252
rect 165614 389240 165620 389252
rect 165672 389280 165678 389292
rect 248322 389280 248328 389292
rect 165672 389252 248328 389280
rect 165672 389240 165678 389252
rect 248322 389240 248328 389252
rect 248380 389240 248386 389292
rect 53742 389172 53748 389224
rect 53800 389212 53806 389224
rect 82998 389212 83004 389224
rect 53800 389184 83004 389212
rect 53800 389172 53806 389184
rect 82998 389172 83004 389184
rect 83056 389172 83062 389224
rect 103146 389172 103152 389224
rect 103204 389212 103210 389224
rect 238754 389212 238760 389224
rect 103204 389184 238760 389212
rect 103204 389172 103210 389184
rect 238754 389172 238760 389184
rect 238812 389212 238818 389224
rect 239950 389212 239956 389224
rect 238812 389184 239956 389212
rect 238812 389172 238818 389184
rect 239950 389172 239956 389184
rect 240008 389172 240014 389224
rect 249150 389172 249156 389224
rect 249208 389212 249214 389224
rect 254210 389212 254216 389224
rect 249208 389184 254216 389212
rect 249208 389172 249214 389184
rect 254210 389172 254216 389184
rect 254268 389172 254274 389224
rect 11698 389104 11704 389156
rect 11756 389144 11762 389156
rect 51442 389144 51448 389156
rect 11756 389116 51448 389144
rect 11756 389104 11762 389116
rect 51442 389104 51448 389116
rect 51500 389144 51506 389156
rect 52362 389144 52368 389156
rect 51500 389116 52368 389144
rect 51500 389104 51506 389116
rect 52362 389104 52368 389116
rect 52420 389104 52426 389156
rect 69658 389104 69664 389156
rect 69716 389144 69722 389156
rect 73706 389144 73712 389156
rect 69716 389116 73712 389144
rect 69716 389104 69722 389116
rect 73706 389104 73712 389116
rect 73764 389104 73770 389156
rect 107838 389104 107844 389156
rect 107896 389144 107902 389156
rect 246390 389144 246396 389156
rect 107896 389116 246396 389144
rect 107896 389104 107902 389116
rect 246390 389104 246396 389116
rect 246448 389144 246454 389156
rect 246574 389144 246580 389156
rect 246448 389116 246580 389144
rect 246448 389104 246454 389116
rect 246574 389104 246580 389116
rect 246632 389104 246638 389156
rect 48222 389036 48228 389088
rect 48280 389076 48286 389088
rect 72510 389076 72516 389088
rect 48280 389048 72516 389076
rect 48280 389036 48286 389048
rect 72510 389036 72516 389048
rect 72568 389036 72574 389088
rect 111978 389036 111984 389088
rect 112036 389076 112042 389088
rect 133874 389076 133880 389088
rect 112036 389048 133880 389076
rect 112036 389036 112042 389048
rect 133874 389036 133880 389048
rect 133932 389076 133938 389088
rect 251818 389076 251824 389088
rect 133932 389048 251824 389076
rect 133932 389036 133938 389048
rect 251818 389036 251824 389048
rect 251876 389036 251882 389088
rect 87598 387880 87604 387932
rect 87656 387920 87662 387932
rect 92014 387920 92020 387932
rect 87656 387892 92020 387920
rect 87656 387880 87662 387892
rect 92014 387880 92020 387892
rect 92072 387880 92078 387932
rect 71130 387812 71136 387864
rect 71188 387852 71194 387864
rect 71682 387852 71688 387864
rect 71188 387824 71688 387852
rect 71188 387812 71194 387824
rect 71682 387812 71688 387824
rect 71740 387812 71746 387864
rect 78122 387812 78128 387864
rect 78180 387852 78186 387864
rect 78582 387852 78588 387864
rect 78180 387824 78588 387852
rect 78180 387812 78186 387824
rect 78582 387812 78588 387824
rect 78640 387812 78646 387864
rect 79962 387812 79968 387864
rect 80020 387852 80026 387864
rect 81526 387852 81532 387864
rect 80020 387824 81532 387852
rect 80020 387812 80026 387824
rect 81526 387812 81532 387824
rect 81584 387812 81590 387864
rect 86218 387812 86224 387864
rect 86276 387852 86282 387864
rect 87782 387852 87788 387864
rect 86276 387824 87788 387852
rect 86276 387812 86282 387824
rect 87782 387812 87788 387824
rect 87840 387812 87846 387864
rect 249242 387812 249248 387864
rect 249300 387852 249306 387864
rect 251358 387852 251364 387864
rect 249300 387824 251364 387852
rect 249300 387812 249306 387824
rect 251358 387812 251364 387824
rect 251416 387812 251422 387864
rect 7558 387744 7564 387796
rect 7616 387784 7622 387796
rect 93946 387784 93952 387796
rect 7616 387756 93952 387784
rect 7616 387744 7622 387756
rect 93946 387744 93952 387756
rect 94004 387784 94010 387796
rect 94498 387784 94504 387796
rect 94004 387756 94504 387784
rect 94004 387744 94010 387756
rect 94498 387744 94504 387756
rect 94556 387744 94562 387796
rect 100386 387744 100392 387796
rect 100444 387784 100450 387796
rect 121546 387784 121552 387796
rect 100444 387756 121552 387784
rect 100444 387744 100450 387756
rect 121546 387744 121552 387756
rect 121604 387784 121610 387796
rect 122190 387784 122196 387796
rect 121604 387756 122196 387784
rect 121604 387744 121610 387756
rect 122190 387744 122196 387756
rect 122248 387744 122254 387796
rect 186038 387132 186044 387184
rect 186096 387172 186102 387184
rect 220998 387172 221004 387184
rect 186096 387144 221004 387172
rect 186096 387132 186102 387144
rect 220998 387132 221004 387144
rect 221056 387132 221062 387184
rect 110414 387064 110420 387116
rect 110472 387104 110478 387116
rect 186958 387104 186964 387116
rect 110472 387076 186964 387104
rect 110472 387064 110478 387076
rect 186958 387064 186964 387076
rect 187016 387064 187022 387116
rect 192662 387064 192668 387116
rect 192720 387104 192726 387116
rect 214006 387104 214012 387116
rect 192720 387076 214012 387104
rect 192720 387064 192726 387076
rect 214006 387064 214012 387076
rect 214064 387104 214070 387116
rect 253474 387104 253480 387116
rect 214064 387076 253480 387104
rect 214064 387064 214070 387076
rect 253474 387064 253480 387076
rect 253532 387064 253538 387116
rect 226334 386996 226340 387048
rect 226392 387036 226398 387048
rect 227254 387036 227260 387048
rect 226392 387008 227260 387036
rect 226392 386996 226398 387008
rect 227254 386996 227260 387008
rect 227312 386996 227318 387048
rect 231210 386384 231216 386436
rect 231268 386424 231274 386436
rect 270494 386424 270500 386436
rect 231268 386396 270500 386424
rect 231268 386384 231274 386396
rect 270494 386384 270500 386396
rect 270552 386384 270558 386436
rect 43990 386316 43996 386368
rect 44048 386356 44054 386368
rect 89254 386356 89260 386368
rect 44048 386328 89260 386356
rect 44048 386316 44054 386328
rect 89254 386316 89260 386328
rect 89312 386316 89318 386368
rect 99650 386316 99656 386368
rect 99708 386356 99714 386368
rect 100846 386356 100852 386368
rect 99708 386328 100852 386356
rect 99708 386316 99714 386328
rect 100846 386316 100852 386328
rect 100904 386316 100910 386368
rect 105170 386316 105176 386368
rect 105228 386356 105234 386368
rect 124306 386356 124312 386368
rect 105228 386328 124312 386356
rect 105228 386316 105234 386328
rect 124306 386316 124312 386328
rect 124364 386356 124370 386368
rect 124858 386356 124864 386368
rect 124364 386328 124864 386356
rect 124364 386316 124370 386328
rect 124858 386316 124864 386328
rect 124916 386316 124922 386368
rect 131758 386316 131764 386368
rect 131816 386356 131822 386368
rect 256878 386356 256884 386368
rect 131816 386328 256884 386356
rect 131816 386316 131822 386328
rect 256878 386316 256884 386328
rect 256936 386316 256942 386368
rect 240778 386248 240784 386300
rect 240836 386288 240842 386300
rect 247034 386288 247040 386300
rect 240836 386260 247040 386288
rect 240836 386248 240842 386260
rect 247034 386248 247040 386260
rect 247092 386248 247098 386300
rect 82078 385636 82084 385688
rect 82136 385676 82142 385688
rect 91094 385676 91100 385688
rect 82136 385648 91100 385676
rect 82136 385636 82142 385648
rect 91094 385636 91100 385648
rect 91152 385636 91158 385688
rect 101950 385636 101956 385688
rect 102008 385676 102014 385688
rect 112714 385676 112720 385688
rect 102008 385648 112720 385676
rect 102008 385636 102014 385648
rect 112714 385636 112720 385648
rect 112772 385636 112778 385688
rect 197998 385636 198004 385688
rect 198056 385676 198062 385688
rect 203886 385676 203892 385688
rect 198056 385648 203892 385676
rect 198056 385636 198062 385648
rect 203886 385636 203892 385648
rect 203944 385636 203950 385688
rect 232498 385024 232504 385076
rect 232556 385064 232562 385076
rect 239030 385064 239036 385076
rect 232556 385036 239036 385064
rect 232556 385024 232562 385036
rect 239030 385024 239036 385036
rect 239088 385024 239094 385076
rect 289906 385024 289912 385076
rect 289964 385064 289970 385076
rect 582558 385064 582564 385076
rect 289964 385036 582564 385064
rect 289964 385024 289970 385036
rect 582558 385024 582564 385036
rect 582616 385024 582622 385076
rect 56502 384956 56508 385008
rect 56560 384996 56566 385008
rect 86218 384996 86224 385008
rect 56560 384968 86224 384996
rect 56560 384956 56566 384968
rect 86218 384956 86224 384968
rect 86276 384956 86282 385008
rect 100938 384956 100944 385008
rect 100996 384996 101002 385008
rect 236638 384996 236644 385008
rect 100996 384968 236644 384996
rect 100996 384956 101002 384968
rect 236638 384956 236644 384968
rect 236696 384956 236702 385008
rect 66162 384888 66168 384940
rect 66220 384928 66226 384940
rect 87598 384928 87604 384940
rect 66220 384900 87604 384928
rect 66220 384888 66226 384900
rect 87598 384888 87604 384900
rect 87656 384888 87662 384940
rect 89162 384888 89168 384940
rect 89220 384928 89226 384940
rect 126882 384928 126888 384940
rect 89220 384900 126888 384928
rect 89220 384888 89226 384900
rect 126882 384888 126888 384900
rect 126940 384888 126946 384940
rect 148318 384888 148324 384940
rect 148376 384928 148382 384940
rect 148962 384928 148968 384940
rect 148376 384900 148968 384928
rect 148376 384888 148382 384900
rect 148962 384888 148968 384900
rect 149020 384928 149026 384940
rect 258166 384928 258172 384940
rect 149020 384900 258172 384928
rect 149020 384888 149026 384900
rect 258166 384888 258172 384900
rect 258224 384888 258230 384940
rect 236638 384276 236644 384328
rect 236696 384316 236702 384328
rect 266538 384316 266544 384328
rect 236696 384288 266544 384316
rect 236696 384276 236702 384288
rect 266538 384276 266544 384288
rect 266596 384276 266602 384328
rect 279418 384276 279424 384328
rect 279476 384316 279482 384328
rect 582926 384316 582932 384328
rect 279476 384288 582932 384316
rect 279476 384276 279482 384288
rect 582926 384276 582932 384288
rect 582984 384276 582990 384328
rect 189810 383596 189816 383648
rect 189868 383636 189874 383648
rect 252738 383636 252744 383648
rect 189868 383608 252744 383636
rect 189868 383596 189874 383608
rect 252738 383596 252744 383608
rect 252796 383636 252802 383648
rect 255314 383636 255320 383648
rect 252796 383608 255320 383636
rect 252796 383596 252802 383608
rect 255314 383596 255320 383608
rect 255372 383596 255378 383648
rect 97902 382916 97908 382968
rect 97960 382956 97966 382968
rect 128354 382956 128360 382968
rect 97960 382928 128360 382956
rect 97960 382916 97966 382928
rect 128354 382916 128360 382928
rect 128412 382916 128418 382968
rect 251818 382916 251824 382968
rect 251876 382956 251882 382968
rect 267826 382956 267832 382968
rect 251876 382928 267832 382956
rect 251876 382916 251882 382928
rect 267826 382916 267832 382928
rect 267884 382916 267890 382968
rect 3510 382236 3516 382288
rect 3568 382276 3574 382288
rect 113174 382276 113180 382288
rect 3568 382248 113180 382276
rect 3568 382236 3574 382248
rect 113174 382236 113180 382248
rect 113232 382276 113238 382288
rect 113450 382276 113456 382288
rect 113232 382248 113456 382276
rect 113232 382236 113238 382248
rect 113450 382236 113456 382248
rect 113508 382236 113514 382288
rect 128354 382236 128360 382288
rect 128412 382276 128418 382288
rect 231854 382276 231860 382288
rect 128412 382248 231860 382276
rect 128412 382236 128418 382248
rect 231854 382236 231860 382248
rect 231912 382236 231918 382288
rect 252738 382276 252744 382288
rect 251836 382248 252744 382276
rect 251836 382220 251864 382248
rect 252738 382236 252744 382248
rect 252796 382236 252802 382288
rect 101030 382168 101036 382220
rect 101088 382208 101094 382220
rect 122098 382208 122104 382220
rect 101088 382180 122104 382208
rect 101088 382168 101094 382180
rect 122098 382168 122104 382180
rect 122156 382168 122162 382220
rect 126882 382168 126888 382220
rect 126940 382208 126946 382220
rect 186038 382208 186044 382220
rect 126940 382180 186044 382208
rect 126940 382168 126946 382180
rect 186038 382168 186044 382180
rect 186096 382168 186102 382220
rect 251818 382168 251824 382220
rect 251876 382168 251882 382220
rect 187510 381556 187516 381608
rect 187568 381596 187574 381608
rect 194594 381596 194600 381608
rect 187568 381568 194600 381596
rect 187568 381556 187574 381568
rect 194594 381556 194600 381568
rect 194652 381556 194658 381608
rect 101398 381488 101404 381540
rect 101456 381528 101462 381540
rect 113542 381528 113548 381540
rect 101456 381500 113548 381528
rect 101456 381488 101462 381500
rect 113542 381488 113548 381500
rect 113600 381488 113606 381540
rect 191742 381488 191748 381540
rect 191800 381528 191806 381540
rect 264974 381528 264980 381540
rect 191800 381500 264980 381528
rect 191800 381488 191806 381500
rect 264974 381488 264980 381500
rect 265032 381488 265038 381540
rect 186038 380876 186044 380928
rect 186096 380916 186102 380928
rect 186314 380916 186320 380928
rect 186096 380888 186320 380916
rect 186096 380876 186102 380888
rect 186314 380876 186320 380888
rect 186372 380876 186378 380928
rect 198734 380876 198740 380928
rect 198792 380916 198798 380928
rect 276014 380916 276020 380928
rect 198792 380888 276020 380916
rect 198792 380876 198798 380888
rect 276014 380876 276020 380888
rect 276072 380876 276078 380928
rect 105538 380808 105544 380860
rect 105596 380848 105602 380860
rect 231210 380848 231216 380860
rect 105596 380820 231216 380848
rect 105596 380808 105602 380820
rect 231210 380808 231216 380820
rect 231268 380808 231274 380860
rect 274726 380808 274732 380860
rect 274784 380848 274790 380860
rect 582374 380848 582380 380860
rect 274784 380820 582380 380848
rect 274784 380808 274790 380820
rect 582374 380808 582380 380820
rect 582432 380808 582438 380860
rect 193398 380740 193404 380792
rect 193456 380780 193462 380792
rect 255590 380780 255596 380792
rect 193456 380752 255596 380780
rect 193456 380740 193462 380752
rect 255590 380740 255596 380752
rect 255648 380740 255654 380792
rect 188982 380264 188988 380316
rect 189040 380304 189046 380316
rect 192570 380304 192576 380316
rect 189040 380276 192576 380304
rect 189040 380264 189046 380276
rect 192570 380264 192576 380276
rect 192628 380264 192634 380316
rect 60550 380196 60556 380248
rect 60608 380236 60614 380248
rect 77478 380236 77484 380248
rect 60608 380208 77484 380236
rect 60608 380196 60614 380208
rect 77478 380196 77484 380208
rect 77536 380196 77542 380248
rect 73154 380128 73160 380180
rect 73212 380168 73218 380180
rect 168374 380168 168380 380180
rect 73212 380140 168380 380168
rect 73212 380128 73218 380140
rect 168374 380128 168380 380140
rect 168432 380128 168438 380180
rect 105998 379448 106004 379500
rect 106056 379488 106062 379500
rect 243078 379488 243084 379500
rect 106056 379460 243084 379488
rect 106056 379448 106062 379460
rect 243078 379448 243084 379460
rect 243136 379448 243142 379500
rect 67542 379380 67548 379432
rect 67600 379420 67606 379432
rect 155954 379420 155960 379432
rect 67600 379392 155960 379420
rect 67600 379380 67606 379392
rect 155954 379380 155960 379392
rect 156012 379420 156018 379432
rect 156598 379420 156604 379432
rect 156012 379392 156604 379420
rect 156012 379380 156018 379392
rect 156598 379380 156604 379392
rect 156656 379380 156662 379432
rect 173066 379380 173072 379432
rect 173124 379420 173130 379432
rect 173710 379420 173716 379432
rect 173124 379392 173716 379420
rect 173124 379380 173130 379392
rect 173710 379380 173716 379392
rect 173768 379420 173774 379432
rect 207014 379420 207020 379432
rect 173768 379392 207020 379420
rect 173768 379380 173774 379392
rect 207014 379380 207020 379392
rect 207072 379380 207078 379432
rect 243078 378972 243084 379024
rect 243136 379012 243142 379024
rect 243538 379012 243544 379024
rect 243136 378984 243544 379012
rect 243136 378972 243142 378984
rect 243538 378972 243544 378984
rect 243596 378972 243602 379024
rect 231854 378768 231860 378820
rect 231912 378808 231918 378820
rect 281718 378808 281724 378820
rect 231912 378780 281724 378808
rect 231912 378768 231918 378780
rect 281718 378768 281724 378780
rect 281776 378768 281782 378820
rect 106918 377476 106924 377528
rect 106976 377516 106982 377528
rect 116026 377516 116032 377528
rect 106976 377488 116032 377516
rect 106976 377476 106982 377488
rect 116026 377476 116032 377488
rect 116084 377476 116090 377528
rect 78582 377408 78588 377460
rect 78640 377448 78646 377460
rect 176470 377448 176476 377460
rect 78640 377420 176476 377448
rect 78640 377408 78646 377420
rect 176470 377408 176476 377420
rect 176528 377448 176534 377460
rect 205634 377448 205640 377460
rect 176528 377420 205640 377448
rect 176528 377408 176534 377420
rect 205634 377408 205640 377420
rect 205692 377408 205698 377460
rect 3418 376660 3424 376712
rect 3476 376700 3482 376712
rect 116118 376700 116124 376712
rect 3476 376672 116124 376700
rect 3476 376660 3482 376672
rect 116118 376660 116124 376672
rect 116176 376660 116182 376712
rect 152458 376660 152464 376712
rect 152516 376700 152522 376712
rect 247034 376700 247040 376712
rect 152516 376672 247040 376700
rect 152516 376660 152522 376672
rect 247034 376660 247040 376672
rect 247092 376700 247098 376712
rect 247678 376700 247684 376712
rect 247092 376672 247684 376700
rect 247092 376660 247098 376672
rect 247678 376660 247684 376672
rect 247736 376660 247742 376712
rect 92474 376592 92480 376644
rect 92532 376632 92538 376644
rect 122926 376632 122932 376644
rect 92532 376604 122932 376632
rect 92532 376592 92538 376604
rect 122926 376592 122932 376604
rect 122984 376632 122990 376644
rect 123478 376632 123484 376644
rect 122984 376604 123484 376632
rect 122984 376592 122990 376604
rect 123478 376592 123484 376604
rect 123536 376592 123542 376644
rect 118602 375980 118608 376032
rect 118660 376020 118666 376032
rect 277486 376020 277492 376032
rect 118660 375992 277492 376020
rect 118660 375980 118666 375992
rect 277486 375980 277492 375992
rect 277544 375980 277550 376032
rect 87598 375300 87604 375352
rect 87656 375340 87662 375352
rect 88242 375340 88248 375352
rect 87656 375312 88248 375340
rect 87656 375300 87662 375312
rect 88242 375300 88248 375312
rect 88300 375340 88306 375352
rect 88300 375312 93854 375340
rect 88300 375300 88306 375312
rect 93826 375272 93854 375312
rect 107470 375300 107476 375352
rect 107528 375340 107534 375352
rect 245746 375340 245752 375352
rect 107528 375312 245752 375340
rect 107528 375300 107534 375312
rect 245746 375300 245752 375312
rect 245804 375300 245810 375352
rect 224954 375272 224960 375284
rect 93826 375244 224960 375272
rect 224954 375232 224960 375244
rect 225012 375232 225018 375284
rect 255682 374620 255688 374672
rect 255740 374660 255746 374672
rect 256786 374660 256792 374672
rect 255740 374632 256792 374660
rect 255740 374620 255746 374632
rect 256786 374620 256792 374632
rect 256844 374660 256850 374672
rect 291286 374660 291292 374672
rect 256844 374632 291292 374660
rect 256844 374620 256850 374632
rect 291286 374620 291292 374632
rect 291344 374620 291350 374672
rect 245746 374552 245752 374604
rect 245804 374592 245810 374604
rect 246298 374592 246304 374604
rect 245804 374564 246304 374592
rect 245804 374552 245810 374564
rect 246298 374552 246304 374564
rect 246356 374552 246362 374604
rect 122190 373940 122196 373992
rect 122248 373980 122254 373992
rect 235994 373980 236000 373992
rect 122248 373952 236000 373980
rect 122248 373940 122254 373952
rect 235994 373940 236000 373952
rect 236052 373940 236058 373992
rect 100570 373260 100576 373312
rect 100628 373300 100634 373312
rect 118602 373300 118608 373312
rect 100628 373272 118608 373300
rect 100628 373260 100634 373272
rect 118602 373260 118608 373272
rect 118660 373260 118666 373312
rect 208486 373260 208492 373312
rect 208544 373300 208550 373312
rect 284386 373300 284392 373312
rect 208544 373272 284392 373300
rect 208544 373260 208550 373272
rect 284386 373260 284392 373272
rect 284444 373260 284450 373312
rect 235994 372580 236000 372632
rect 236052 372620 236058 372632
rect 236638 372620 236644 372632
rect 236052 372592 236644 372620
rect 236052 372580 236058 372592
rect 236638 372580 236644 372592
rect 236696 372580 236702 372632
rect 111794 372512 111800 372564
rect 111852 372552 111858 372564
rect 112530 372552 112536 372564
rect 111852 372524 112536 372552
rect 111852 372512 111858 372524
rect 112530 372512 112536 372524
rect 112588 372552 112594 372564
rect 252646 372552 252652 372564
rect 112588 372524 252652 372552
rect 112588 372512 112594 372524
rect 252646 372512 252652 372524
rect 252704 372512 252710 372564
rect 75914 372444 75920 372496
rect 75972 372484 75978 372496
rect 197998 372484 198004 372496
rect 75972 372456 198004 372484
rect 75972 372444 75978 372456
rect 197998 372444 198004 372456
rect 198056 372444 198062 372496
rect 209774 371832 209780 371884
rect 209832 371872 209838 371884
rect 278866 371872 278872 371884
rect 209832 371844 278872 371872
rect 209832 371832 209838 371844
rect 278866 371832 278872 371844
rect 278924 371832 278930 371884
rect 114462 371152 114468 371204
rect 114520 371192 114526 371204
rect 259638 371192 259644 371204
rect 114520 371164 259644 371192
rect 114520 371152 114526 371164
rect 259638 371152 259644 371164
rect 259696 371192 259702 371204
rect 260742 371192 260748 371204
rect 259696 371164 260748 371192
rect 259696 371152 259702 371164
rect 260742 371152 260748 371164
rect 260800 371152 260806 371204
rect 104158 370540 104164 370592
rect 104216 370580 104222 370592
rect 113174 370580 113180 370592
rect 104216 370552 113180 370580
rect 104216 370540 104222 370552
rect 113174 370540 113180 370552
rect 113232 370580 113238 370592
rect 114462 370580 114468 370592
rect 113232 370552 114468 370580
rect 113232 370540 113238 370552
rect 114462 370540 114468 370552
rect 114520 370540 114526 370592
rect 94038 370472 94044 370524
rect 94096 370512 94102 370524
rect 107654 370512 107660 370524
rect 94096 370484 107660 370512
rect 94096 370472 94102 370484
rect 107654 370472 107660 370484
rect 107712 370472 107718 370524
rect 155218 370472 155224 370524
rect 155276 370512 155282 370524
rect 252462 370512 252468 370524
rect 155276 370484 252468 370512
rect 155276 370472 155282 370484
rect 252462 370472 252468 370484
rect 252520 370512 252526 370524
rect 255406 370512 255412 370524
rect 252520 370484 255412 370512
rect 252520 370472 252526 370484
rect 255406 370472 255412 370484
rect 255464 370472 255470 370524
rect 260742 370472 260748 370524
rect 260800 370512 260806 370524
rect 281810 370512 281816 370524
rect 260800 370484 281816 370512
rect 260800 370472 260806 370484
rect 281810 370472 281816 370484
rect 281868 370472 281874 370524
rect 196066 369180 196072 369232
rect 196124 369220 196130 369232
rect 240226 369220 240232 369232
rect 196124 369192 240232 369220
rect 196124 369180 196130 369192
rect 240226 369180 240232 369192
rect 240284 369180 240290 369232
rect 102134 369112 102140 369164
rect 102192 369152 102198 369164
rect 137462 369152 137468 369164
rect 102192 369124 137468 369152
rect 102192 369112 102198 369124
rect 137462 369112 137468 369124
rect 137520 369152 137526 369164
rect 232498 369152 232504 369164
rect 137520 369124 232504 369152
rect 137520 369112 137526 369124
rect 232498 369112 232504 369124
rect 232556 369112 232562 369164
rect 130470 368432 130476 368484
rect 130528 368472 130534 368484
rect 231118 368472 231124 368484
rect 130528 368444 231124 368472
rect 130528 368432 130534 368444
rect 231118 368432 231124 368444
rect 231176 368432 231182 368484
rect 89070 367820 89076 367872
rect 89128 367860 89134 367872
rect 128998 367860 129004 367872
rect 89128 367832 129004 367860
rect 89128 367820 89134 367832
rect 128998 367820 129004 367832
rect 129056 367820 129062 367872
rect 232498 367820 232504 367872
rect 232556 367860 232562 367872
rect 262214 367860 262220 367872
rect 232556 367832 262220 367860
rect 232556 367820 232562 367832
rect 262214 367820 262220 367832
rect 262272 367820 262278 367872
rect 74626 367752 74632 367804
rect 74684 367792 74690 367804
rect 152550 367792 152556 367804
rect 74684 367764 152556 367792
rect 74684 367752 74690 367764
rect 152550 367752 152556 367764
rect 152608 367792 152614 367804
rect 201494 367792 201500 367804
rect 152608 367764 201500 367792
rect 152608 367752 152614 367764
rect 201494 367752 201500 367764
rect 201552 367752 201558 367804
rect 254578 367752 254584 367804
rect 254636 367792 254642 367804
rect 582742 367792 582748 367804
rect 254636 367764 582748 367792
rect 254636 367752 254642 367764
rect 582742 367752 582748 367764
rect 582800 367752 582806 367804
rect 204254 367004 204260 367056
rect 204312 367044 204318 367056
rect 582466 367044 582472 367056
rect 204312 367016 582472 367044
rect 204312 367004 204318 367016
rect 582466 367004 582472 367016
rect 582524 367004 582530 367056
rect 107746 366392 107752 366444
rect 107804 366432 107810 366444
rect 180794 366432 180800 366444
rect 107804 366404 180800 366432
rect 107804 366392 107810 366404
rect 180794 366392 180800 366404
rect 180852 366432 180858 366444
rect 181346 366432 181352 366444
rect 180852 366404 181352 366432
rect 180852 366392 180858 366404
rect 181346 366392 181352 366404
rect 181404 366392 181410 366444
rect 45370 366324 45376 366376
rect 45428 366364 45434 366376
rect 75914 366364 75920 366376
rect 45428 366336 75920 366364
rect 45428 366324 45434 366336
rect 75914 366324 75920 366336
rect 75972 366324 75978 366376
rect 82814 366324 82820 366376
rect 82872 366364 82878 366376
rect 156598 366364 156604 366376
rect 82872 366336 156604 366364
rect 82872 366324 82878 366336
rect 156598 366324 156604 366336
rect 156656 366364 156662 366376
rect 213914 366364 213920 366376
rect 156656 366336 213920 366364
rect 156656 366324 156662 366336
rect 213914 366324 213920 366336
rect 213972 366324 213978 366376
rect 63310 365644 63316 365696
rect 63368 365684 63374 365696
rect 184290 365684 184296 365696
rect 63368 365656 184296 365684
rect 63368 365644 63374 365656
rect 184290 365644 184296 365656
rect 184348 365644 184354 365696
rect 220722 365644 220728 365696
rect 220780 365684 220786 365696
rect 240778 365684 240784 365696
rect 220780 365656 240784 365684
rect 220780 365644 220786 365656
rect 240778 365644 240784 365656
rect 240836 365644 240842 365696
rect 182910 364964 182916 365016
rect 182968 365004 182974 365016
rect 229094 365004 229100 365016
rect 182968 364976 229100 365004
rect 182968 364964 182974 364976
rect 229094 364964 229100 364976
rect 229152 364964 229158 365016
rect 193398 363740 193404 363792
rect 193456 363780 193462 363792
rect 195974 363780 195980 363792
rect 193456 363752 195980 363780
rect 193456 363740 193462 363752
rect 195974 363740 195980 363752
rect 196032 363740 196038 363792
rect 253842 363780 253848 363792
rect 238726 363752 253848 363780
rect 151170 363672 151176 363724
rect 151228 363712 151234 363724
rect 238726 363712 238754 363752
rect 253842 363740 253848 363752
rect 253900 363780 253906 363792
rect 255498 363780 255504 363792
rect 253900 363752 255504 363780
rect 253900 363740 253906 363752
rect 255498 363740 255504 363752
rect 255556 363740 255562 363792
rect 151228 363684 238754 363712
rect 151228 363672 151234 363684
rect 71682 363604 71688 363656
rect 71740 363644 71746 363656
rect 193398 363644 193404 363656
rect 71740 363616 193404 363644
rect 71740 363604 71746 363616
rect 193398 363604 193404 363616
rect 193456 363604 193462 363656
rect 116578 362856 116584 362908
rect 116636 362896 116642 362908
rect 252554 362896 252560 362908
rect 116636 362868 252560 362896
rect 116636 362856 116642 362868
rect 252554 362856 252560 362868
rect 252612 362856 252618 362908
rect 86218 362788 86224 362840
rect 86276 362828 86282 362840
rect 219526 362828 219532 362840
rect 86276 362800 219532 362828
rect 86276 362788 86282 362800
rect 219526 362788 219532 362800
rect 219584 362828 219590 362840
rect 220078 362828 220084 362840
rect 219584 362800 220084 362828
rect 219584 362788 219590 362800
rect 220078 362788 220084 362800
rect 220136 362788 220142 362840
rect 85574 361496 85580 361548
rect 85632 361536 85638 361548
rect 216674 361536 216680 361548
rect 85632 361508 216680 361536
rect 85632 361496 85638 361508
rect 216674 361496 216680 361508
rect 216732 361496 216738 361548
rect 123478 361428 123484 361480
rect 123536 361468 123542 361480
rect 226426 361468 226432 361480
rect 123536 361440 226432 361468
rect 123536 361428 123542 361440
rect 226426 361428 226432 361440
rect 226484 361428 226490 361480
rect 232590 360816 232596 360868
rect 232648 360856 232654 360868
rect 263778 360856 263784 360868
rect 232648 360828 263784 360856
rect 232648 360816 232654 360828
rect 263778 360816 263784 360828
rect 263836 360816 263842 360868
rect 226426 360204 226432 360256
rect 226484 360244 226490 360256
rect 226978 360244 226984 360256
rect 226484 360216 226984 360244
rect 226484 360204 226490 360216
rect 226978 360204 226984 360216
rect 227036 360204 227042 360256
rect 94498 359524 94504 359576
rect 94556 359564 94562 359576
rect 124214 359564 124220 359576
rect 94556 359536 124220 359564
rect 94556 359524 94562 359536
rect 124214 359524 124220 359536
rect 124272 359564 124278 359576
rect 125042 359564 125048 359576
rect 124272 359536 125048 359564
rect 124272 359524 124278 359536
rect 125042 359524 125048 359536
rect 125100 359524 125106 359576
rect 56410 359456 56416 359508
rect 56468 359496 56474 359508
rect 184382 359496 184388 359508
rect 56468 359468 184388 359496
rect 56468 359456 56474 359468
rect 184382 359456 184388 359468
rect 184440 359456 184446 359508
rect 215386 359456 215392 359508
rect 215444 359496 215450 359508
rect 242894 359496 242900 359508
rect 215444 359468 242900 359496
rect 215444 359456 215450 359468
rect 242894 359456 242900 359468
rect 242952 359456 242958 359508
rect 125042 358776 125048 358828
rect 125100 358816 125106 358828
rect 226334 358816 226340 358828
rect 125100 358788 226340 358816
rect 125100 358776 125106 358788
rect 226334 358776 226340 358788
rect 226392 358776 226398 358828
rect 84194 358708 84200 358760
rect 84252 358748 84258 358760
rect 215294 358748 215300 358760
rect 84252 358720 215300 358748
rect 84252 358708 84258 358720
rect 215294 358708 215300 358720
rect 215352 358748 215358 358760
rect 215938 358748 215944 358760
rect 215352 358720 215944 358748
rect 215352 358708 215358 358720
rect 215938 358708 215944 358720
rect 215996 358708 216002 358760
rect 2774 358436 2780 358488
rect 2832 358476 2838 358488
rect 4798 358476 4804 358488
rect 2832 358448 4804 358476
rect 2832 358436 2838 358448
rect 4798 358436 4804 358448
rect 4856 358436 4862 358488
rect 103514 357348 103520 357400
rect 103572 357388 103578 357400
rect 240134 357388 240140 357400
rect 103572 357360 240140 357388
rect 103572 357348 103578 357360
rect 240134 357348 240140 357360
rect 240192 357388 240198 357400
rect 240778 357388 240784 357400
rect 240192 357360 240784 357388
rect 240192 357348 240198 357360
rect 240778 357348 240784 357360
rect 240836 357348 240842 357400
rect 226334 356668 226340 356720
rect 226392 356708 226398 356720
rect 262214 356708 262220 356720
rect 226392 356680 262220 356708
rect 226392 356668 226398 356680
rect 262214 356668 262220 356680
rect 262272 356668 262278 356720
rect 128998 355988 129004 356040
rect 129056 356028 129062 356040
rect 220906 356028 220912 356040
rect 129056 356000 220912 356028
rect 129056 355988 129062 356000
rect 220906 355988 220912 356000
rect 220964 356028 220970 356040
rect 221550 356028 221556 356040
rect 220964 356000 221556 356028
rect 220964 355988 220970 356000
rect 221550 355988 221556 356000
rect 221608 355988 221614 356040
rect 75730 355308 75736 355360
rect 75788 355348 75794 355360
rect 193306 355348 193312 355360
rect 75788 355320 193312 355348
rect 75788 355308 75794 355320
rect 193306 355308 193312 355320
rect 193364 355348 193370 355360
rect 202874 355348 202880 355360
rect 193364 355320 202880 355348
rect 193364 355308 193370 355320
rect 202874 355308 202880 355320
rect 202932 355308 202938 355360
rect 79962 354628 79968 354680
rect 80020 354668 80026 354680
rect 211154 354668 211160 354680
rect 80020 354640 211160 354668
rect 80020 354628 80026 354640
rect 211154 354628 211160 354640
rect 211212 354628 211218 354680
rect 81526 353948 81532 354000
rect 81584 353988 81590 354000
rect 102134 353988 102140 354000
rect 81584 353960 102140 353988
rect 81584 353948 81590 353960
rect 102134 353948 102140 353960
rect 102192 353988 102198 354000
rect 212534 353988 212540 354000
rect 102192 353960 212540 353988
rect 102192 353948 102198 353960
rect 212534 353948 212540 353960
rect 212592 353948 212598 354000
rect 222194 353268 222200 353320
rect 222252 353308 222258 353320
rect 231118 353308 231124 353320
rect 222252 353280 231124 353308
rect 222252 353268 222258 353280
rect 231118 353268 231124 353280
rect 231176 353268 231182 353320
rect 249702 353268 249708 353320
rect 249760 353308 249766 353320
rect 252554 353308 252560 353320
rect 249760 353280 252560 353308
rect 249760 353268 249766 353280
rect 252554 353268 252560 353280
rect 252612 353268 252618 353320
rect 111058 353200 111064 353252
rect 111116 353240 111122 353252
rect 249242 353240 249248 353252
rect 111116 353212 249248 353240
rect 111116 353200 111122 353212
rect 249242 353200 249248 353212
rect 249300 353200 249306 353252
rect 110506 352860 110512 352912
rect 110564 352900 110570 352912
rect 111058 352900 111064 352912
rect 110564 352872 111064 352900
rect 110564 352860 110570 352872
rect 111058 352860 111064 352872
rect 111116 352860 111122 352912
rect 155862 352520 155868 352572
rect 155920 352560 155926 352572
rect 194594 352560 194600 352572
rect 155920 352532 194600 352560
rect 155920 352520 155926 352532
rect 194594 352520 194600 352532
rect 194652 352560 194658 352572
rect 222838 352560 222844 352572
rect 194652 352532 222844 352560
rect 194652 352520 194658 352532
rect 222838 352520 222844 352532
rect 222896 352520 222902 352572
rect 95142 351840 95148 351892
rect 95200 351880 95206 351892
rect 182174 351880 182180 351892
rect 95200 351852 182180 351880
rect 95200 351840 95206 351852
rect 182174 351840 182180 351852
rect 182232 351880 182238 351892
rect 182910 351880 182916 351892
rect 182232 351852 182916 351880
rect 182232 351840 182238 351852
rect 182910 351840 182916 351852
rect 182968 351840 182974 351892
rect 186958 351840 186964 351892
rect 187016 351880 187022 351892
rect 187510 351880 187516 351892
rect 187016 351852 187516 351880
rect 187016 351840 187022 351852
rect 187510 351840 187516 351852
rect 187568 351880 187574 351892
rect 249794 351880 249800 351892
rect 187568 351852 249800 351880
rect 187568 351840 187574 351852
rect 249794 351840 249800 351852
rect 249852 351840 249858 351892
rect 195238 349868 195244 349920
rect 195296 349908 195302 349920
rect 249150 349908 249156 349920
rect 195296 349880 249156 349908
rect 195296 349868 195302 349880
rect 249150 349868 249156 349880
rect 249208 349868 249214 349920
rect 154482 349800 154488 349852
rect 154540 349840 154546 349852
rect 270586 349840 270592 349852
rect 154540 349812 270592 349840
rect 154540 349800 154546 349812
rect 270586 349800 270592 349812
rect 270644 349800 270650 349852
rect 196618 348372 196624 348424
rect 196676 348412 196682 348424
rect 238018 348412 238024 348424
rect 196676 348384 238024 348412
rect 196676 348372 196682 348384
rect 238018 348372 238024 348384
rect 238076 348372 238082 348424
rect 67450 347760 67456 347812
rect 67508 347800 67514 347812
rect 294046 347800 294052 347812
rect 67508 347772 294052 347800
rect 67508 347760 67514 347772
rect 294046 347760 294052 347772
rect 294104 347760 294110 347812
rect 123570 346468 123576 346520
rect 123628 346508 123634 346520
rect 211154 346508 211160 346520
rect 123628 346480 211160 346508
rect 123628 346468 123634 346480
rect 211154 346468 211160 346480
rect 211212 346508 211218 346520
rect 211798 346508 211804 346520
rect 211212 346480 211804 346508
rect 211212 346468 211218 346480
rect 211798 346468 211804 346480
rect 211856 346468 211862 346520
rect 142982 346400 142988 346452
rect 143040 346440 143046 346452
rect 234798 346440 234804 346452
rect 143040 346412 234804 346440
rect 143040 346400 143046 346412
rect 234798 346400 234804 346412
rect 234856 346400 234862 346452
rect 141602 345108 141608 345160
rect 141660 345148 141666 345160
rect 234706 345148 234712 345160
rect 141660 345120 234712 345148
rect 141660 345108 141666 345120
rect 234706 345108 234712 345120
rect 234764 345108 234770 345160
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 11698 345080 11704 345092
rect 3384 345052 11704 345080
rect 3384 345040 3390 345052
rect 11698 345040 11704 345052
rect 11756 345040 11762 345092
rect 88978 345040 88984 345092
rect 89036 345080 89042 345092
rect 292574 345080 292580 345092
rect 89036 345052 292580 345080
rect 89036 345040 89042 345052
rect 292574 345040 292580 345052
rect 292632 345040 292638 345092
rect 141418 343680 141424 343732
rect 141476 343720 141482 343732
rect 142062 343720 142068 343732
rect 141476 343692 142068 343720
rect 141476 343680 141482 343692
rect 142062 343680 142068 343692
rect 142120 343720 142126 343732
rect 291378 343720 291384 343732
rect 142120 343692 291384 343720
rect 142120 343680 142126 343692
rect 291378 343680 291384 343692
rect 291436 343680 291442 343732
rect 37182 343612 37188 343664
rect 37240 343652 37246 343664
rect 204254 343652 204260 343664
rect 37240 343624 204260 343652
rect 37240 343612 37246 343624
rect 204254 343612 204260 343624
rect 204312 343612 204318 343664
rect 172422 342864 172428 342916
rect 172480 342904 172486 342916
rect 183462 342904 183468 342916
rect 172480 342876 183468 342904
rect 172480 342864 172486 342876
rect 183462 342864 183468 342876
rect 183520 342904 183526 342916
rect 224218 342904 224224 342916
rect 183520 342876 224224 342904
rect 183520 342864 183526 342876
rect 224218 342864 224224 342876
rect 224276 342864 224282 342916
rect 227714 342864 227720 342916
rect 227772 342904 227778 342916
rect 253198 342904 253204 342916
rect 227772 342876 253204 342904
rect 227772 342864 227778 342876
rect 253198 342864 253204 342876
rect 253256 342864 253262 342916
rect 88242 342252 88248 342304
rect 88300 342292 88306 342304
rect 233970 342292 233976 342304
rect 88300 342264 233976 342292
rect 88300 342252 88306 342264
rect 233970 342252 233976 342264
rect 234028 342252 234034 342304
rect 184750 341504 184756 341556
rect 184808 341544 184814 341556
rect 208394 341544 208400 341556
rect 184808 341516 208400 341544
rect 184808 341504 184814 341516
rect 208394 341504 208400 341516
rect 208452 341504 208458 341556
rect 244366 341504 244372 341556
rect 244424 341544 244430 341556
rect 263594 341544 263600 341556
rect 244424 341516 263600 341544
rect 244424 341504 244430 341516
rect 263594 341504 263600 341516
rect 263652 341504 263658 341556
rect 130470 340892 130476 340944
rect 130528 340932 130534 340944
rect 244366 340932 244372 340944
rect 130528 340904 244372 340932
rect 130528 340892 130534 340904
rect 244366 340892 244372 340904
rect 244424 340892 244430 340944
rect 170950 340144 170956 340196
rect 171008 340184 171014 340196
rect 244274 340184 244280 340196
rect 171008 340156 244280 340184
rect 171008 340144 171014 340156
rect 244274 340144 244280 340156
rect 244332 340144 244338 340196
rect 159542 339464 159548 339516
rect 159600 339504 159606 339516
rect 295518 339504 295524 339516
rect 159600 339476 295524 339504
rect 159600 339464 159606 339476
rect 295518 339464 295524 339476
rect 295576 339464 295582 339516
rect 124858 338172 124864 338224
rect 124916 338212 124922 338224
rect 229094 338212 229100 338224
rect 124916 338184 229100 338212
rect 124916 338172 124922 338184
rect 229094 338172 229100 338184
rect 229152 338172 229158 338224
rect 112438 338104 112444 338156
rect 112496 338144 112502 338156
rect 238754 338144 238760 338156
rect 112496 338116 238760 338144
rect 112496 338104 112502 338116
rect 238754 338104 238760 338116
rect 238812 338144 238818 338156
rect 239398 338144 239404 338156
rect 238812 338116 239404 338144
rect 238812 338104 238818 338116
rect 239398 338104 239404 338116
rect 239456 338104 239462 338156
rect 184842 337424 184848 337476
rect 184900 337464 184906 337476
rect 232590 337464 232596 337476
rect 184900 337436 232596 337464
rect 184900 337424 184906 337436
rect 232590 337424 232596 337436
rect 232648 337424 232654 337476
rect 223482 337356 223488 337408
rect 223540 337396 223546 337408
rect 272058 337396 272064 337408
rect 223540 337368 272064 337396
rect 223540 337356 223546 337368
rect 272058 337356 272064 337368
rect 272116 337356 272122 337408
rect 42702 336744 42708 336796
rect 42760 336784 42766 336796
rect 221458 336784 221464 336796
rect 42760 336756 221464 336784
rect 42760 336744 42766 336756
rect 221458 336744 221464 336756
rect 221516 336744 221522 336796
rect 190362 335996 190368 336048
rect 190420 336036 190426 336048
rect 280246 336036 280252 336048
rect 190420 336008 280252 336036
rect 190420 335996 190426 336008
rect 280246 335996 280252 336008
rect 280304 335996 280310 336048
rect 108942 335724 108948 335776
rect 109000 335764 109006 335776
rect 112530 335764 112536 335776
rect 109000 335736 112536 335764
rect 109000 335724 109006 335736
rect 112530 335724 112536 335736
rect 112588 335724 112594 335776
rect 155310 335316 155316 335368
rect 155368 335356 155374 335368
rect 251818 335356 251824 335368
rect 155368 335328 251824 335356
rect 155368 335316 155374 335328
rect 251818 335316 251824 335328
rect 251876 335316 251882 335368
rect 184290 334568 184296 334620
rect 184348 334608 184354 334620
rect 274726 334608 274732 334620
rect 184348 334580 274732 334608
rect 184348 334568 184354 334580
rect 274726 334568 274732 334580
rect 274784 334568 274790 334620
rect 145650 333956 145656 334008
rect 145708 333996 145714 334008
rect 247034 333996 247040 334008
rect 145708 333968 247040 333996
rect 145708 333956 145714 333968
rect 247034 333956 247040 333968
rect 247092 333996 247098 334008
rect 247678 333996 247684 334008
rect 247092 333968 247684 333996
rect 247092 333956 247098 333968
rect 247678 333956 247684 333968
rect 247736 333956 247742 334008
rect 183462 333208 183468 333260
rect 183520 333248 183526 333260
rect 232498 333248 232504 333260
rect 183520 333220 232504 333248
rect 183520 333208 183526 333220
rect 232498 333208 232504 333220
rect 232556 333208 232562 333260
rect 152642 332596 152648 332648
rect 152700 332636 152706 332648
rect 233142 332636 233148 332648
rect 152700 332608 233148 332636
rect 152700 332596 152706 332608
rect 233142 332596 233148 332608
rect 233200 332636 233206 332648
rect 233878 332636 233884 332648
rect 233200 332608 233884 332636
rect 233200 332596 233206 332608
rect 233878 332596 233884 332608
rect 233936 332596 233942 332648
rect 174630 331304 174636 331356
rect 174688 331344 174694 331356
rect 242894 331344 242900 331356
rect 174688 331316 242900 331344
rect 174688 331304 174694 331316
rect 242894 331304 242900 331316
rect 242952 331304 242958 331356
rect 173618 331236 173624 331288
rect 173676 331276 173682 331288
rect 245654 331276 245660 331288
rect 173676 331248 245660 331276
rect 173676 331236 173682 331248
rect 245654 331236 245660 331248
rect 245712 331236 245718 331288
rect 246390 330488 246396 330540
rect 246448 330528 246454 330540
rect 270586 330528 270592 330540
rect 246448 330500 270592 330528
rect 246448 330488 246454 330500
rect 270586 330488 270592 330500
rect 270644 330488 270650 330540
rect 177482 329876 177488 329928
rect 177540 329916 177546 329928
rect 177942 329916 177948 329928
rect 177540 329888 177948 329916
rect 177540 329876 177546 329888
rect 177942 329876 177948 329888
rect 178000 329916 178006 329928
rect 232498 329916 232504 329928
rect 178000 329888 232504 329916
rect 178000 329876 178006 329888
rect 232498 329876 232504 329888
rect 232556 329876 232562 329928
rect 177298 329808 177304 329860
rect 177356 329848 177362 329860
rect 240226 329848 240232 329860
rect 177356 329820 240232 329848
rect 177356 329808 177362 329820
rect 240226 329808 240232 329820
rect 240284 329808 240290 329860
rect 166350 329332 166356 329384
rect 166408 329372 166414 329384
rect 166902 329372 166908 329384
rect 166408 329344 166908 329372
rect 166408 329332 166414 329344
rect 166902 329332 166908 329344
rect 166960 329332 166966 329384
rect 115198 329128 115204 329180
rect 115256 329168 115262 329180
rect 115842 329168 115848 329180
rect 115256 329140 115848 329168
rect 115256 329128 115262 329140
rect 115842 329128 115848 329140
rect 115900 329128 115906 329180
rect 115842 328516 115848 328568
rect 115900 328556 115906 328568
rect 192570 328556 192576 328568
rect 115900 328528 192576 328556
rect 115900 328516 115906 328528
rect 192570 328516 192576 328528
rect 192628 328516 192634 328568
rect 166350 328448 166356 328500
rect 166408 328488 166414 328500
rect 256786 328488 256792 328500
rect 166408 328460 256792 328488
rect 166408 328448 166414 328460
rect 256786 328448 256792 328460
rect 256844 328448 256850 328500
rect 242802 328040 242808 328092
rect 242860 328080 242866 328092
rect 244366 328080 244372 328092
rect 242860 328052 244372 328080
rect 242860 328040 242866 328052
rect 244366 328040 244372 328052
rect 244424 328040 244430 328092
rect 253842 327768 253848 327820
rect 253900 327808 253906 327820
rect 265250 327808 265256 327820
rect 253900 327780 265256 327808
rect 253900 327768 253906 327780
rect 265250 327768 265256 327780
rect 265308 327768 265314 327820
rect 181990 327700 181996 327752
rect 182048 327740 182054 327752
rect 192478 327740 192484 327752
rect 182048 327712 192484 327740
rect 182048 327700 182054 327712
rect 192478 327700 192484 327712
rect 192536 327700 192542 327752
rect 141694 327088 141700 327140
rect 141752 327128 141758 327140
rect 189074 327128 189080 327140
rect 141752 327100 189080 327128
rect 141752 327088 141758 327100
rect 189074 327088 189080 327100
rect 189132 327088 189138 327140
rect 170398 326340 170404 326392
rect 170456 326380 170462 326392
rect 184198 326380 184204 326392
rect 170456 326352 184204 326380
rect 170456 326340 170462 326352
rect 184198 326340 184204 326352
rect 184256 326340 184262 326392
rect 188338 326340 188344 326392
rect 188396 326380 188402 326392
rect 227070 326380 227076 326392
rect 188396 326352 227076 326380
rect 188396 326340 188402 326352
rect 227070 326340 227076 326352
rect 227128 326340 227134 326392
rect 236638 326340 236644 326392
rect 236696 326380 236702 326392
rect 259822 326380 259828 326392
rect 236696 326352 259828 326380
rect 236696 326340 236702 326352
rect 259822 326340 259828 326352
rect 259880 326340 259886 326392
rect 261478 326340 261484 326392
rect 261536 326380 261542 326392
rect 283098 326380 283104 326392
rect 261536 326352 283104 326380
rect 261536 326340 261542 326352
rect 283098 326340 283104 326352
rect 283156 326340 283162 326392
rect 163590 325660 163596 325712
rect 163648 325700 163654 325712
rect 242986 325700 242992 325712
rect 163648 325672 242992 325700
rect 163648 325660 163654 325672
rect 242986 325660 242992 325672
rect 243044 325660 243050 325712
rect 239398 324912 239404 324964
rect 239456 324952 239462 324964
rect 249794 324952 249800 324964
rect 239456 324924 249800 324952
rect 239456 324912 239462 324924
rect 249794 324912 249800 324924
rect 249852 324912 249858 324964
rect 159358 324300 159364 324352
rect 159416 324340 159422 324352
rect 259730 324340 259736 324352
rect 159416 324312 259736 324340
rect 159416 324300 159422 324312
rect 259730 324300 259736 324312
rect 259788 324300 259794 324352
rect 144270 323620 144276 323672
rect 144328 323660 144334 323672
rect 159358 323660 159364 323672
rect 144328 323632 159364 323660
rect 144328 323620 144334 323632
rect 159358 323620 159364 323632
rect 159416 323620 159422 323672
rect 162394 323620 162400 323672
rect 162452 323660 162458 323672
rect 259454 323660 259460 323672
rect 162452 323632 259460 323660
rect 162452 323620 162458 323632
rect 259454 323620 259460 323632
rect 259512 323620 259518 323672
rect 108390 323552 108396 323604
rect 108448 323592 108454 323604
rect 120718 323592 120724 323604
rect 108448 323564 120724 323592
rect 108448 323552 108454 323564
rect 120718 323552 120724 323564
rect 120776 323592 120782 323604
rect 273530 323592 273536 323604
rect 120776 323564 273536 323592
rect 120776 323552 120782 323564
rect 273530 323552 273536 323564
rect 273588 323552 273594 323604
rect 125686 322872 125692 322924
rect 125744 322912 125750 322924
rect 276106 322912 276112 322924
rect 125744 322884 276112 322912
rect 125744 322872 125750 322884
rect 276106 322872 276112 322884
rect 276164 322872 276170 322924
rect 104250 322260 104256 322312
rect 104308 322300 104314 322312
rect 125686 322300 125692 322312
rect 104308 322272 125692 322300
rect 104308 322260 104314 322272
rect 125686 322260 125692 322272
rect 125744 322260 125750 322312
rect 86218 322192 86224 322244
rect 86276 322232 86282 322244
rect 166258 322232 166264 322244
rect 86276 322204 166264 322232
rect 86276 322192 86282 322204
rect 166258 322192 166264 322204
rect 166316 322232 166322 322244
rect 258074 322232 258080 322244
rect 166316 322204 258080 322232
rect 166316 322192 166322 322204
rect 258074 322192 258080 322204
rect 258132 322192 258138 322244
rect 193122 320900 193128 320952
rect 193180 320940 193186 320952
rect 216674 320940 216680 320952
rect 193180 320912 216680 320940
rect 193180 320900 193186 320912
rect 216674 320900 216680 320912
rect 216732 320900 216738 320952
rect 226978 320900 226984 320952
rect 227036 320940 227042 320952
rect 262398 320940 262404 320952
rect 227036 320912 262404 320940
rect 227036 320900 227042 320912
rect 262398 320900 262404 320912
rect 262456 320900 262462 320952
rect 126882 320832 126888 320884
rect 126940 320872 126946 320884
rect 136634 320872 136640 320884
rect 126940 320844 136640 320872
rect 126940 320832 126946 320844
rect 136634 320832 136640 320844
rect 136692 320872 136698 320884
rect 263594 320872 263600 320884
rect 136692 320844 263600 320872
rect 136692 320832 136698 320844
rect 263594 320832 263600 320844
rect 263652 320832 263658 320884
rect 268378 320832 268384 320884
rect 268436 320872 268442 320884
rect 286410 320872 286416 320884
rect 268436 320844 286416 320872
rect 268436 320832 268442 320844
rect 286410 320832 286416 320844
rect 286468 320832 286474 320884
rect 104342 320220 104348 320272
rect 104400 320260 104406 320272
rect 126882 320260 126888 320272
rect 104400 320232 126888 320260
rect 104400 320220 104406 320232
rect 126882 320220 126888 320232
rect 126940 320220 126946 320272
rect 75822 320152 75828 320204
rect 75880 320192 75886 320204
rect 108298 320192 108304 320204
rect 75880 320164 108304 320192
rect 75880 320152 75886 320164
rect 108298 320152 108304 320164
rect 108356 320152 108362 320204
rect 175918 319472 175924 319524
rect 175976 319512 175982 319524
rect 176562 319512 176568 319524
rect 175976 319484 176568 319512
rect 175976 319472 175982 319484
rect 176562 319472 176568 319484
rect 176620 319472 176626 319524
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 15838 319444 15844 319456
rect 4120 319416 15844 319444
rect 4120 319404 4126 319416
rect 15838 319404 15844 319416
rect 15896 319404 15902 319456
rect 97994 319404 98000 319456
rect 98052 319444 98058 319456
rect 141418 319444 141424 319456
rect 98052 319416 141424 319444
rect 98052 319404 98058 319416
rect 141418 319404 141424 319416
rect 141476 319404 141482 319456
rect 182082 319404 182088 319456
rect 182140 319444 182146 319456
rect 215294 319444 215300 319456
rect 182140 319416 215300 319444
rect 182140 319404 182146 319416
rect 215294 319404 215300 319416
rect 215352 319404 215358 319456
rect 233970 319404 233976 319456
rect 234028 319444 234034 319456
rect 276198 319444 276204 319456
rect 234028 319416 276204 319444
rect 234028 319404 234034 319416
rect 276198 319404 276204 319416
rect 276256 319404 276262 319456
rect 259362 319336 259368 319388
rect 259420 319376 259426 319388
rect 263778 319376 263784 319388
rect 259420 319348 263784 319376
rect 259420 319336 259426 319348
rect 263778 319336 263784 319348
rect 263836 319336 263842 319388
rect 175918 318792 175924 318844
rect 175976 318832 175982 318844
rect 246482 318832 246488 318844
rect 175976 318804 246488 318832
rect 175976 318792 175982 318804
rect 246482 318792 246488 318804
rect 246540 318792 246546 318844
rect 71958 318044 71964 318096
rect 72016 318084 72022 318096
rect 88978 318084 88984 318096
rect 72016 318056 88984 318084
rect 72016 318044 72022 318056
rect 88978 318044 88984 318056
rect 89036 318044 89042 318096
rect 103422 318044 103428 318096
rect 103480 318084 103486 318096
rect 114554 318084 114560 318096
rect 103480 318056 114560 318084
rect 103480 318044 103486 318056
rect 114554 318044 114560 318056
rect 114612 318044 114618 318096
rect 144822 317500 144828 317552
rect 144880 317540 144886 317552
rect 197446 317540 197452 317552
rect 144880 317512 197452 317540
rect 144880 317500 144886 317512
rect 197446 317500 197452 317512
rect 197504 317500 197510 317552
rect 142798 317432 142804 317484
rect 142856 317472 142862 317484
rect 261018 317472 261024 317484
rect 142856 317444 261024 317472
rect 142856 317432 142862 317444
rect 261018 317432 261024 317444
rect 261076 317432 261082 317484
rect 184198 317364 184204 317416
rect 184256 317404 184262 317416
rect 184658 317404 184664 317416
rect 184256 317376 184664 317404
rect 184256 317364 184262 317376
rect 184658 317364 184664 317376
rect 184716 317364 184722 317416
rect 214006 316752 214012 316804
rect 214064 316792 214070 316804
rect 214558 316792 214564 316804
rect 214064 316764 214564 316792
rect 214064 316752 214070 316764
rect 214558 316752 214564 316764
rect 214616 316752 214622 316804
rect 119338 316684 119344 316736
rect 119396 316724 119402 316736
rect 190454 316724 190460 316736
rect 119396 316696 190460 316724
rect 119396 316684 119402 316696
rect 190454 316684 190460 316696
rect 190512 316684 190518 316736
rect 215294 316684 215300 316736
rect 215352 316724 215358 316736
rect 254670 316724 254676 316736
rect 215352 316696 254676 316724
rect 215352 316684 215358 316696
rect 254670 316684 254676 316696
rect 254728 316724 254734 316736
rect 579614 316724 579620 316736
rect 254728 316696 579620 316724
rect 254728 316684 254734 316696
rect 579614 316684 579620 316696
rect 579672 316684 579678 316736
rect 87598 316616 87604 316668
rect 87656 316656 87662 316668
rect 88242 316656 88248 316668
rect 87656 316628 88248 316656
rect 87656 316616 87662 316628
rect 88242 316616 88248 316628
rect 88300 316616 88306 316668
rect 192478 316072 192484 316124
rect 192536 316112 192542 316124
rect 214558 316112 214564 316124
rect 192536 316084 214564 316112
rect 192536 316072 192542 316084
rect 214558 316072 214564 316084
rect 214616 316072 214622 316124
rect 88242 316004 88248 316056
rect 88300 316044 88306 316056
rect 110506 316044 110512 316056
rect 88300 316016 110512 316044
rect 88300 316004 88306 316016
rect 110506 316004 110512 316016
rect 110564 316004 110570 316056
rect 184658 316004 184664 316056
rect 184716 316044 184722 316056
rect 257338 316044 257344 316056
rect 184716 316016 257344 316044
rect 184716 316004 184722 316016
rect 257338 316004 257344 316016
rect 257396 316004 257402 316056
rect 228358 315256 228364 315308
rect 228416 315296 228422 315308
rect 265066 315296 265072 315308
rect 228416 315268 265072 315296
rect 228416 315256 228422 315268
rect 265066 315256 265072 315268
rect 265124 315256 265130 315308
rect 190454 315188 190460 315240
rect 190512 315228 190518 315240
rect 191558 315228 191564 315240
rect 190512 315200 191564 315228
rect 190512 315188 190518 315200
rect 191558 315188 191564 315200
rect 191616 315228 191622 315240
rect 195238 315228 195244 315240
rect 191616 315200 195244 315228
rect 191616 315188 191622 315200
rect 195238 315188 195244 315200
rect 195296 315188 195302 315240
rect 178678 314644 178684 314696
rect 178736 314684 178742 314696
rect 179322 314684 179328 314696
rect 178736 314656 179328 314684
rect 178736 314644 178742 314656
rect 179322 314644 179328 314656
rect 179380 314684 179386 314696
rect 226334 314684 226340 314696
rect 179380 314656 226340 314684
rect 179380 314644 179386 314656
rect 226334 314644 226340 314656
rect 226392 314644 226398 314696
rect 216030 313896 216036 313948
rect 216088 313936 216094 313948
rect 236546 313936 236552 313948
rect 216088 313908 236552 313936
rect 216088 313896 216094 313908
rect 236546 313896 236552 313908
rect 236604 313896 236610 313948
rect 239398 313896 239404 313948
rect 239456 313936 239462 313948
rect 269390 313936 269396 313948
rect 239456 313908 269396 313936
rect 239456 313896 239462 313908
rect 269390 313896 269396 313908
rect 269448 313896 269454 313948
rect 167638 313352 167644 313404
rect 167696 313392 167702 313404
rect 208394 313392 208400 313404
rect 167696 313364 208400 313392
rect 167696 313352 167702 313364
rect 208394 313352 208400 313364
rect 208452 313352 208458 313404
rect 164878 313284 164884 313336
rect 164936 313324 164942 313336
rect 211338 313324 211344 313336
rect 164936 313296 211344 313324
rect 164936 313284 164942 313296
rect 211338 313284 211344 313296
rect 211396 313284 211402 313336
rect 238662 313284 238668 313336
rect 238720 313324 238726 313336
rect 279050 313324 279056 313336
rect 238720 313296 279056 313324
rect 238720 313284 238726 313296
rect 279050 313284 279056 313296
rect 279108 313284 279114 313336
rect 246482 312536 246488 312588
rect 246540 312576 246546 312588
rect 273254 312576 273260 312588
rect 246540 312548 273260 312576
rect 246540 312536 246546 312548
rect 273254 312536 273260 312548
rect 273312 312536 273318 312588
rect 185578 311924 185584 311976
rect 185636 311964 185642 311976
rect 186130 311964 186136 311976
rect 185636 311936 186136 311964
rect 185636 311924 185642 311936
rect 186130 311924 186136 311936
rect 186188 311964 186194 311976
rect 262490 311964 262496 311976
rect 186188 311936 262496 311964
rect 186188 311924 186194 311936
rect 262490 311924 262496 311936
rect 262548 311924 262554 311976
rect 151262 311856 151268 311908
rect 151320 311896 151326 311908
rect 231854 311896 231860 311908
rect 151320 311868 231860 311896
rect 151320 311856 151326 311868
rect 231854 311856 231860 311868
rect 231912 311856 231918 311908
rect 218054 311108 218060 311160
rect 218112 311148 218118 311160
rect 249610 311148 249616 311160
rect 218112 311120 249616 311148
rect 218112 311108 218118 311120
rect 249610 311108 249616 311120
rect 249668 311108 249674 311160
rect 181438 310564 181444 310616
rect 181496 310604 181502 310616
rect 267734 310604 267740 310616
rect 181496 310576 267740 310604
rect 181496 310564 181502 310576
rect 267734 310564 267740 310576
rect 267792 310564 267798 310616
rect 115842 310496 115848 310548
rect 115900 310536 115906 310548
rect 217410 310536 217416 310548
rect 115900 310508 217416 310536
rect 115900 310496 115906 310508
rect 217410 310496 217416 310508
rect 217468 310496 217474 310548
rect 57606 310428 57612 310480
rect 57664 310468 57670 310480
rect 57882 310468 57888 310480
rect 57664 310440 57888 310468
rect 57664 310428 57670 310440
rect 57882 310428 57888 310440
rect 57940 310428 57946 310480
rect 112530 310428 112536 310480
rect 112588 310468 112594 310480
rect 114646 310468 114652 310480
rect 112588 310440 114652 310468
rect 112588 310428 112594 310440
rect 114646 310428 114652 310440
rect 114704 310428 114710 310480
rect 168374 310428 168380 310480
rect 168432 310468 168438 310480
rect 169018 310468 169024 310480
rect 168432 310440 169024 310468
rect 168432 310428 168438 310440
rect 169018 310428 169024 310440
rect 169076 310428 169082 310480
rect 57514 309884 57520 309936
rect 57572 309924 57578 309936
rect 80054 309924 80060 309936
rect 57572 309896 80060 309924
rect 57572 309884 57578 309896
rect 80054 309884 80060 309896
rect 80112 309884 80118 309936
rect 57882 309748 57888 309800
rect 57940 309788 57946 309800
rect 168374 309788 168380 309800
rect 57940 309760 168380 309788
rect 57940 309748 57946 309760
rect 168374 309748 168380 309760
rect 168432 309748 168438 309800
rect 187050 309204 187056 309256
rect 187108 309244 187114 309256
rect 259546 309244 259552 309256
rect 187108 309216 259552 309244
rect 187108 309204 187114 309216
rect 259546 309204 259552 309216
rect 259604 309204 259610 309256
rect 170398 309136 170404 309188
rect 170456 309176 170462 309188
rect 271874 309176 271880 309188
rect 170456 309148 271880 309176
rect 170456 309136 170462 309148
rect 271874 309136 271880 309148
rect 271932 309136 271938 309188
rect 184566 309068 184572 309120
rect 184624 309108 184630 309120
rect 187694 309108 187700 309120
rect 184624 309080 187700 309108
rect 184624 309068 184630 309080
rect 187694 309068 187700 309080
rect 187752 309068 187758 309120
rect 84194 308388 84200 308440
rect 84252 308428 84258 308440
rect 151170 308428 151176 308440
rect 84252 308400 151176 308428
rect 84252 308388 84258 308400
rect 151170 308388 151176 308400
rect 151228 308388 151234 308440
rect 223574 308388 223580 308440
rect 223632 308428 223638 308440
rect 255958 308428 255964 308440
rect 223632 308400 255964 308428
rect 223632 308388 223638 308400
rect 255958 308388 255964 308400
rect 256016 308388 256022 308440
rect 4062 307776 4068 307828
rect 4120 307816 4126 307828
rect 7558 307816 7564 307828
rect 4120 307788 7564 307816
rect 4120 307776 4126 307788
rect 7558 307776 7564 307788
rect 7616 307776 7622 307828
rect 148318 307776 148324 307828
rect 148376 307816 148382 307828
rect 216030 307816 216036 307828
rect 148376 307788 216036 307816
rect 148376 307776 148382 307788
rect 216030 307776 216036 307788
rect 216088 307776 216094 307828
rect 251818 307776 251824 307828
rect 251876 307816 251882 307828
rect 282914 307816 282920 307828
rect 251876 307788 282920 307816
rect 251876 307776 251882 307788
rect 282914 307776 282920 307788
rect 282972 307776 282978 307828
rect 233234 307096 233240 307148
rect 233292 307136 233298 307148
rect 252554 307136 252560 307148
rect 233292 307108 252560 307136
rect 233292 307096 233298 307108
rect 252554 307096 252560 307108
rect 252612 307096 252618 307148
rect 199378 307028 199384 307080
rect 199436 307068 199442 307080
rect 203978 307068 203984 307080
rect 199436 307040 203984 307068
rect 199436 307028 199442 307040
rect 203978 307028 203984 307040
rect 204036 307028 204042 307080
rect 226334 307028 226340 307080
rect 226392 307068 226398 307080
rect 262306 307068 262312 307080
rect 226392 307040 262312 307068
rect 226392 307028 226398 307040
rect 262306 307028 262312 307040
rect 262364 307028 262370 307080
rect 253198 306552 253204 306604
rect 253256 306592 253262 306604
rect 258258 306592 258264 306604
rect 253256 306564 258264 306592
rect 253256 306552 253262 306564
rect 258258 306552 258264 306564
rect 258316 306552 258322 306604
rect 152458 306416 152464 306468
rect 152516 306456 152522 306468
rect 214190 306456 214196 306468
rect 152516 306428 214196 306456
rect 152516 306416 152522 306428
rect 214190 306416 214196 306428
rect 214248 306416 214254 306468
rect 9582 306348 9588 306400
rect 9640 306388 9646 306400
rect 197354 306388 197360 306400
rect 9640 306360 197360 306388
rect 9640 306348 9646 306360
rect 197354 306348 197360 306360
rect 197412 306348 197418 306400
rect 213270 305736 213276 305788
rect 213328 305776 213334 305788
rect 231578 305776 231584 305788
rect 213328 305748 231584 305776
rect 213328 305736 213334 305748
rect 231578 305736 231584 305748
rect 231636 305736 231642 305788
rect 222838 305600 222844 305652
rect 222896 305640 222902 305652
rect 246022 305640 246028 305652
rect 222896 305612 246028 305640
rect 222896 305600 222902 305612
rect 246022 305600 246028 305612
rect 246080 305600 246086 305652
rect 191374 305056 191380 305108
rect 191432 305096 191438 305108
rect 193306 305096 193312 305108
rect 191432 305068 193312 305096
rect 191432 305056 191438 305068
rect 193306 305056 193312 305068
rect 193364 305056 193370 305108
rect 193490 305056 193496 305108
rect 193548 305096 193554 305108
rect 202782 305096 202788 305108
rect 193548 305068 202788 305096
rect 193548 305056 193554 305068
rect 202782 305056 202788 305068
rect 202840 305056 202846 305108
rect 249242 305056 249248 305108
rect 249300 305096 249306 305108
rect 249702 305096 249708 305108
rect 249300 305068 249708 305096
rect 249300 305056 249306 305068
rect 249702 305056 249708 305068
rect 249760 305096 249766 305108
rect 278774 305096 278780 305108
rect 249760 305068 278780 305096
rect 249760 305056 249766 305068
rect 278774 305056 278780 305068
rect 278832 305056 278838 305108
rect 137278 304988 137284 305040
rect 137336 305028 137342 305040
rect 216582 305028 216588 305040
rect 137336 305000 216588 305028
rect 137336 304988 137342 305000
rect 216582 304988 216588 305000
rect 216640 304988 216646 305040
rect 240042 304988 240048 305040
rect 240100 305028 240106 305040
rect 270678 305028 270684 305040
rect 240100 305000 270684 305028
rect 240100 304988 240106 305000
rect 270678 304988 270684 305000
rect 270736 304988 270742 305040
rect 218698 304920 218704 304972
rect 218756 304960 218762 304972
rect 220814 304960 220820 304972
rect 218756 304932 220820 304960
rect 218756 304920 218762 304932
rect 220814 304920 220820 304932
rect 220872 304920 220878 304972
rect 97902 304308 97908 304360
rect 97960 304348 97966 304360
rect 108390 304348 108396 304360
rect 97960 304320 108396 304348
rect 97960 304308 97966 304320
rect 108390 304308 108396 304320
rect 108448 304308 108454 304360
rect 123478 304308 123484 304360
rect 123536 304348 123542 304360
rect 151078 304348 151084 304360
rect 123536 304320 151084 304348
rect 123536 304308 123542 304320
rect 151078 304308 151084 304320
rect 151136 304308 151142 304360
rect 151354 304308 151360 304360
rect 151412 304348 151418 304360
rect 164878 304348 164884 304360
rect 151412 304320 164884 304348
rect 151412 304308 151418 304320
rect 164878 304308 164884 304320
rect 164936 304308 164942 304360
rect 226978 304308 226984 304360
rect 227036 304348 227042 304360
rect 236362 304348 236368 304360
rect 227036 304320 236368 304348
rect 227036 304308 227042 304320
rect 236362 304308 236368 304320
rect 236420 304308 236426 304360
rect 60458 304240 60464 304292
rect 60516 304280 60522 304292
rect 170490 304280 170496 304292
rect 60516 304252 170496 304280
rect 60516 304240 60522 304252
rect 170490 304240 170496 304252
rect 170548 304240 170554 304292
rect 213178 304240 213184 304292
rect 213236 304280 213242 304292
rect 223206 304280 223212 304292
rect 213236 304252 223212 304280
rect 213236 304240 213242 304252
rect 223206 304240 223212 304252
rect 223264 304240 223270 304292
rect 231118 304240 231124 304292
rect 231176 304280 231182 304292
rect 253198 304280 253204 304292
rect 231176 304252 253204 304280
rect 231176 304240 231182 304252
rect 253198 304240 253204 304252
rect 253256 304240 253262 304292
rect 226518 303764 226524 303816
rect 226576 303804 226582 303816
rect 231026 303804 231032 303816
rect 226576 303776 231032 303804
rect 226576 303764 226582 303776
rect 231026 303764 231032 303776
rect 231084 303764 231090 303816
rect 186038 303696 186044 303748
rect 186096 303736 186102 303748
rect 196250 303736 196256 303748
rect 186096 303708 196256 303736
rect 186096 303696 186102 303708
rect 196250 303696 196256 303708
rect 196308 303696 196314 303748
rect 221458 303696 221464 303748
rect 221516 303736 221522 303748
rect 224402 303736 224408 303748
rect 221516 303708 224408 303736
rect 221516 303696 221522 303708
rect 224402 303696 224408 303708
rect 224460 303696 224466 303748
rect 193214 303628 193220 303680
rect 193272 303668 193278 303680
rect 193582 303668 193588 303680
rect 193272 303640 193588 303668
rect 193272 303628 193278 303640
rect 193582 303628 193588 303640
rect 193640 303628 193646 303680
rect 211338 303628 211344 303680
rect 211396 303668 211402 303680
rect 212166 303668 212172 303680
rect 211396 303640 212172 303668
rect 211396 303628 211402 303640
rect 212166 303628 212172 303640
rect 212224 303628 212230 303680
rect 215938 303628 215944 303680
rect 215996 303668 216002 303680
rect 217226 303668 217232 303680
rect 215996 303640 217232 303668
rect 215996 303628 216002 303640
rect 217226 303628 217232 303640
rect 217284 303628 217290 303680
rect 220906 303628 220912 303680
rect 220964 303668 220970 303680
rect 221734 303668 221740 303680
rect 220964 303640 221740 303668
rect 220964 303628 220970 303640
rect 221734 303628 221740 303640
rect 221792 303628 221798 303680
rect 222930 303628 222936 303680
rect 222988 303668 222994 303680
rect 226242 303668 226248 303680
rect 222988 303640 226248 303668
rect 222988 303628 222994 303640
rect 226242 303628 226248 303640
rect 226300 303628 226306 303680
rect 243078 303628 243084 303680
rect 243136 303668 243142 303680
rect 243814 303668 243820 303680
rect 243136 303640 243820 303668
rect 243136 303628 243142 303640
rect 243814 303628 243820 303640
rect 243872 303628 243878 303680
rect 248414 303628 248420 303680
rect 248472 303668 248478 303680
rect 248966 303668 248972 303680
rect 248472 303640 248972 303668
rect 248472 303628 248478 303640
rect 248966 303628 248972 303640
rect 249024 303668 249030 303680
rect 265158 303668 265164 303680
rect 249024 303640 265164 303668
rect 249024 303628 249030 303640
rect 265158 303628 265164 303640
rect 265216 303628 265222 303680
rect 176654 302880 176660 302932
rect 176712 302920 176718 302932
rect 177390 302920 177396 302932
rect 176712 302892 177396 302920
rect 176712 302880 176718 302892
rect 177390 302880 177396 302892
rect 177448 302920 177454 302932
rect 192662 302920 192668 302932
rect 177448 302892 192668 302920
rect 177448 302880 177454 302892
rect 192662 302880 192668 302892
rect 192720 302880 192726 302932
rect 197354 302880 197360 302932
rect 197412 302920 197418 302932
rect 211246 302920 211252 302932
rect 197412 302892 211252 302920
rect 197412 302880 197418 302892
rect 211246 302880 211252 302892
rect 211304 302880 211310 302932
rect 233142 302880 233148 302932
rect 233200 302920 233206 302932
rect 254118 302920 254124 302932
rect 233200 302892 254124 302920
rect 233200 302880 233206 302892
rect 254118 302880 254124 302892
rect 254176 302880 254182 302932
rect 257430 302880 257436 302932
rect 257488 302920 257494 302932
rect 261110 302920 261116 302932
rect 257488 302892 261116 302920
rect 257488 302880 257494 302892
rect 261110 302880 261116 302892
rect 261168 302880 261174 302932
rect 87690 302268 87696 302320
rect 87748 302308 87754 302320
rect 176654 302308 176660 302320
rect 87748 302280 176660 302308
rect 87748 302268 87754 302280
rect 176654 302268 176660 302280
rect 176712 302268 176718 302320
rect 192570 302268 192576 302320
rect 192628 302308 192634 302320
rect 218422 302308 218428 302320
rect 192628 302280 218428 302308
rect 192628 302268 192634 302280
rect 218422 302268 218428 302280
rect 218480 302268 218486 302320
rect 15838 302200 15844 302252
rect 15896 302240 15902 302252
rect 197998 302240 198004 302252
rect 15896 302212 198004 302240
rect 15896 302200 15902 302212
rect 197998 302200 198004 302212
rect 198056 302200 198062 302252
rect 247678 302200 247684 302252
rect 247736 302240 247742 302252
rect 281534 302240 281540 302252
rect 247736 302212 281540 302240
rect 247736 302200 247742 302212
rect 281534 302200 281540 302212
rect 281592 302200 281598 302252
rect 252462 302132 252468 302184
rect 252520 302172 252526 302184
rect 258442 302172 258448 302184
rect 252520 302144 258448 302172
rect 252520 302132 252526 302144
rect 258442 302132 258448 302144
rect 258500 302132 258506 302184
rect 240870 301656 240876 301708
rect 240928 301656 240934 301708
rect 73062 301452 73068 301504
rect 73120 301492 73126 301504
rect 173618 301492 173624 301504
rect 73120 301464 173624 301492
rect 73120 301452 73126 301464
rect 173618 301452 173624 301464
rect 173676 301492 173682 301504
rect 176102 301492 176108 301504
rect 173676 301464 176108 301492
rect 173676 301452 173682 301464
rect 176102 301452 176108 301464
rect 176160 301452 176166 301504
rect 240888 301492 240916 301656
rect 252922 301492 252928 301504
rect 240888 301464 252928 301492
rect 252922 301452 252928 301464
rect 252980 301452 252986 301504
rect 193306 301044 193312 301096
rect 193364 301084 193370 301096
rect 195238 301084 195244 301096
rect 193364 301056 195244 301084
rect 193364 301044 193370 301056
rect 195238 301044 195244 301056
rect 195296 301044 195302 301096
rect 245102 301084 245108 301096
rect 238726 301056 245108 301084
rect 188522 300976 188528 301028
rect 188580 301016 188586 301028
rect 206922 301016 206928 301028
rect 188580 300988 206928 301016
rect 188580 300976 188586 300988
rect 206922 300976 206928 300988
rect 206980 300976 206986 301028
rect 178862 300908 178868 300960
rect 178920 300948 178926 300960
rect 192478 300948 192484 300960
rect 178920 300920 192484 300948
rect 178920 300908 178926 300920
rect 192478 300908 192484 300920
rect 192536 300908 192542 300960
rect 199470 300908 199476 300960
rect 199528 300908 199534 300960
rect 214558 300908 214564 300960
rect 214616 300908 214622 300960
rect 191466 300772 191472 300824
rect 191524 300812 191530 300824
rect 199488 300812 199516 300908
rect 214576 300880 214604 300908
rect 238726 300880 238754 301056
rect 245102 301044 245108 301056
rect 245160 301044 245166 301096
rect 242066 300976 242072 301028
rect 242124 300976 242130 301028
rect 214576 300852 238754 300880
rect 191524 300784 199516 300812
rect 242084 300812 242112 300976
rect 258718 300908 258724 300960
rect 258776 300948 258782 300960
rect 259454 300948 259460 300960
rect 258776 300920 259460 300948
rect 258776 300908 258782 300920
rect 259454 300908 259460 300920
rect 259512 300908 259518 300960
rect 255406 300840 255412 300892
rect 255464 300880 255470 300892
rect 278038 300880 278044 300892
rect 255464 300852 278044 300880
rect 255464 300840 255470 300852
rect 278038 300840 278044 300852
rect 278096 300840 278102 300892
rect 252462 300812 252468 300824
rect 242084 300784 252468 300812
rect 191524 300772 191530 300784
rect 252462 300772 252468 300784
rect 252520 300772 252526 300824
rect 124950 300092 124956 300144
rect 125008 300132 125014 300144
rect 159450 300132 159456 300144
rect 125008 300104 159456 300132
rect 125008 300092 125014 300104
rect 159450 300092 159456 300104
rect 159508 300132 159514 300144
rect 164234 300132 164240 300144
rect 159508 300104 164240 300132
rect 159508 300092 159514 300104
rect 164234 300092 164240 300104
rect 164292 300092 164298 300144
rect 255774 299548 255780 299600
rect 255832 299588 255838 299600
rect 259362 299588 259368 299600
rect 255832 299560 259368 299588
rect 255832 299548 255838 299560
rect 259362 299548 259368 299560
rect 259420 299548 259426 299600
rect 164234 299480 164240 299532
rect 164292 299520 164298 299532
rect 191742 299520 191748 299532
rect 164292 299492 191748 299520
rect 164292 299480 164298 299492
rect 191742 299480 191748 299492
rect 191800 299480 191806 299532
rect 255406 299480 255412 299532
rect 255464 299520 255470 299532
rect 288710 299520 288716 299532
rect 255464 299492 288716 299520
rect 255464 299480 255470 299492
rect 288710 299480 288716 299492
rect 288768 299480 288774 299532
rect 281350 299412 281356 299464
rect 281408 299452 281414 299464
rect 580166 299452 580172 299464
rect 281408 299424 580172 299452
rect 281408 299412 281414 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 191006 298840 191012 298852
rect 190426 298812 191012 298840
rect 92842 298732 92848 298784
rect 92900 298772 92906 298784
rect 130470 298772 130476 298784
rect 92900 298744 130476 298772
rect 92900 298732 92906 298744
rect 130470 298732 130476 298744
rect 130528 298732 130534 298784
rect 170490 298732 170496 298784
rect 170548 298772 170554 298784
rect 187510 298772 187516 298784
rect 170548 298744 187516 298772
rect 170548 298732 170554 298744
rect 187510 298732 187516 298744
rect 187568 298772 187574 298784
rect 190426 298772 190454 298812
rect 191006 298800 191012 298812
rect 191064 298800 191070 298852
rect 275278 298800 275284 298852
rect 275336 298840 275342 298852
rect 280246 298840 280252 298852
rect 275336 298812 280252 298840
rect 275336 298800 275342 298812
rect 280246 298800 280252 298812
rect 280304 298840 280310 298852
rect 281350 298840 281356 298852
rect 280304 298812 281356 298840
rect 280304 298800 280310 298812
rect 281350 298800 281356 298812
rect 281408 298800 281414 298852
rect 187568 298744 190454 298772
rect 187568 298732 187574 298744
rect 259362 298732 259368 298784
rect 259420 298772 259426 298784
rect 293954 298772 293960 298784
rect 259420 298744 293960 298772
rect 259420 298732 259426 298744
rect 293954 298732 293960 298744
rect 294012 298732 294018 298784
rect 257338 298188 257344 298240
rect 257396 298228 257402 298240
rect 258166 298228 258172 298240
rect 257396 298200 258172 298228
rect 257396 298188 257402 298200
rect 258166 298188 258172 298200
rect 258224 298188 258230 298240
rect 255406 298120 255412 298172
rect 255464 298160 255470 298172
rect 266630 298160 266636 298172
rect 255464 298132 266636 298160
rect 255464 298120 255470 298132
rect 266630 298120 266636 298132
rect 266688 298120 266694 298172
rect 164142 298052 164148 298104
rect 164200 298092 164206 298104
rect 191742 298092 191748 298104
rect 164200 298064 191748 298092
rect 164200 298052 164206 298064
rect 191742 298052 191748 298064
rect 191800 298052 191806 298104
rect 255406 297712 255412 297764
rect 255464 297752 255470 297764
rect 259454 297752 259460 297764
rect 255464 297724 259460 297752
rect 255464 297712 255470 297724
rect 259454 297712 259460 297724
rect 259512 297712 259518 297764
rect 91186 297372 91192 297424
rect 91244 297412 91250 297424
rect 104342 297412 104348 297424
rect 91244 297384 104348 297412
rect 91244 297372 91250 297384
rect 104342 297372 104348 297384
rect 104400 297372 104406 297424
rect 117222 297372 117228 297424
rect 117280 297412 117286 297424
rect 164142 297412 164148 297424
rect 117280 297384 164148 297412
rect 117280 297372 117286 297384
rect 164142 297372 164148 297384
rect 164200 297372 164206 297424
rect 253290 296692 253296 296744
rect 253348 296732 253354 296744
rect 296714 296732 296720 296744
rect 253348 296704 296720 296732
rect 253348 296692 253354 296704
rect 296714 296692 296720 296704
rect 296772 296692 296778 296744
rect 255498 296080 255504 296132
rect 255556 296120 255562 296132
rect 255682 296120 255688 296132
rect 255556 296092 255688 296120
rect 255556 296080 255562 296092
rect 255682 296080 255688 296092
rect 255740 296080 255746 296132
rect 130562 296012 130568 296064
rect 130620 296052 130626 296064
rect 191558 296052 191564 296064
rect 130620 296024 191564 296052
rect 130620 296012 130626 296024
rect 191558 296012 191564 296024
rect 191616 296012 191622 296064
rect 78582 295944 78588 295996
rect 78640 295984 78646 295996
rect 78640 295956 180794 295984
rect 78640 295944 78646 295956
rect 180766 295916 180794 295956
rect 255498 295944 255504 295996
rect 255556 295984 255562 295996
rect 265250 295984 265256 295996
rect 255556 295956 265256 295984
rect 255556 295944 255562 295956
rect 265250 295944 265256 295956
rect 265308 295984 265314 295996
rect 284478 295984 284484 295996
rect 265308 295956 284484 295984
rect 265308 295944 265314 295956
rect 284478 295944 284484 295956
rect 284536 295944 284542 295996
rect 189074 295916 189080 295928
rect 180766 295888 189080 295916
rect 189074 295876 189080 295888
rect 189132 295916 189138 295928
rect 189718 295916 189724 295928
rect 189132 295888 189724 295916
rect 189132 295876 189138 295888
rect 189718 295876 189724 295888
rect 189776 295876 189782 295928
rect 77386 295332 77392 295384
rect 77444 295372 77450 295384
rect 78582 295372 78588 295384
rect 77444 295344 78588 295372
rect 77444 295332 77450 295344
rect 78582 295332 78588 295344
rect 78640 295332 78646 295384
rect 191282 295332 191288 295384
rect 191340 295372 191346 295384
rect 193398 295372 193404 295384
rect 191340 295344 193404 295372
rect 191340 295332 191346 295344
rect 193398 295332 193404 295344
rect 193456 295332 193462 295384
rect 86954 294652 86960 294704
rect 87012 294692 87018 294704
rect 152642 294692 152648 294704
rect 87012 294664 152648 294692
rect 87012 294652 87018 294664
rect 152642 294652 152648 294664
rect 152700 294652 152706 294704
rect 19242 294584 19248 294636
rect 19300 294624 19306 294636
rect 149698 294624 149704 294636
rect 19300 294596 149704 294624
rect 19300 294584 19306 294596
rect 149698 294584 149704 294596
rect 149756 294584 149762 294636
rect 152734 294584 152740 294636
rect 152792 294624 152798 294636
rect 189902 294624 189908 294636
rect 152792 294596 189908 294624
rect 152792 294584 152798 294596
rect 189902 294584 189908 294596
rect 189960 294584 189966 294636
rect 255406 294584 255412 294636
rect 255464 294624 255470 294636
rect 258258 294624 258264 294636
rect 255464 294596 258264 294624
rect 255464 294584 255470 294596
rect 258258 294584 258264 294596
rect 258316 294624 258322 294636
rect 280338 294624 280344 294636
rect 258316 294596 280344 294624
rect 258316 294584 258322 294596
rect 280338 294584 280344 294596
rect 280396 294584 280402 294636
rect 255406 293972 255412 294024
rect 255464 294012 255470 294024
rect 277578 294012 277584 294024
rect 255464 293984 277584 294012
rect 255464 293972 255470 293984
rect 277578 293972 277584 293984
rect 277636 293972 277642 294024
rect 93762 293904 93768 293956
rect 93820 293944 93826 293956
rect 117222 293944 117228 293956
rect 93820 293916 117228 293944
rect 93820 293904 93826 293916
rect 117222 293904 117228 293916
rect 117280 293904 117286 293956
rect 138014 293904 138020 293956
rect 138072 293944 138078 293956
rect 143626 293944 143632 293956
rect 138072 293916 143632 293944
rect 138072 293904 138078 293916
rect 143626 293904 143632 293916
rect 143684 293944 143690 293956
rect 155770 293944 155776 293956
rect 143684 293916 155776 293944
rect 143684 293904 143690 293916
rect 155770 293904 155776 293916
rect 155828 293944 155834 293956
rect 191190 293944 191196 293956
rect 155828 293916 191196 293944
rect 155828 293904 155834 293916
rect 191190 293904 191196 293916
rect 191248 293904 191254 293956
rect 253842 293904 253848 293956
rect 253900 293944 253906 293956
rect 269114 293944 269120 293956
rect 253900 293916 269120 293944
rect 253900 293904 253906 293916
rect 269114 293904 269120 293916
rect 269172 293904 269178 293956
rect 58986 293224 58992 293276
rect 59044 293264 59050 293276
rect 78674 293264 78680 293276
rect 59044 293236 78680 293264
rect 59044 293224 59050 293236
rect 78674 293224 78680 293236
rect 78732 293224 78738 293276
rect 96706 293224 96712 293276
rect 96764 293264 96770 293276
rect 141694 293264 141700 293276
rect 96764 293236 141700 293264
rect 96764 293224 96770 293236
rect 141694 293224 141700 293236
rect 141752 293224 141758 293276
rect 166902 293224 166908 293276
rect 166960 293264 166966 293276
rect 187694 293264 187700 293276
rect 166960 293236 187700 293264
rect 166960 293224 166966 293236
rect 187694 293224 187700 293236
rect 187752 293224 187758 293276
rect 255498 293224 255504 293276
rect 255556 293264 255562 293276
rect 258442 293264 258448 293276
rect 255556 293236 258448 293264
rect 255556 293224 255562 293236
rect 258442 293224 258448 293236
rect 258500 293264 258506 293276
rect 289998 293264 290004 293276
rect 258500 293236 290004 293264
rect 258500 293224 258506 293236
rect 289998 293224 290004 293236
rect 290056 293224 290062 293276
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 14458 292584 14464 292596
rect 3568 292556 14464 292584
rect 3568 292544 3574 292556
rect 14458 292544 14464 292556
rect 14516 292544 14522 292596
rect 65794 291796 65800 291848
rect 65852 291836 65858 291848
rect 86218 291836 86224 291848
rect 65852 291808 86224 291836
rect 65852 291796 65858 291808
rect 86218 291796 86224 291808
rect 86276 291796 86282 291848
rect 163682 291796 163688 291848
rect 163740 291836 163746 291848
rect 178954 291836 178960 291848
rect 163740 291808 178960 291836
rect 163740 291796 163746 291808
rect 178954 291796 178960 291808
rect 179012 291796 179018 291848
rect 256418 291796 256424 291848
rect 256476 291836 256482 291848
rect 264974 291836 264980 291848
rect 256476 291808 264980 291836
rect 256476 291796 256482 291808
rect 264974 291796 264980 291808
rect 265032 291796 265038 291848
rect 253842 291728 253848 291780
rect 253900 291768 253906 291780
rect 256602 291768 256608 291780
rect 253900 291740 256608 291768
rect 253900 291728 253906 291740
rect 256602 291728 256608 291740
rect 256660 291728 256666 291780
rect 104894 291292 104900 291304
rect 89686 291264 104900 291292
rect 85850 291184 85856 291236
rect 85908 291224 85914 291236
rect 86770 291224 86776 291236
rect 85908 291196 86776 291224
rect 85908 291184 85914 291196
rect 86770 291184 86776 291196
rect 86828 291224 86834 291236
rect 89686 291224 89714 291264
rect 104894 291252 104900 291264
rect 104952 291252 104958 291304
rect 86828 291196 89714 291224
rect 86828 291184 86834 291196
rect 95142 291184 95148 291236
rect 95200 291224 95206 291236
rect 127710 291224 127716 291236
rect 95200 291196 127716 291224
rect 95200 291184 95206 291196
rect 127710 291184 127716 291196
rect 127768 291184 127774 291236
rect 256510 291048 256516 291100
rect 256568 291088 256574 291100
rect 263870 291088 263876 291100
rect 256568 291060 263876 291088
rect 256568 291048 256574 291060
rect 263870 291048 263876 291060
rect 263928 291048 263934 291100
rect 98454 290504 98460 290556
rect 98512 290544 98518 290556
rect 138014 290544 138020 290556
rect 98512 290516 138020 290544
rect 98512 290504 98518 290516
rect 138014 290504 138020 290516
rect 138072 290504 138078 290556
rect 173158 290504 173164 290556
rect 173216 290544 173222 290556
rect 184198 290544 184204 290556
rect 173216 290516 184204 290544
rect 173216 290504 173222 290516
rect 184198 290504 184204 290516
rect 184256 290504 184262 290556
rect 33778 290436 33784 290488
rect 33836 290476 33842 290488
rect 87598 290476 87604 290488
rect 33836 290448 87604 290476
rect 33836 290436 33842 290448
rect 87598 290436 87604 290448
rect 87656 290436 87662 290488
rect 106182 290436 106188 290488
rect 106240 290476 106246 290488
rect 177482 290476 177488 290488
rect 106240 290448 177488 290476
rect 106240 290436 106246 290448
rect 177482 290436 177488 290448
rect 177540 290436 177546 290488
rect 71866 289824 71872 289876
rect 71924 289864 71930 289876
rect 104986 289864 104992 289876
rect 71924 289836 104992 289864
rect 71924 289824 71930 289836
rect 104986 289824 104992 289836
rect 105044 289864 105050 289876
rect 106182 289864 106188 289876
rect 105044 289836 106188 289864
rect 105044 289824 105050 289836
rect 106182 289824 106188 289836
rect 106240 289824 106246 289876
rect 177574 289824 177580 289876
rect 177632 289864 177638 289876
rect 191742 289864 191748 289876
rect 177632 289836 191748 289864
rect 177632 289824 177638 289836
rect 191742 289824 191748 289836
rect 191800 289824 191806 289876
rect 79962 289756 79968 289808
rect 80020 289796 80026 289808
rect 173802 289796 173808 289808
rect 80020 289768 173808 289796
rect 80020 289756 80026 289768
rect 173802 289756 173808 289768
rect 173860 289796 173866 289808
rect 191650 289796 191656 289808
rect 173860 289768 191656 289796
rect 173860 289756 173866 289768
rect 191650 289756 191656 289768
rect 191708 289756 191714 289808
rect 61838 289076 61844 289128
rect 61896 289116 61902 289128
rect 77478 289116 77484 289128
rect 61896 289088 77484 289116
rect 61896 289076 61902 289088
rect 77478 289076 77484 289088
rect 77536 289116 77542 289128
rect 80146 289116 80152 289128
rect 77536 289088 80152 289116
rect 77536 289076 77542 289088
rect 80146 289076 80152 289088
rect 80204 289076 80210 289128
rect 180702 289076 180708 289128
rect 180760 289116 180766 289128
rect 184198 289116 184204 289128
rect 180760 289088 184204 289116
rect 180760 289076 180766 289088
rect 184198 289076 184204 289088
rect 184256 289076 184262 289128
rect 255958 288872 255964 288924
rect 256016 288912 256022 288924
rect 259730 288912 259736 288924
rect 256016 288884 259736 288912
rect 256016 288872 256022 288884
rect 259730 288872 259736 288884
rect 259788 288872 259794 288924
rect 97534 288396 97540 288448
rect 97592 288436 97598 288448
rect 97902 288436 97908 288448
rect 97592 288408 97908 288436
rect 97592 288396 97598 288408
rect 97902 288396 97908 288408
rect 97960 288436 97966 288448
rect 109034 288436 109040 288448
rect 97960 288408 109040 288436
rect 97960 288396 97966 288408
rect 109034 288396 109040 288408
rect 109092 288396 109098 288448
rect 259362 288396 259368 288448
rect 259420 288436 259426 288448
rect 261110 288436 261116 288448
rect 259420 288408 261116 288436
rect 259420 288396 259426 288408
rect 261110 288396 261116 288408
rect 261168 288396 261174 288448
rect 255866 288328 255872 288380
rect 255924 288368 255930 288380
rect 276106 288368 276112 288380
rect 255924 288340 276112 288368
rect 255924 288328 255930 288340
rect 276106 288328 276112 288340
rect 276164 288328 276170 288380
rect 255774 288260 255780 288312
rect 255832 288300 255838 288312
rect 258074 288300 258080 288312
rect 255832 288272 258080 288300
rect 255832 288260 255838 288272
rect 258074 288260 258080 288272
rect 258132 288260 258138 288312
rect 116486 287716 116492 287768
rect 116544 287756 116550 287768
rect 184842 287756 184848 287768
rect 116544 287728 184848 287756
rect 116544 287716 116550 287728
rect 184842 287716 184848 287728
rect 184900 287756 184906 287768
rect 191742 287756 191748 287768
rect 184900 287728 191748 287756
rect 184900 287716 184906 287728
rect 191742 287716 191748 287728
rect 191800 287716 191806 287768
rect 78582 287648 78588 287700
rect 78640 287688 78646 287700
rect 186958 287688 186964 287700
rect 78640 287660 186964 287688
rect 78640 287648 78646 287660
rect 186958 287648 186964 287660
rect 187016 287648 187022 287700
rect 87874 287036 87880 287088
rect 87932 287076 87938 287088
rect 88150 287076 88156 287088
rect 87932 287048 88156 287076
rect 87932 287036 87938 287048
rect 88150 287036 88156 287048
rect 88208 287076 88214 287088
rect 104342 287076 104348 287088
rect 88208 287048 104348 287076
rect 88208 287036 88214 287048
rect 104342 287036 104348 287048
rect 104400 287036 104406 287088
rect 276750 287036 276756 287088
rect 276808 287076 276814 287088
rect 279050 287076 279056 287088
rect 276808 287048 279056 287076
rect 276808 287036 276814 287048
rect 279050 287036 279056 287048
rect 279108 287036 279114 287088
rect 61930 286968 61936 287020
rect 61988 287008 61994 287020
rect 65978 287008 65984 287020
rect 61988 286980 65984 287008
rect 61988 286968 61994 286980
rect 65978 286968 65984 286980
rect 66036 286968 66042 287020
rect 95786 286968 95792 287020
rect 95844 287008 95850 287020
rect 97534 287008 97540 287020
rect 95844 286980 97540 287008
rect 95844 286968 95850 286980
rect 97534 286968 97540 286980
rect 97592 286968 97598 287020
rect 127710 286968 127716 287020
rect 127768 287008 127774 287020
rect 142890 287008 142896 287020
rect 127768 286980 142896 287008
rect 127768 286968 127774 286980
rect 142890 286968 142896 286980
rect 142948 286968 142954 287020
rect 256602 286628 256608 286680
rect 256660 286668 256666 286680
rect 261018 286668 261024 286680
rect 256660 286640 261024 286668
rect 256660 286628 256666 286640
rect 261018 286628 261024 286640
rect 261076 286628 261082 286680
rect 75730 286288 75736 286340
rect 75788 286328 75794 286340
rect 185578 286328 185584 286340
rect 75788 286300 185584 286328
rect 75788 286288 75794 286300
rect 185578 286288 185584 286300
rect 185636 286288 185642 286340
rect 90910 286220 90916 286272
rect 90968 286260 90974 286272
rect 94498 286260 94504 286272
rect 90968 286232 94504 286260
rect 90968 286220 90974 286232
rect 94498 286220 94504 286232
rect 94556 286220 94562 286272
rect 85298 285880 85304 285932
rect 85356 285920 85362 285932
rect 87690 285920 87696 285932
rect 85356 285892 87696 285920
rect 85356 285880 85362 285892
rect 87690 285880 87696 285892
rect 87748 285880 87754 285932
rect 81250 285852 81256 285864
rect 80026 285824 81256 285852
rect 68646 285744 68652 285796
rect 68704 285784 68710 285796
rect 80026 285784 80054 285824
rect 81250 285812 81256 285824
rect 81308 285852 81314 285864
rect 83458 285852 83464 285864
rect 81308 285824 83464 285852
rect 81308 285812 81314 285824
rect 83458 285812 83464 285824
rect 83516 285812 83522 285864
rect 68704 285756 80054 285784
rect 68704 285744 68710 285756
rect 71314 285676 71320 285728
rect 71372 285716 71378 285728
rect 72418 285716 72424 285728
rect 71372 285688 72424 285716
rect 71372 285676 71378 285688
rect 72418 285676 72424 285688
rect 72476 285676 72482 285728
rect 74810 285676 74816 285728
rect 74868 285716 74874 285728
rect 75822 285716 75828 285728
rect 74868 285688 75828 285716
rect 74868 285676 74874 285688
rect 75822 285676 75828 285688
rect 75880 285676 75886 285728
rect 79226 285676 79232 285728
rect 79284 285716 79290 285728
rect 79962 285716 79968 285728
rect 79284 285688 79968 285716
rect 79284 285676 79290 285688
rect 79962 285676 79968 285688
rect 80020 285676 80026 285728
rect 256418 285676 256424 285728
rect 256476 285716 256482 285728
rect 262490 285716 262496 285728
rect 256476 285688 262496 285716
rect 256476 285676 256482 285688
rect 262490 285676 262496 285688
rect 262548 285716 262554 285728
rect 263962 285716 263968 285728
rect 262548 285688 263968 285716
rect 262548 285676 262554 285688
rect 263962 285676 263968 285688
rect 264020 285676 264026 285728
rect 256602 285608 256608 285660
rect 256660 285648 256666 285660
rect 263594 285648 263600 285660
rect 256660 285620 263600 285648
rect 256660 285608 256666 285620
rect 263594 285608 263600 285620
rect 263652 285608 263658 285660
rect 140038 284996 140044 285048
rect 140096 285036 140102 285048
rect 149790 285036 149796 285048
rect 140096 285008 149796 285036
rect 140096 284996 140102 285008
rect 149790 284996 149796 285008
rect 149848 284996 149854 285048
rect 75914 284928 75920 284980
rect 75972 284968 75978 284980
rect 76374 284968 76380 284980
rect 75972 284940 76380 284968
rect 75972 284928 75978 284940
rect 76374 284928 76380 284940
rect 76432 284928 76438 284980
rect 149698 284928 149704 284980
rect 149756 284968 149762 284980
rect 180150 284968 180156 284980
rect 149756 284940 180156 284968
rect 149756 284928 149762 284940
rect 180150 284928 180156 284940
rect 180208 284928 180214 284980
rect 266630 284792 266636 284844
rect 266688 284832 266694 284844
rect 267826 284832 267832 284844
rect 266688 284804 267832 284832
rect 266688 284792 266694 284804
rect 267826 284792 267832 284804
rect 267884 284792 267890 284844
rect 53558 284452 53564 284504
rect 53616 284492 53622 284504
rect 71314 284492 71320 284504
rect 53616 284464 71320 284492
rect 53616 284452 53622 284464
rect 71314 284452 71320 284464
rect 71372 284452 71378 284504
rect 70854 284384 70860 284436
rect 70912 284424 70918 284436
rect 99374 284424 99380 284436
rect 70912 284396 99380 284424
rect 70912 284384 70918 284396
rect 99374 284384 99380 284396
rect 99432 284384 99438 284436
rect 67358 284316 67364 284368
rect 67416 284356 67422 284368
rect 160094 284356 160100 284368
rect 67416 284328 160100 284356
rect 67416 284316 67422 284328
rect 160094 284316 160100 284328
rect 160152 284316 160158 284368
rect 167822 284316 167828 284368
rect 167880 284356 167886 284368
rect 191742 284356 191748 284368
rect 167880 284328 191748 284356
rect 167880 284316 167886 284328
rect 191742 284316 191748 284328
rect 191800 284316 191806 284368
rect 149054 284248 149060 284300
rect 149112 284288 149118 284300
rect 149112 284260 180794 284288
rect 149112 284248 149118 284260
rect 180766 284220 180794 284260
rect 256602 284248 256608 284300
rect 256660 284288 256666 284300
rect 294046 284288 294052 284300
rect 256660 284260 294052 284288
rect 256660 284248 256666 284260
rect 294046 284248 294052 284260
rect 294104 284248 294110 284300
rect 191742 284220 191748 284232
rect 180766 284192 191748 284220
rect 191742 284180 191748 284192
rect 191800 284180 191806 284232
rect 256326 284180 256332 284232
rect 256384 284220 256390 284232
rect 273254 284220 273260 284232
rect 256384 284192 273260 284220
rect 256384 284180 256390 284192
rect 273254 284180 273260 284192
rect 273312 284180 273318 284232
rect 88288 283704 88294 283756
rect 88346 283744 88352 283756
rect 89530 283744 89536 283756
rect 88346 283716 89536 283744
rect 88346 283704 88352 283716
rect 89530 283704 89536 283716
rect 89588 283704 89594 283756
rect 92704 283704 92710 283756
rect 92762 283744 92768 283756
rect 93762 283744 93768 283756
rect 92762 283716 93768 283744
rect 92762 283704 92768 283716
rect 93762 283704 93768 283716
rect 93820 283704 93826 283756
rect 96890 283364 96896 283416
rect 96948 283404 96954 283416
rect 97258 283404 97264 283416
rect 96948 283376 97264 283404
rect 96948 283364 96954 283376
rect 97258 283364 97264 283376
rect 97316 283364 97322 283416
rect 184658 283228 184664 283280
rect 184716 283268 184722 283280
rect 187694 283268 187700 283280
rect 184716 283240 187700 283268
rect 184716 283228 184722 283240
rect 187694 283228 187700 283240
rect 187752 283228 187758 283280
rect 86862 283024 86868 283076
rect 86920 283064 86926 283076
rect 98914 283064 98920 283076
rect 86920 283036 98920 283064
rect 86920 283024 86926 283036
rect 98914 283024 98920 283036
rect 98972 283024 98978 283076
rect 63218 282956 63224 283008
rect 63276 282996 63282 283008
rect 76006 282996 76012 283008
rect 63276 282968 76012 282996
rect 63276 282956 63282 282968
rect 76006 282956 76012 282968
rect 76064 282956 76070 283008
rect 94130 282956 94136 283008
rect 94188 282996 94194 283008
rect 98822 282996 98828 283008
rect 94188 282968 98828 282996
rect 94188 282956 94194 282968
rect 98822 282956 98828 282968
rect 98880 282956 98886 283008
rect 56410 282888 56416 282940
rect 56468 282928 56474 282940
rect 66254 282928 66260 282940
rect 56468 282900 66260 282928
rect 56468 282888 56474 282900
rect 66254 282888 66260 282900
rect 66312 282888 66318 282940
rect 68830 282888 68836 282940
rect 68888 282928 68894 282940
rect 173802 282928 173808 282940
rect 68888 282900 173808 282928
rect 68888 282888 68894 282900
rect 173802 282888 173808 282900
rect 173860 282928 173866 282940
rect 175918 282928 175924 282940
rect 173860 282900 175924 282928
rect 173860 282888 173866 282900
rect 175918 282888 175924 282900
rect 175976 282888 175982 282940
rect 119338 282820 119344 282872
rect 119396 282860 119402 282872
rect 124950 282860 124956 282872
rect 119396 282832 124956 282860
rect 119396 282820 119402 282832
rect 124950 282820 124956 282832
rect 125008 282820 125014 282872
rect 44082 282140 44088 282192
rect 44140 282180 44146 282192
rect 63494 282180 63500 282192
rect 44140 282152 63500 282180
rect 44140 282140 44146 282152
rect 63494 282140 63500 282152
rect 63552 282140 63558 282192
rect 135898 282140 135904 282192
rect 135956 282180 135962 282192
rect 191834 282180 191840 282192
rect 135956 282152 191840 282180
rect 135956 282140 135962 282152
rect 191834 282140 191840 282152
rect 191892 282140 191898 282192
rect 255498 282140 255504 282192
rect 255556 282180 255562 282192
rect 259822 282180 259828 282192
rect 255556 282152 259828 282180
rect 255556 282140 255562 282152
rect 259822 282140 259828 282152
rect 259880 282180 259886 282192
rect 263686 282180 263692 282192
rect 259880 282152 263692 282180
rect 259880 282140 259886 282152
rect 263686 282140 263692 282152
rect 263744 282140 263750 282192
rect 63494 281596 63500 281648
rect 63552 281636 63558 281648
rect 64598 281636 64604 281648
rect 63552 281608 64604 281636
rect 63552 281596 63558 281608
rect 64598 281596 64604 281608
rect 64656 281636 64662 281648
rect 102778 281636 102784 281648
rect 64656 281608 102784 281636
rect 64656 281596 64662 281608
rect 102778 281596 102784 281608
rect 102836 281596 102842 281648
rect 100754 281528 100760 281580
rect 100812 281568 100818 281580
rect 180334 281568 180340 281580
rect 100812 281540 180340 281568
rect 100812 281528 100818 281540
rect 180334 281528 180340 281540
rect 180392 281528 180398 281580
rect 181530 281528 181536 281580
rect 181588 281568 181594 281580
rect 190454 281568 190460 281580
rect 181588 281540 190460 281568
rect 181588 281528 181594 281540
rect 190454 281528 190460 281540
rect 190512 281528 190518 281580
rect 255314 281460 255320 281512
rect 255372 281500 255378 281512
rect 281810 281500 281816 281512
rect 255372 281472 281816 281500
rect 255372 281460 255378 281472
rect 281810 281460 281816 281472
rect 281868 281460 281874 281512
rect 255498 281392 255504 281444
rect 255556 281432 255562 281444
rect 262306 281432 262312 281444
rect 255556 281404 262312 281432
rect 255556 281392 255562 281404
rect 262306 281392 262312 281404
rect 262364 281392 262370 281444
rect 119338 280848 119344 280900
rect 119396 280888 119402 280900
rect 155310 280888 155316 280900
rect 119396 280860 155316 280888
rect 119396 280848 119402 280860
rect 155310 280848 155316 280860
rect 155368 280848 155374 280900
rect 176470 280848 176476 280900
rect 176528 280888 176534 280900
rect 190546 280888 190552 280900
rect 176528 280860 190552 280888
rect 176528 280848 176534 280860
rect 190546 280848 190552 280860
rect 190604 280848 190610 280900
rect 99374 280780 99380 280832
rect 99432 280820 99438 280832
rect 162670 280820 162676 280832
rect 99432 280792 162676 280820
rect 99432 280780 99438 280792
rect 162670 280780 162676 280792
rect 162728 280820 162734 280832
rect 178678 280820 178684 280832
rect 162728 280792 178684 280820
rect 162728 280780 162734 280792
rect 178678 280780 178684 280792
rect 178736 280780 178742 280832
rect 4798 280168 4804 280220
rect 4856 280208 4862 280220
rect 67542 280208 67548 280220
rect 4856 280180 67548 280208
rect 4856 280168 4862 280180
rect 67542 280168 67548 280180
rect 67600 280208 67606 280220
rect 68830 280208 68836 280220
rect 67600 280180 68836 280208
rect 67600 280168 67606 280180
rect 68830 280168 68836 280180
rect 68888 280168 68894 280220
rect 100846 280100 100852 280152
rect 100904 280140 100910 280152
rect 162118 280140 162124 280152
rect 100904 280112 162124 280140
rect 100904 280100 100910 280112
rect 162118 280100 162124 280112
rect 162176 280100 162182 280152
rect 165522 280100 165528 280152
rect 165580 280140 165586 280152
rect 175274 280140 175280 280152
rect 165580 280112 175280 280140
rect 165580 280100 165586 280112
rect 175274 280100 175280 280112
rect 175332 280100 175338 280152
rect 255498 280100 255504 280152
rect 255556 280140 255562 280152
rect 291378 280140 291384 280152
rect 255556 280112 291384 280140
rect 255556 280100 255562 280112
rect 291378 280100 291384 280112
rect 291436 280100 291442 280152
rect 159450 280032 159456 280084
rect 159508 280072 159514 280084
rect 160094 280072 160100 280084
rect 159508 280044 160100 280072
rect 159508 280032 159514 280044
rect 160094 280032 160100 280044
rect 160152 280072 160158 280084
rect 190454 280072 190460 280084
rect 160152 280044 190460 280072
rect 160152 280032 160158 280044
rect 190454 280032 190460 280044
rect 190512 280032 190518 280084
rect 3418 279624 3424 279676
rect 3476 279664 3482 279676
rect 7650 279664 7656 279676
rect 3476 279636 7656 279664
rect 3476 279624 3482 279636
rect 7650 279624 7656 279636
rect 7708 279624 7714 279676
rect 7558 279420 7564 279472
rect 7616 279460 7622 279472
rect 37090 279460 37096 279472
rect 7616 279432 37096 279460
rect 7616 279420 7622 279432
rect 37090 279420 37096 279432
rect 37148 279460 37154 279472
rect 60458 279460 60464 279472
rect 37148 279432 60464 279460
rect 37148 279420 37154 279432
rect 60458 279420 60464 279432
rect 60516 279460 60522 279472
rect 66806 279460 66812 279472
rect 60516 279432 66812 279460
rect 60516 279420 60522 279432
rect 66806 279420 66812 279432
rect 66864 279420 66870 279472
rect 179322 279420 179328 279472
rect 179380 279460 179386 279472
rect 191282 279460 191288 279472
rect 179380 279432 191288 279460
rect 179380 279420 179386 279432
rect 191282 279420 191288 279432
rect 191340 279420 191346 279472
rect 262306 279420 262312 279472
rect 262364 279460 262370 279472
rect 270586 279460 270592 279472
rect 262364 279432 270592 279460
rect 262364 279420 262370 279432
rect 270586 279420 270592 279432
rect 270644 279420 270650 279472
rect 255314 278740 255320 278792
rect 255372 278780 255378 278792
rect 262306 278780 262312 278792
rect 255372 278752 262312 278780
rect 255372 278740 255378 278752
rect 262306 278740 262312 278752
rect 262364 278740 262370 278792
rect 64598 278672 64604 278724
rect 64656 278712 64662 278724
rect 66806 278712 66812 278724
rect 64656 278684 66812 278712
rect 64656 278672 64662 278684
rect 66806 278672 66812 278684
rect 66864 278672 66870 278724
rect 100754 278604 100760 278656
rect 100812 278644 100818 278656
rect 104434 278644 104440 278656
rect 100812 278616 104440 278644
rect 100812 278604 100818 278616
rect 104434 278604 104440 278616
rect 104492 278604 104498 278656
rect 112806 278060 112812 278112
rect 112864 278100 112870 278112
rect 116578 278100 116584 278112
rect 112864 278072 116584 278100
rect 112864 278060 112870 278072
rect 116578 278060 116584 278072
rect 116636 278060 116642 278112
rect 144178 278060 144184 278112
rect 144236 278100 144242 278112
rect 167638 278100 167644 278112
rect 144236 278072 167644 278100
rect 144236 278060 144242 278072
rect 167638 278060 167644 278072
rect 167696 278060 167702 278112
rect 255498 278060 255504 278112
rect 255556 278100 255562 278112
rect 266538 278100 266544 278112
rect 255556 278072 266544 278100
rect 255556 278060 255562 278072
rect 266538 278060 266544 278072
rect 266596 278060 266602 278112
rect 112622 277992 112628 278044
rect 112680 278032 112686 278044
rect 152550 278032 152556 278044
rect 112680 278004 152556 278032
rect 112680 277992 112686 278004
rect 152550 277992 152556 278004
rect 152608 278032 152614 278044
rect 190270 278032 190276 278044
rect 152608 278004 190276 278032
rect 152608 277992 152614 278004
rect 190270 277992 190276 278004
rect 190328 278032 190334 278044
rect 190454 278032 190460 278044
rect 190328 278004 190460 278032
rect 190328 277992 190334 278004
rect 190454 277992 190460 278004
rect 190512 277992 190518 278044
rect 258074 277992 258080 278044
rect 258132 278032 258138 278044
rect 295518 278032 295524 278044
rect 258132 278004 295524 278032
rect 258132 277992 258138 278004
rect 295518 277992 295524 278004
rect 295576 277992 295582 278044
rect 52362 277312 52368 277364
rect 52420 277352 52426 277364
rect 66806 277352 66812 277364
rect 52420 277324 66812 277352
rect 52420 277312 52426 277324
rect 66806 277312 66812 277324
rect 66864 277312 66870 277364
rect 100754 277312 100760 277364
rect 100812 277352 100818 277364
rect 123478 277352 123484 277364
rect 100812 277324 123484 277352
rect 100812 277312 100818 277324
rect 123478 277312 123484 277324
rect 123536 277312 123542 277364
rect 255314 277312 255320 277364
rect 255372 277352 255378 277364
rect 271966 277352 271972 277364
rect 255372 277324 271972 277352
rect 255372 277312 255378 277324
rect 271966 277312 271972 277324
rect 272024 277312 272030 277364
rect 255498 277244 255504 277296
rect 255556 277284 255562 277296
rect 267734 277284 267740 277296
rect 255556 277256 267740 277284
rect 255556 277244 255562 277256
rect 267734 277244 267740 277256
rect 267792 277244 267798 277296
rect 98914 276632 98920 276684
rect 98972 276672 98978 276684
rect 176654 276672 176660 276684
rect 98972 276644 176660 276672
rect 98972 276632 98978 276644
rect 176654 276632 176660 276644
rect 176712 276632 176718 276684
rect 63310 276020 63316 276072
rect 63368 276060 63374 276072
rect 67634 276060 67640 276072
rect 63368 276032 67640 276060
rect 63368 276020 63374 276032
rect 67634 276020 67640 276032
rect 67692 276020 67698 276072
rect 148502 276020 148508 276072
rect 148560 276060 148566 276072
rect 190454 276060 190460 276072
rect 148560 276032 190460 276060
rect 148560 276020 148566 276032
rect 190454 276020 190460 276032
rect 190512 276020 190518 276072
rect 57882 275952 57888 276004
rect 57940 275992 57946 276004
rect 66806 275992 66812 276004
rect 57940 275964 66812 275992
rect 57940 275952 57946 275964
rect 66806 275952 66812 275964
rect 66864 275952 66870 276004
rect 176654 275952 176660 276004
rect 176712 275992 176718 276004
rect 177850 275992 177856 276004
rect 176712 275964 177856 275992
rect 176712 275952 176718 275964
rect 177850 275952 177856 275964
rect 177908 275992 177914 276004
rect 181438 275992 181444 276004
rect 177908 275964 181444 275992
rect 177908 275952 177914 275964
rect 181438 275952 181444 275964
rect 181496 275952 181502 276004
rect 255314 275952 255320 276004
rect 255372 275992 255378 276004
rect 270494 275992 270500 276004
rect 255372 275964 270500 275992
rect 255372 275952 255378 275964
rect 270494 275952 270500 275964
rect 270552 275952 270558 276004
rect 255498 275476 255504 275528
rect 255556 275516 255562 275528
rect 258074 275516 258080 275528
rect 255556 275488 258080 275516
rect 255556 275476 255562 275488
rect 258074 275476 258080 275488
rect 258132 275476 258138 275528
rect 101674 275340 101680 275392
rect 101732 275380 101738 275392
rect 136082 275380 136088 275392
rect 101732 275352 136088 275380
rect 101732 275340 101738 275352
rect 136082 275340 136088 275352
rect 136140 275340 136146 275392
rect 57698 275272 57704 275324
rect 57756 275312 57762 275324
rect 66438 275312 66444 275324
rect 57756 275284 66444 275312
rect 57756 275272 57762 275284
rect 66438 275272 66444 275284
rect 66496 275312 66502 275324
rect 66714 275312 66720 275324
rect 66496 275284 66720 275312
rect 66496 275272 66502 275284
rect 66714 275272 66720 275284
rect 66772 275272 66778 275324
rect 100938 275272 100944 275324
rect 100996 275312 101002 275324
rect 169202 275312 169208 275324
rect 100996 275284 169208 275312
rect 100996 275272 101002 275284
rect 169202 275272 169208 275284
rect 169260 275272 169266 275324
rect 259362 275272 259368 275324
rect 259420 275312 259426 275324
rect 292574 275312 292580 275324
rect 259420 275284 292580 275312
rect 259420 275272 259426 275284
rect 292574 275272 292580 275284
rect 292632 275272 292638 275324
rect 184842 274728 184848 274780
rect 184900 274768 184906 274780
rect 186406 274768 186412 274780
rect 184900 274740 186412 274768
rect 184900 274728 184906 274740
rect 186406 274728 186412 274740
rect 186464 274728 186470 274780
rect 187050 274728 187056 274780
rect 187108 274768 187114 274780
rect 190546 274768 190552 274780
rect 187108 274740 190552 274768
rect 187108 274728 187114 274740
rect 190546 274728 190552 274740
rect 190604 274728 190610 274780
rect 171962 274660 171968 274712
rect 172020 274700 172026 274712
rect 190454 274700 190460 274712
rect 172020 274672 190460 274700
rect 172020 274660 172026 274672
rect 190454 274660 190460 274672
rect 190512 274660 190518 274712
rect 100754 274592 100760 274644
rect 100812 274632 100818 274644
rect 170398 274632 170404 274644
rect 100812 274604 170404 274632
rect 100812 274592 100818 274604
rect 170398 274592 170404 274604
rect 170456 274592 170462 274644
rect 255314 274592 255320 274644
rect 255372 274632 255378 274644
rect 281718 274632 281724 274644
rect 255372 274604 281724 274632
rect 255372 274592 255378 274604
rect 281718 274592 281724 274604
rect 281776 274592 281782 274644
rect 100846 274524 100852 274576
rect 100904 274564 100910 274576
rect 135990 274564 135996 274576
rect 100904 274536 135996 274564
rect 100904 274524 100910 274536
rect 135990 274524 135996 274536
rect 136048 274524 136054 274576
rect 255498 274252 255504 274304
rect 255556 274292 255562 274304
rect 259270 274292 259276 274304
rect 255556 274264 259276 274292
rect 255556 274252 255562 274264
rect 259270 274252 259276 274264
rect 259328 274292 259334 274304
rect 259546 274292 259552 274304
rect 259328 274264 259552 274292
rect 259328 274252 259334 274264
rect 259546 274252 259552 274264
rect 259604 274252 259610 274304
rect 145742 273912 145748 273964
rect 145800 273952 145806 273964
rect 159542 273952 159548 273964
rect 145800 273924 159548 273952
rect 145800 273912 145806 273924
rect 159542 273912 159548 273924
rect 159600 273912 159606 273964
rect 58894 273300 58900 273352
rect 58952 273340 58958 273352
rect 60642 273340 60648 273352
rect 58952 273312 60648 273340
rect 58952 273300 58958 273312
rect 60642 273300 60648 273312
rect 60700 273340 60706 273352
rect 66806 273340 66812 273352
rect 60700 273312 66812 273340
rect 60700 273300 60706 273312
rect 66806 273300 66812 273312
rect 66864 273300 66870 273352
rect 182910 273232 182916 273284
rect 182968 273272 182974 273284
rect 190454 273272 190460 273284
rect 182968 273244 190460 273272
rect 182968 273232 182974 273244
rect 190454 273232 190460 273244
rect 190512 273232 190518 273284
rect 100754 273164 100760 273216
rect 100812 273204 100818 273216
rect 129734 273204 129740 273216
rect 100812 273176 129740 273204
rect 100812 273164 100818 273176
rect 129734 273164 129740 273176
rect 129792 273164 129798 273216
rect 278682 272960 278688 273012
rect 278740 273000 278746 273012
rect 281718 273000 281724 273012
rect 278740 272972 281724 273000
rect 278740 272960 278746 272972
rect 281718 272960 281724 272972
rect 281776 272960 281782 273012
rect 255498 272892 255504 272944
rect 255556 272932 255562 272944
rect 259362 272932 259368 272944
rect 255556 272904 259368 272932
rect 255556 272892 255562 272904
rect 259362 272892 259368 272904
rect 259420 272892 259426 272944
rect 146938 272552 146944 272604
rect 146996 272592 147002 272604
rect 173158 272592 173164 272604
rect 146996 272564 173164 272592
rect 146996 272552 147002 272564
rect 173158 272552 173164 272564
rect 173216 272552 173222 272604
rect 100018 272484 100024 272536
rect 100076 272524 100082 272536
rect 115934 272524 115940 272536
rect 100076 272496 115940 272524
rect 100076 272484 100082 272496
rect 115934 272484 115940 272496
rect 115992 272484 115998 272536
rect 129734 272484 129740 272536
rect 129792 272524 129798 272536
rect 159542 272524 159548 272536
rect 129792 272496 159548 272524
rect 129792 272484 129798 272496
rect 159542 272484 159548 272496
rect 159600 272484 159606 272536
rect 61654 271940 61660 271992
rect 61712 271980 61718 271992
rect 61930 271980 61936 271992
rect 61712 271952 61936 271980
rect 61712 271940 61718 271952
rect 61930 271940 61936 271952
rect 61988 271980 61994 271992
rect 66806 271980 66812 271992
rect 61988 271952 66812 271980
rect 61988 271940 61994 271952
rect 66806 271940 66812 271952
rect 66864 271940 66870 271992
rect 181438 271872 181444 271924
rect 181496 271912 181502 271924
rect 190822 271912 190828 271924
rect 181496 271884 190828 271912
rect 181496 271872 181502 271884
rect 190822 271872 190828 271884
rect 190880 271872 190886 271924
rect 101122 271804 101128 271856
rect 101180 271844 101186 271856
rect 101858 271844 101864 271856
rect 101180 271816 101864 271844
rect 101180 271804 101186 271816
rect 101858 271804 101864 271816
rect 101916 271844 101922 271856
rect 128722 271844 128728 271856
rect 101916 271816 128728 271844
rect 101916 271804 101922 271816
rect 128722 271804 128728 271816
rect 128780 271804 128786 271856
rect 271966 271804 271972 271856
rect 272024 271844 272030 271856
rect 276014 271844 276020 271856
rect 272024 271816 276020 271844
rect 272024 271804 272030 271816
rect 276014 271804 276020 271816
rect 276072 271804 276078 271856
rect 128722 271192 128728 271244
rect 128780 271232 128786 271244
rect 129642 271232 129648 271244
rect 128780 271204 129648 271232
rect 128780 271192 128786 271204
rect 129642 271192 129648 271204
rect 129700 271232 129706 271244
rect 135990 271232 135996 271244
rect 129700 271204 135996 271232
rect 129700 271192 129706 271204
rect 135990 271192 135996 271204
rect 136048 271192 136054 271244
rect 137370 271192 137376 271244
rect 137428 271232 137434 271244
rect 188522 271232 188528 271244
rect 137428 271204 188528 271232
rect 137428 271192 137434 271204
rect 188522 271192 188528 271204
rect 188580 271192 188586 271244
rect 98822 271124 98828 271176
rect 98880 271164 98886 271176
rect 155310 271164 155316 271176
rect 98880 271136 155316 271164
rect 98880 271124 98886 271136
rect 155310 271124 155316 271136
rect 155368 271124 155374 271176
rect 255498 270920 255504 270972
rect 255556 270960 255562 270972
rect 258718 270960 258724 270972
rect 255556 270932 258724 270960
rect 255556 270920 255562 270932
rect 258718 270920 258724 270932
rect 258776 270920 258782 270972
rect 63402 270580 63408 270632
rect 63460 270620 63466 270632
rect 64598 270620 64604 270632
rect 63460 270592 64604 270620
rect 63460 270580 63466 270592
rect 64598 270580 64604 270592
rect 64656 270620 64662 270632
rect 66806 270620 66812 270632
rect 64656 270592 66812 270620
rect 64656 270580 64662 270592
rect 66806 270580 66812 270592
rect 66864 270580 66870 270632
rect 188430 270580 188436 270632
rect 188488 270620 188494 270632
rect 191650 270620 191656 270632
rect 188488 270592 191656 270620
rect 188488 270580 188494 270592
rect 191650 270580 191656 270592
rect 191708 270580 191714 270632
rect 255498 270512 255504 270564
rect 255556 270552 255562 270564
rect 271966 270552 271972 270564
rect 255556 270524 271972 270552
rect 255556 270512 255562 270524
rect 271966 270512 271972 270524
rect 272024 270512 272030 270564
rect 57238 270444 57244 270496
rect 57296 270484 57302 270496
rect 57790 270484 57796 270496
rect 57296 270456 57796 270484
rect 57296 270444 57302 270456
rect 57790 270444 57796 270456
rect 57848 270484 57854 270496
rect 66622 270484 66628 270496
rect 57848 270456 66628 270484
rect 57848 270444 57854 270456
rect 66622 270444 66628 270456
rect 66680 270444 66686 270496
rect 100754 270444 100760 270496
rect 100812 270484 100818 270496
rect 112530 270484 112536 270496
rect 100812 270456 112536 270484
rect 100812 270444 100818 270456
rect 112530 270444 112536 270456
rect 112588 270444 112594 270496
rect 255314 270444 255320 270496
rect 255372 270484 255378 270496
rect 277486 270484 277492 270496
rect 255372 270456 277492 270484
rect 255372 270444 255378 270456
rect 277486 270444 277492 270456
rect 277544 270444 277550 270496
rect 255498 270376 255504 270428
rect 255556 270416 255562 270428
rect 262398 270416 262404 270428
rect 255556 270388 262404 270416
rect 255556 270376 255562 270388
rect 262398 270376 262404 270388
rect 262456 270416 262462 270428
rect 262674 270416 262680 270428
rect 262456 270388 262680 270416
rect 262456 270376 262462 270388
rect 262674 270376 262680 270388
rect 262732 270376 262738 270428
rect 152642 269832 152648 269884
rect 152700 269872 152706 269884
rect 171778 269872 171784 269884
rect 152700 269844 171784 269872
rect 152700 269832 152706 269844
rect 171778 269832 171784 269844
rect 171836 269832 171842 269884
rect 98730 269764 98736 269816
rect 98788 269804 98794 269816
rect 160922 269804 160928 269816
rect 98788 269776 160928 269804
rect 98788 269764 98794 269776
rect 160922 269764 160928 269776
rect 160980 269764 160986 269816
rect 187142 269152 187148 269204
rect 187200 269192 187206 269204
rect 191558 269192 191564 269204
rect 187200 269164 191564 269192
rect 187200 269152 187206 269164
rect 191558 269152 191564 269164
rect 191616 269152 191622 269204
rect 53282 269084 53288 269136
rect 53340 269124 53346 269136
rect 57238 269124 57244 269136
rect 53340 269096 57244 269124
rect 53340 269084 53346 269096
rect 57238 269084 57244 269096
rect 57296 269084 57302 269136
rect 170582 269084 170588 269136
rect 170640 269124 170646 269136
rect 190822 269124 190828 269136
rect 170640 269096 190828 269124
rect 170640 269084 170646 269096
rect 190822 269084 190828 269096
rect 190880 269084 190886 269136
rect 262674 269084 262680 269136
rect 262732 269124 262738 269136
rect 269298 269124 269304 269136
rect 262732 269096 269304 269124
rect 262732 269084 262738 269096
rect 269298 269084 269304 269096
rect 269356 269084 269362 269136
rect 267826 269016 267832 269068
rect 267884 269056 267890 269068
rect 270770 269056 270776 269068
rect 267884 269028 270776 269056
rect 267884 269016 267890 269028
rect 270770 269016 270776 269028
rect 270828 269016 270834 269068
rect 166810 268608 166816 268660
rect 166868 268648 166874 268660
rect 168374 268648 168380 268660
rect 166868 268620 168380 268648
rect 166868 268608 166874 268620
rect 168374 268608 168380 268620
rect 168432 268608 168438 268660
rect 100110 268404 100116 268456
rect 100168 268444 100174 268456
rect 134702 268444 134708 268456
rect 100168 268416 134708 268444
rect 100168 268404 100174 268416
rect 134702 268404 134708 268416
rect 134760 268404 134766 268456
rect 145558 268404 145564 268456
rect 145616 268444 145622 268456
rect 173250 268444 173256 268456
rect 145616 268416 173256 268444
rect 145616 268404 145622 268416
rect 173250 268404 173256 268416
rect 173308 268404 173314 268456
rect 113818 268336 113824 268388
rect 113876 268376 113882 268388
rect 166350 268376 166356 268388
rect 113876 268348 166356 268376
rect 113876 268336 113882 268348
rect 166350 268336 166356 268348
rect 166408 268336 166414 268388
rect 100754 267996 100760 268048
rect 100812 268036 100818 268048
rect 104250 268036 104256 268048
rect 100812 268008 104256 268036
rect 100812 267996 100818 268008
rect 104250 267996 104256 268008
rect 104308 267996 104314 268048
rect 255498 267792 255504 267844
rect 255556 267832 255562 267844
rect 267826 267832 267832 267844
rect 255556 267804 267832 267832
rect 255556 267792 255562 267804
rect 267826 267792 267832 267804
rect 267884 267792 267890 267844
rect 54938 267724 54944 267776
rect 54996 267764 55002 267776
rect 57790 267764 57796 267776
rect 54996 267736 57796 267764
rect 54996 267724 55002 267736
rect 57790 267724 57796 267736
rect 57848 267764 57854 267776
rect 66806 267764 66812 267776
rect 57848 267736 66812 267764
rect 57848 267724 57854 267736
rect 66806 267724 66812 267736
rect 66864 267724 66870 267776
rect 173158 267724 173164 267776
rect 173216 267764 173222 267776
rect 191650 267764 191656 267776
rect 173216 267736 191656 267764
rect 173216 267724 173222 267736
rect 191650 267724 191656 267736
rect 191708 267724 191714 267776
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 33778 267696 33784 267708
rect 3568 267668 33784 267696
rect 3568 267656 3574 267668
rect 33778 267656 33784 267668
rect 33836 267656 33842 267708
rect 291286 267656 291292 267708
rect 291344 267696 291350 267708
rect 580258 267696 580264 267708
rect 291344 267668 580264 267696
rect 291344 267656 291350 267668
rect 580258 267656 580264 267668
rect 580316 267656 580322 267708
rect 174538 267112 174544 267164
rect 174596 267152 174602 267164
rect 180794 267152 180800 267164
rect 174596 267124 180800 267152
rect 174596 267112 174602 267124
rect 180794 267112 180800 267124
rect 180852 267112 180858 267164
rect 102226 266976 102232 267028
rect 102284 267016 102290 267028
rect 115198 267016 115204 267028
rect 102284 266988 115204 267016
rect 102284 266976 102290 266988
rect 115198 266976 115204 266988
rect 115256 266976 115262 267028
rect 175182 266976 175188 267028
rect 175240 267016 175246 267028
rect 189074 267016 189080 267028
rect 175240 266988 189080 267016
rect 175240 266976 175246 266988
rect 189074 266976 189080 266988
rect 189132 266976 189138 267028
rect 257338 266976 257344 267028
rect 257396 267016 257402 267028
rect 291286 267016 291292 267028
rect 257396 266988 291292 267016
rect 257396 266976 257402 266988
rect 291286 266976 291292 266988
rect 291344 266976 291350 267028
rect 62022 266364 62028 266416
rect 62080 266404 62086 266416
rect 64782 266404 64788 266416
rect 62080 266376 64788 266404
rect 62080 266364 62086 266376
rect 64782 266364 64788 266376
rect 64840 266404 64846 266416
rect 66806 266404 66812 266416
rect 64840 266376 66812 266404
rect 64840 266364 64846 266376
rect 66806 266364 66812 266376
rect 66864 266364 66870 266416
rect 100754 266364 100760 266416
rect 100812 266404 100818 266416
rect 147122 266404 147128 266416
rect 100812 266376 147128 266404
rect 100812 266364 100818 266376
rect 147122 266364 147128 266376
rect 147180 266364 147186 266416
rect 255314 266364 255320 266416
rect 255372 266404 255378 266416
rect 262398 266404 262404 266416
rect 255372 266376 262404 266404
rect 255372 266364 255378 266376
rect 262398 266364 262404 266376
rect 262456 266364 262462 266416
rect 255498 266296 255504 266348
rect 255556 266336 255562 266348
rect 265066 266336 265072 266348
rect 255556 266308 265072 266336
rect 255556 266296 255562 266308
rect 265066 266296 265072 266308
rect 265124 266296 265130 266348
rect 117314 266024 117320 266076
rect 117372 266064 117378 266076
rect 123478 266064 123484 266076
rect 117372 266036 123484 266064
rect 117372 266024 117378 266036
rect 123478 266024 123484 266036
rect 123536 266024 123542 266076
rect 130470 265616 130476 265668
rect 130528 265656 130534 265668
rect 147030 265656 147036 265668
rect 130528 265628 147036 265656
rect 130528 265616 130534 265628
rect 147030 265616 147036 265628
rect 147088 265616 147094 265668
rect 266722 265616 266728 265668
rect 266780 265656 266786 265668
rect 280154 265656 280160 265668
rect 266780 265628 280160 265656
rect 266780 265616 266786 265628
rect 280154 265616 280160 265628
rect 280212 265616 280218 265668
rect 52270 265004 52276 265056
rect 52328 265044 52334 265056
rect 54846 265044 54852 265056
rect 52328 265016 54852 265044
rect 52328 265004 52334 265016
rect 54846 265004 54852 265016
rect 54904 265004 54910 265056
rect 163498 265004 163504 265056
rect 163556 265044 163562 265056
rect 190822 265044 190828 265056
rect 163556 265016 190828 265044
rect 163556 265004 163562 265016
rect 190822 265004 190828 265016
rect 190880 265004 190886 265056
rect 64782 264936 64788 264988
rect 64840 264976 64846 264988
rect 66530 264976 66536 264988
rect 64840 264948 66536 264976
rect 64840 264936 64846 264948
rect 66530 264936 66536 264948
rect 66588 264936 66594 264988
rect 100754 264936 100760 264988
rect 100812 264976 100818 264988
rect 138842 264976 138848 264988
rect 100812 264948 138848 264976
rect 100812 264936 100818 264948
rect 138842 264936 138848 264948
rect 138900 264936 138906 264988
rect 157978 264936 157984 264988
rect 158036 264976 158042 264988
rect 191650 264976 191656 264988
rect 158036 264948 191656 264976
rect 158036 264936 158042 264948
rect 191650 264936 191656 264948
rect 191708 264936 191714 264988
rect 255498 264936 255504 264988
rect 255556 264976 255562 264988
rect 266446 264976 266452 264988
rect 255556 264948 266452 264976
rect 255556 264936 255562 264948
rect 266446 264936 266452 264948
rect 266504 264976 266510 264988
rect 266722 264976 266728 264988
rect 266504 264948 266728 264976
rect 266504 264936 266510 264948
rect 266722 264936 266728 264948
rect 266780 264936 266786 264988
rect 147674 264868 147680 264920
rect 147732 264908 147738 264920
rect 148962 264908 148968 264920
rect 147732 264880 148968 264908
rect 147732 264868 147738 264880
rect 148962 264868 148968 264880
rect 149020 264908 149026 264920
rect 181530 264908 181536 264920
rect 149020 264880 181536 264908
rect 149020 264868 149026 264880
rect 181530 264868 181536 264880
rect 181588 264868 181594 264920
rect 131758 264256 131764 264308
rect 131816 264296 131822 264308
rect 151354 264296 151360 264308
rect 131816 264268 151360 264296
rect 131816 264256 131822 264268
rect 151354 264256 151360 264268
rect 151412 264256 151418 264308
rect 53650 264188 53656 264240
rect 53708 264228 53714 264240
rect 66254 264228 66260 264240
rect 53708 264200 66260 264228
rect 53708 264188 53714 264200
rect 66254 264188 66260 264200
rect 66312 264188 66318 264240
rect 100938 264188 100944 264240
rect 100996 264228 101002 264240
rect 147674 264228 147680 264240
rect 100996 264200 147680 264228
rect 100996 264188 101002 264200
rect 147674 264188 147680 264200
rect 147732 264188 147738 264240
rect 276934 264188 276940 264240
rect 276992 264228 276998 264240
rect 284570 264228 284576 264240
rect 276992 264200 284576 264228
rect 276992 264188 276998 264200
rect 284570 264188 284576 264200
rect 284628 264188 284634 264240
rect 59170 263644 59176 263696
rect 59228 263684 59234 263696
rect 66806 263684 66812 263696
rect 59228 263656 66812 263684
rect 59228 263644 59234 263656
rect 66806 263644 66812 263656
rect 66864 263644 66870 263696
rect 255314 263644 255320 263696
rect 255372 263684 255378 263696
rect 260834 263684 260840 263696
rect 255372 263656 260840 263684
rect 255372 263644 255378 263656
rect 260834 263644 260840 263656
rect 260892 263644 260898 263696
rect 100846 263576 100852 263628
rect 100904 263616 100910 263628
rect 104434 263616 104440 263628
rect 100904 263588 104440 263616
rect 100904 263576 100910 263588
rect 104434 263576 104440 263588
rect 104492 263576 104498 263628
rect 164878 263576 164884 263628
rect 164936 263616 164942 263628
rect 191650 263616 191656 263628
rect 164936 263588 191656 263616
rect 164936 263576 164942 263588
rect 191650 263576 191656 263588
rect 191708 263576 191714 263628
rect 255498 263576 255504 263628
rect 255556 263616 255562 263628
rect 276014 263616 276020 263628
rect 255556 263588 276020 263616
rect 255556 263576 255562 263588
rect 276014 263576 276020 263588
rect 276072 263616 276078 263628
rect 276934 263616 276940 263628
rect 276072 263588 276940 263616
rect 276072 263576 276078 263588
rect 276934 263576 276940 263588
rect 276992 263576 276998 263628
rect 100754 263508 100760 263560
rect 100812 263548 100818 263560
rect 145650 263548 145656 263560
rect 100812 263520 145656 263548
rect 100812 263508 100818 263520
rect 145650 263508 145656 263520
rect 145708 263508 145714 263560
rect 273346 262828 273352 262880
rect 273404 262868 273410 262880
rect 281258 262868 281264 262880
rect 273404 262840 281264 262868
rect 273404 262828 273410 262840
rect 281258 262828 281264 262840
rect 281316 262828 281322 262880
rect 256418 262284 256424 262336
rect 256476 262324 256482 262336
rect 265342 262324 265348 262336
rect 256476 262296 265348 262324
rect 256476 262284 256482 262296
rect 265342 262284 265348 262296
rect 265400 262324 265406 262336
rect 265802 262324 265808 262336
rect 265400 262296 265808 262324
rect 265400 262284 265406 262296
rect 265802 262284 265808 262296
rect 265860 262284 265866 262336
rect 7742 262216 7748 262268
rect 7800 262256 7806 262268
rect 65886 262256 65892 262268
rect 7800 262228 65892 262256
rect 7800 262216 7806 262228
rect 65886 262216 65892 262228
rect 65944 262256 65950 262268
rect 66530 262256 66536 262268
rect 65944 262228 66536 262256
rect 65944 262216 65950 262228
rect 66530 262216 66536 262228
rect 66588 262216 66594 262268
rect 167638 262216 167644 262268
rect 167696 262256 167702 262268
rect 191650 262256 191656 262268
rect 167696 262228 191656 262256
rect 167696 262216 167702 262228
rect 191650 262216 191656 262228
rect 191708 262216 191714 262268
rect 280798 262148 280804 262200
rect 280856 262188 280862 262200
rect 281258 262188 281264 262200
rect 280856 262160 281264 262188
rect 280856 262148 280862 262160
rect 281258 262148 281264 262160
rect 281316 262188 281322 262200
rect 287330 262188 287336 262200
rect 281316 262160 287336 262188
rect 281316 262148 281322 262160
rect 287330 262148 287336 262160
rect 287388 262148 287394 262200
rect 52362 261536 52368 261588
rect 52420 261576 52426 261588
rect 61010 261576 61016 261588
rect 52420 261548 61016 261576
rect 52420 261536 52426 261548
rect 61010 261536 61016 261548
rect 61068 261576 61074 261588
rect 61746 261576 61752 261588
rect 61068 261548 61752 261576
rect 61068 261536 61074 261548
rect 61746 261536 61752 261548
rect 61804 261536 61810 261588
rect 104342 261536 104348 261588
rect 104400 261576 104406 261588
rect 117958 261576 117964 261588
rect 104400 261548 117964 261576
rect 104400 261536 104406 261548
rect 117958 261536 117964 261548
rect 118016 261536 118022 261588
rect 124950 261536 124956 261588
rect 125008 261576 125014 261588
rect 169570 261576 169576 261588
rect 125008 261548 169576 261576
rect 125008 261536 125014 261548
rect 169570 261536 169576 261548
rect 169628 261576 169634 261588
rect 169628 261548 171134 261576
rect 169628 261536 169634 261548
rect 7558 261468 7564 261520
rect 7616 261508 7622 261520
rect 67082 261508 67088 261520
rect 7616 261480 67088 261508
rect 7616 261468 7622 261480
rect 67082 261468 67088 261480
rect 67140 261468 67146 261520
rect 103422 261468 103428 261520
rect 103480 261508 103486 261520
rect 106274 261508 106280 261520
rect 103480 261480 106280 261508
rect 103480 261468 103486 261480
rect 106274 261468 106280 261480
rect 106332 261468 106338 261520
rect 113082 261468 113088 261520
rect 113140 261508 113146 261520
rect 166258 261508 166264 261520
rect 113140 261480 166264 261508
rect 113140 261468 113146 261480
rect 166258 261468 166264 261480
rect 166316 261468 166322 261520
rect 171106 261508 171134 261548
rect 258718 261536 258724 261588
rect 258776 261576 258782 261588
rect 279050 261576 279056 261588
rect 258776 261548 279056 261576
rect 258776 261536 258782 261548
rect 279050 261536 279056 261548
rect 279108 261536 279114 261588
rect 182818 261508 182824 261520
rect 171106 261480 182824 261508
rect 182818 261468 182824 261480
rect 182876 261468 182882 261520
rect 256602 261468 256608 261520
rect 256660 261508 256666 261520
rect 280246 261508 280252 261520
rect 256660 261480 280252 261508
rect 256660 261468 256666 261480
rect 280246 261468 280252 261480
rect 280304 261508 280310 261520
rect 281442 261508 281448 261520
rect 280304 261480 281448 261508
rect 280304 261468 280310 261480
rect 281442 261468 281448 261480
rect 281500 261468 281506 261520
rect 178678 260856 178684 260908
rect 178736 260896 178742 260908
rect 191650 260896 191656 260908
rect 178736 260868 191656 260896
rect 178736 260856 178742 260868
rect 191650 260856 191656 260868
rect 191708 260856 191714 260908
rect 281442 260856 281448 260908
rect 281500 260896 281506 260908
rect 295334 260896 295340 260908
rect 281500 260868 295340 260896
rect 281500 260856 281506 260868
rect 295334 260856 295340 260868
rect 295392 260856 295398 260908
rect 50890 260176 50896 260228
rect 50948 260216 50954 260228
rect 65794 260216 65800 260228
rect 50948 260188 65800 260216
rect 50948 260176 50954 260188
rect 65794 260176 65800 260188
rect 65852 260216 65858 260228
rect 66530 260216 66536 260228
rect 65852 260188 66536 260216
rect 65852 260176 65858 260188
rect 66530 260176 66536 260188
rect 66588 260176 66594 260228
rect 39942 260108 39948 260160
rect 40000 260148 40006 260160
rect 60458 260148 60464 260160
rect 40000 260120 60464 260148
rect 40000 260108 40006 260120
rect 60458 260108 60464 260120
rect 60516 260108 60522 260160
rect 256602 260108 256608 260160
rect 256660 260148 256666 260160
rect 263226 260148 263232 260160
rect 256660 260120 263232 260148
rect 256660 260108 256666 260120
rect 263226 260108 263232 260120
rect 263284 260108 263290 260160
rect 285674 260108 285680 260160
rect 285732 260148 285738 260160
rect 288526 260148 288532 260160
rect 285732 260120 288532 260148
rect 285732 260108 285738 260120
rect 288526 260108 288532 260120
rect 288584 260108 288590 260160
rect 100754 259496 100760 259548
rect 100812 259536 100818 259548
rect 155402 259536 155408 259548
rect 100812 259508 155408 259536
rect 100812 259496 100818 259508
rect 155402 259496 155408 259508
rect 155460 259496 155466 259548
rect 177298 259496 177304 259548
rect 177356 259536 177362 259548
rect 191650 259536 191656 259548
rect 177356 259508 191656 259536
rect 177356 259496 177362 259508
rect 191650 259496 191656 259508
rect 191708 259496 191714 259548
rect 100846 259428 100852 259480
rect 100904 259468 100910 259480
rect 185670 259468 185676 259480
rect 100904 259440 185676 259468
rect 100904 259428 100910 259440
rect 185670 259428 185676 259440
rect 185728 259428 185734 259480
rect 258718 259428 258724 259480
rect 258776 259468 258782 259480
rect 285674 259468 285680 259480
rect 258776 259440 285680 259468
rect 258776 259428 258782 259440
rect 285674 259428 285680 259440
rect 285732 259428 285738 259480
rect 101398 259360 101404 259412
rect 101456 259400 101462 259412
rect 154482 259400 154488 259412
rect 101456 259372 154488 259400
rect 101456 259360 101462 259372
rect 154482 259360 154488 259372
rect 154540 259360 154546 259412
rect 104802 258816 104808 258868
rect 104860 258856 104866 258868
rect 111058 258856 111064 258868
rect 104860 258828 111064 258856
rect 104860 258816 104866 258828
rect 111058 258816 111064 258828
rect 111116 258816 111122 258868
rect 46842 258748 46848 258800
rect 46900 258788 46906 258800
rect 64506 258788 64512 258800
rect 46900 258760 64512 258788
rect 46900 258748 46906 258760
rect 64506 258748 64512 258760
rect 64564 258788 64570 258800
rect 66346 258788 66352 258800
rect 64564 258760 66352 258788
rect 64564 258748 64570 258760
rect 66346 258748 66352 258760
rect 66404 258748 66410 258800
rect 255958 258748 255964 258800
rect 256016 258788 256022 258800
rect 265066 258788 265072 258800
rect 256016 258760 265072 258788
rect 256016 258748 256022 258760
rect 265066 258748 265072 258760
rect 265124 258748 265130 258800
rect 41138 258680 41144 258732
rect 41196 258720 41202 258732
rect 66254 258720 66260 258732
rect 41196 258692 66260 258720
rect 41196 258680 41202 258692
rect 66254 258680 66260 258692
rect 66312 258680 66318 258732
rect 156690 258680 156696 258732
rect 156748 258720 156754 258732
rect 171870 258720 171876 258732
rect 156748 258692 171876 258720
rect 156748 258680 156754 258692
rect 171870 258680 171876 258692
rect 171928 258680 171934 258732
rect 256602 258680 256608 258732
rect 256660 258720 256666 258732
rect 271874 258720 271880 258732
rect 256660 258692 271880 258720
rect 256660 258680 256666 258692
rect 271874 258680 271880 258692
rect 271932 258680 271938 258732
rect 274726 258680 274732 258732
rect 274784 258720 274790 258732
rect 287146 258720 287152 258732
rect 274784 258692 287152 258720
rect 274784 258680 274790 258692
rect 287146 258680 287152 258692
rect 287204 258680 287210 258732
rect 265066 258612 265072 258664
rect 265124 258652 265130 258664
rect 265342 258652 265348 258664
rect 265124 258624 265348 258652
rect 265124 258612 265130 258624
rect 265342 258612 265348 258624
rect 265400 258612 265406 258664
rect 174538 258068 174544 258120
rect 174596 258108 174602 258120
rect 190454 258108 190460 258120
rect 174596 258080 190460 258108
rect 174596 258068 174602 258080
rect 190454 258068 190460 258080
rect 190512 258068 190518 258120
rect 50798 258000 50804 258052
rect 50856 258040 50862 258052
rect 66438 258040 66444 258052
rect 50856 258012 66444 258040
rect 50856 258000 50862 258012
rect 66438 258000 66444 258012
rect 66496 258000 66502 258052
rect 100754 258000 100760 258052
rect 100812 258040 100818 258052
rect 104158 258040 104164 258052
rect 100812 258012 104164 258040
rect 100812 258000 100818 258012
rect 104158 258000 104164 258012
rect 104216 258000 104222 258052
rect 256326 258000 256332 258052
rect 256384 258040 256390 258052
rect 258718 258040 258724 258052
rect 256384 258012 258724 258040
rect 256384 258000 256390 258012
rect 258718 258000 258724 258012
rect 258776 258000 258782 258052
rect 267734 258000 267740 258052
rect 267792 258040 267798 258052
rect 288618 258040 288624 258052
rect 267792 258012 288624 258040
rect 267792 258000 267798 258012
rect 288618 258000 288624 258012
rect 288676 258000 288682 258052
rect 66346 257932 66352 257984
rect 66404 257972 66410 257984
rect 68186 257972 68192 257984
rect 66404 257944 68192 257972
rect 66404 257932 66410 257944
rect 68186 257932 68192 257944
rect 68244 257932 68250 257984
rect 102042 257388 102048 257440
rect 102100 257428 102106 257440
rect 130562 257428 130568 257440
rect 102100 257400 130568 257428
rect 102100 257388 102106 257400
rect 130562 257388 130568 257400
rect 130620 257388 130626 257440
rect 256602 257388 256608 257440
rect 256660 257428 256666 257440
rect 267734 257428 267740 257440
rect 256660 257400 267740 257428
rect 256660 257388 256666 257400
rect 267734 257388 267740 257400
rect 267792 257388 267798 257440
rect 44082 257320 44088 257372
rect 44140 257360 44146 257372
rect 50798 257360 50804 257372
rect 44140 257332 50804 257360
rect 44140 257320 44146 257332
rect 50798 257320 50804 257332
rect 50856 257320 50862 257372
rect 113910 257320 113916 257372
rect 113968 257360 113974 257372
rect 184290 257360 184296 257372
rect 113968 257332 184296 257360
rect 113968 257320 113974 257332
rect 184290 257320 184296 257332
rect 184348 257320 184354 257372
rect 258166 257320 258172 257372
rect 258224 257360 258230 257372
rect 286226 257360 286232 257372
rect 258224 257332 286232 257360
rect 258224 257320 258230 257332
rect 286226 257320 286232 257332
rect 286284 257320 286290 257372
rect 175918 256708 175924 256760
rect 175976 256748 175982 256760
rect 191650 256748 191656 256760
rect 175976 256720 191656 256748
rect 175976 256708 175982 256720
rect 191650 256708 191656 256720
rect 191708 256708 191714 256760
rect 286226 256708 286232 256760
rect 286284 256748 286290 256760
rect 287146 256748 287152 256760
rect 286284 256720 287152 256748
rect 286284 256708 286290 256720
rect 287146 256708 287152 256720
rect 287204 256708 287210 256760
rect 286318 256640 286324 256692
rect 286376 256680 286382 256692
rect 580902 256680 580908 256692
rect 286376 256652 580908 256680
rect 286376 256640 286382 256652
rect 580902 256640 580908 256652
rect 580960 256640 580966 256692
rect 184198 256164 184204 256216
rect 184256 256204 184262 256216
rect 192662 256204 192668 256216
rect 184256 256176 192668 256204
rect 184256 256164 184262 256176
rect 192662 256164 192668 256176
rect 192720 256164 192726 256216
rect 41230 255960 41236 256012
rect 41288 256000 41294 256012
rect 53466 256000 53472 256012
rect 41288 255972 53472 256000
rect 41288 255960 41294 255972
rect 53466 255960 53472 255972
rect 53524 256000 53530 256012
rect 59998 256000 60004 256012
rect 53524 255972 60004 256000
rect 53524 255960 53530 255972
rect 59998 255960 60004 255972
rect 60056 255960 60062 256012
rect 100846 255960 100852 256012
rect 100904 256000 100910 256012
rect 178862 256000 178868 256012
rect 100904 255972 178868 256000
rect 100904 255960 100910 255972
rect 178862 255960 178868 255972
rect 178920 255960 178926 256012
rect 256602 255960 256608 256012
rect 256660 256000 256666 256012
rect 276382 256000 276388 256012
rect 256660 255972 276388 256000
rect 256660 255960 256666 255972
rect 276382 255960 276388 255972
rect 276440 256000 276446 256012
rect 278958 256000 278964 256012
rect 276440 255972 278964 256000
rect 276440 255960 276446 255972
rect 278958 255960 278964 255972
rect 279016 255960 279022 256012
rect 278038 255824 278044 255876
rect 278096 255864 278102 255876
rect 285674 255864 285680 255876
rect 278096 255836 285680 255864
rect 278096 255824 278102 255836
rect 285674 255824 285680 255836
rect 285732 255824 285738 255876
rect 63126 255416 63132 255468
rect 63184 255456 63190 255468
rect 66254 255456 66260 255468
rect 63184 255428 66260 255456
rect 63184 255416 63190 255428
rect 66254 255416 66260 255428
rect 66312 255416 66318 255468
rect 100754 255280 100760 255332
rect 100812 255320 100818 255332
rect 164970 255320 164976 255332
rect 100812 255292 164976 255320
rect 100812 255280 100818 255292
rect 164970 255280 164976 255292
rect 165028 255280 165034 255332
rect 180150 255280 180156 255332
rect 180208 255320 180214 255332
rect 190638 255320 190644 255332
rect 180208 255292 190644 255320
rect 180208 255280 180214 255292
rect 190638 255280 190644 255292
rect 190696 255280 190702 255332
rect 256602 255280 256608 255332
rect 256660 255320 256666 255332
rect 262490 255320 262496 255332
rect 256660 255292 262496 255320
rect 256660 255280 256666 255292
rect 262490 255280 262496 255292
rect 262548 255280 262554 255332
rect 48130 255212 48136 255264
rect 48188 255252 48194 255264
rect 66806 255252 66812 255264
rect 48188 255224 66812 255252
rect 48188 255212 48194 255224
rect 66806 255212 66812 255224
rect 66864 255212 66870 255264
rect 137462 255212 137468 255264
rect 137520 255252 137526 255264
rect 177574 255252 177580 255264
rect 137520 255224 177580 255252
rect 137520 255212 137526 255224
rect 177574 255212 177580 255224
rect 177632 255212 177638 255264
rect 2774 255144 2780 255196
rect 2832 255184 2838 255196
rect 4798 255184 4804 255196
rect 2832 255156 4804 255184
rect 2832 255144 2838 255156
rect 4798 255144 4804 255156
rect 4856 255144 4862 255196
rect 100754 254872 100760 254924
rect 100812 254912 100818 254924
rect 104250 254912 104256 254924
rect 100812 254884 104256 254912
rect 100812 254872 100818 254884
rect 104250 254872 104256 254884
rect 104308 254872 104314 254924
rect 256602 254600 256608 254652
rect 256660 254640 256666 254652
rect 274726 254640 274732 254652
rect 256660 254612 274732 254640
rect 256660 254600 256666 254612
rect 274726 254600 274732 254612
rect 274784 254600 274790 254652
rect 59998 254532 60004 254584
rect 60056 254572 60062 254584
rect 66806 254572 66812 254584
rect 60056 254544 66812 254572
rect 60056 254532 60062 254544
rect 66806 254532 66812 254544
rect 66864 254532 66870 254584
rect 115290 254532 115296 254584
rect 115348 254572 115354 254584
rect 137462 254572 137468 254584
rect 115348 254544 137468 254572
rect 115348 254532 115354 254544
rect 137462 254532 137468 254544
rect 137520 254532 137526 254584
rect 171042 254532 171048 254584
rect 171100 254572 171106 254584
rect 176010 254572 176016 254584
rect 171100 254544 176016 254572
rect 171100 254532 171106 254544
rect 176010 254532 176016 254544
rect 176068 254532 176074 254584
rect 259362 254532 259368 254584
rect 259420 254572 259426 254584
rect 289906 254572 289912 254584
rect 259420 254544 289912 254572
rect 259420 254532 259426 254544
rect 289906 254532 289912 254544
rect 289964 254532 289970 254584
rect 185578 253988 185584 254040
rect 185636 254028 185642 254040
rect 191650 254028 191656 254040
rect 185636 254000 191656 254028
rect 185636 253988 185642 254000
rect 191650 253988 191656 254000
rect 191708 253988 191714 254040
rect 46842 253920 46848 253972
rect 46900 253960 46906 253972
rect 48130 253960 48136 253972
rect 46900 253932 48136 253960
rect 46900 253920 46906 253932
rect 48130 253920 48136 253932
rect 48188 253920 48194 253972
rect 100754 253920 100760 253972
rect 100812 253960 100818 253972
rect 115198 253960 115204 253972
rect 100812 253932 115204 253960
rect 100812 253920 100818 253932
rect 115198 253920 115204 253932
rect 115256 253920 115262 253972
rect 182818 253920 182824 253972
rect 182876 253960 182882 253972
rect 191558 253960 191564 253972
rect 182876 253932 191564 253960
rect 182876 253920 182882 253932
rect 191558 253920 191564 253932
rect 191616 253920 191622 253972
rect 111058 253240 111064 253292
rect 111116 253280 111122 253292
rect 122190 253280 122196 253292
rect 111116 253252 122196 253280
rect 111116 253240 111122 253252
rect 122190 253240 122196 253252
rect 122248 253240 122254 253292
rect 7650 253172 7656 253224
rect 7708 253212 7714 253224
rect 66990 253212 66996 253224
rect 7708 253184 66996 253212
rect 7708 253172 7714 253184
rect 66990 253172 66996 253184
rect 67048 253212 67054 253224
rect 67358 253212 67364 253224
rect 67048 253184 67364 253212
rect 67048 253172 67054 253184
rect 67358 253172 67364 253184
rect 67416 253172 67422 253224
rect 108390 253172 108396 253224
rect 108448 253212 108454 253224
rect 123570 253212 123576 253224
rect 108448 253184 123576 253212
rect 108448 253172 108454 253184
rect 123570 253172 123576 253184
rect 123628 253172 123634 253224
rect 138658 253172 138664 253224
rect 138716 253212 138722 253224
rect 162302 253212 162308 253224
rect 138716 253184 162308 253212
rect 138716 253172 138722 253184
rect 162302 253172 162308 253184
rect 162360 253172 162366 253224
rect 254118 253036 254124 253088
rect 254176 253076 254182 253088
rect 259362 253076 259368 253088
rect 254176 253048 259368 253076
rect 254176 253036 254182 253048
rect 259362 253036 259368 253048
rect 259420 253036 259426 253088
rect 158162 252764 158168 252816
rect 158220 252804 158226 252816
rect 161014 252804 161020 252816
rect 158220 252776 161020 252804
rect 158220 252764 158226 252776
rect 161014 252764 161020 252776
rect 161072 252764 161078 252816
rect 100754 252560 100760 252612
rect 100812 252600 100818 252612
rect 111150 252600 111156 252612
rect 100812 252572 111156 252600
rect 100812 252560 100818 252572
rect 111150 252560 111156 252572
rect 111208 252560 111214 252612
rect 170398 252560 170404 252612
rect 170456 252600 170462 252612
rect 191650 252600 191656 252612
rect 170456 252572 191656 252600
rect 170456 252560 170462 252572
rect 191650 252560 191656 252572
rect 191708 252560 191714 252612
rect 255774 252560 255780 252612
rect 255832 252600 255838 252612
rect 258350 252600 258356 252612
rect 255832 252572 258356 252600
rect 255832 252560 255838 252572
rect 258350 252560 258356 252572
rect 258408 252560 258414 252612
rect 273346 252560 273352 252612
rect 273404 252600 273410 252612
rect 275278 252600 275284 252612
rect 273404 252572 275284 252600
rect 273404 252560 273410 252572
rect 275278 252560 275284 252572
rect 275336 252560 275342 252612
rect 100846 252492 100852 252544
rect 100904 252532 100910 252544
rect 119338 252532 119344 252544
rect 100904 252504 119344 252532
rect 100904 252492 100910 252504
rect 119338 252492 119344 252504
rect 119396 252492 119402 252544
rect 116762 251880 116768 251932
rect 116820 251920 116826 251932
rect 158162 251920 158168 251932
rect 116820 251892 158168 251920
rect 116820 251880 116826 251892
rect 158162 251880 158168 251892
rect 158220 251880 158226 251932
rect 55030 251812 55036 251864
rect 55088 251852 55094 251864
rect 66070 251852 66076 251864
rect 55088 251824 66076 251852
rect 55088 251812 55094 251824
rect 66070 251812 66076 251824
rect 66128 251852 66134 251864
rect 66622 251852 66628 251864
rect 66128 251824 66628 251852
rect 66128 251812 66134 251824
rect 66622 251812 66628 251824
rect 66680 251812 66686 251864
rect 129182 251812 129188 251864
rect 129240 251852 129246 251864
rect 180242 251852 180248 251864
rect 129240 251824 180248 251852
rect 129240 251812 129246 251824
rect 180242 251812 180248 251824
rect 180300 251852 180306 251864
rect 189810 251852 189816 251864
rect 180300 251824 189816 251852
rect 180300 251812 180306 251824
rect 189810 251812 189816 251824
rect 189868 251812 189874 251864
rect 190362 251812 190368 251864
rect 190420 251852 190426 251864
rect 193214 251852 193220 251864
rect 190420 251824 193220 251852
rect 190420 251812 190426 251824
rect 193214 251812 193220 251824
rect 193272 251812 193278 251864
rect 270402 251812 270408 251864
rect 270460 251852 270466 251864
rect 582466 251852 582472 251864
rect 270460 251824 582472 251852
rect 270460 251812 270466 251824
rect 582466 251812 582472 251824
rect 582524 251812 582530 251864
rect 100754 251336 100760 251388
rect 100812 251376 100818 251388
rect 103514 251376 103520 251388
rect 100812 251348 103520 251376
rect 100812 251336 100818 251348
rect 103514 251336 103520 251348
rect 103572 251336 103578 251388
rect 256418 251268 256424 251320
rect 256476 251308 256482 251320
rect 269390 251308 269396 251320
rect 256476 251280 269396 251308
rect 256476 251268 256482 251280
rect 269390 251268 269396 251280
rect 269448 251308 269454 251320
rect 270402 251308 270408 251320
rect 269448 251280 270408 251308
rect 269448 251268 269454 251280
rect 270402 251268 270408 251280
rect 270460 251268 270466 251320
rect 166258 251200 166264 251252
rect 166316 251240 166322 251252
rect 191650 251240 191656 251252
rect 166316 251212 191656 251240
rect 166316 251200 166322 251212
rect 191650 251200 191656 251212
rect 191708 251200 191714 251252
rect 256602 251200 256608 251252
rect 256660 251240 256666 251252
rect 271874 251240 271880 251252
rect 256660 251212 271880 251240
rect 256660 251200 256666 251212
rect 271874 251200 271880 251212
rect 271932 251200 271938 251252
rect 60550 250724 60556 250776
rect 60608 250764 60614 250776
rect 66806 250764 66812 250776
rect 60608 250736 66812 250764
rect 60608 250724 60614 250736
rect 66806 250724 66812 250736
rect 66864 250724 66870 250776
rect 100754 250520 100760 250572
rect 100812 250560 100818 250572
rect 106918 250560 106924 250572
rect 100812 250532 106924 250560
rect 100812 250520 100818 250532
rect 106918 250520 106924 250532
rect 106976 250520 106982 250572
rect 102778 250452 102784 250504
rect 102836 250492 102842 250504
rect 153838 250492 153844 250504
rect 102836 250464 153844 250492
rect 102836 250452 102842 250464
rect 153838 250452 153844 250464
rect 153896 250452 153902 250504
rect 256602 250452 256608 250504
rect 256660 250492 256666 250504
rect 273346 250492 273352 250504
rect 256660 250464 273352 250492
rect 256660 250452 256666 250464
rect 273346 250452 273352 250464
rect 273404 250452 273410 250504
rect 256694 250316 256700 250368
rect 256752 250356 256758 250368
rect 257338 250356 257344 250368
rect 256752 250328 257344 250356
rect 256752 250316 256758 250328
rect 257338 250316 257344 250328
rect 257396 250316 257402 250368
rect 169018 249772 169024 249824
rect 169076 249812 169082 249824
rect 190638 249812 190644 249824
rect 169076 249784 190644 249812
rect 169076 249772 169082 249784
rect 190638 249772 190644 249784
rect 190696 249772 190702 249824
rect 100938 249704 100944 249756
rect 100996 249744 101002 249756
rect 108482 249744 108488 249756
rect 100996 249716 108488 249744
rect 100996 249704 101002 249716
rect 108482 249704 108488 249716
rect 108540 249744 108546 249756
rect 108942 249744 108948 249756
rect 108540 249716 108948 249744
rect 108540 249704 108546 249716
rect 108942 249704 108948 249716
rect 109000 249704 109006 249756
rect 162118 249704 162124 249756
rect 162176 249744 162182 249756
rect 163682 249744 163688 249756
rect 162176 249716 163688 249744
rect 162176 249704 162182 249716
rect 163682 249704 163688 249716
rect 163740 249704 163746 249756
rect 108482 249092 108488 249144
rect 108540 249132 108546 249144
rect 129090 249132 129096 249144
rect 108540 249104 129096 249132
rect 108540 249092 108546 249104
rect 129090 249092 129096 249104
rect 129148 249132 129154 249144
rect 148502 249132 148508 249144
rect 129148 249104 148508 249132
rect 129148 249092 129154 249104
rect 148502 249092 148508 249104
rect 148560 249092 148566 249144
rect 120810 249024 120816 249076
rect 120868 249064 120874 249076
rect 160830 249064 160836 249076
rect 120868 249036 160836 249064
rect 120868 249024 120874 249036
rect 160830 249024 160836 249036
rect 160888 249024 160894 249076
rect 256602 248480 256608 248532
rect 256660 248520 256666 248532
rect 278038 248520 278044 248532
rect 256660 248492 278044 248520
rect 256660 248480 256666 248492
rect 278038 248480 278044 248492
rect 278096 248480 278102 248532
rect 53374 248412 53380 248464
rect 53432 248452 53438 248464
rect 57882 248452 57888 248464
rect 53432 248424 57888 248452
rect 53432 248412 53438 248424
rect 57882 248412 57888 248424
rect 57940 248452 57946 248464
rect 66806 248452 66812 248464
rect 57940 248424 66812 248452
rect 57940 248412 57946 248424
rect 66806 248412 66812 248424
rect 66864 248412 66870 248464
rect 188338 248412 188344 248464
rect 188396 248452 188402 248464
rect 190822 248452 190828 248464
rect 188396 248424 190828 248452
rect 188396 248412 188402 248424
rect 190822 248412 190828 248424
rect 190880 248412 190886 248464
rect 256234 248412 256240 248464
rect 256292 248452 256298 248464
rect 291286 248452 291292 248464
rect 256292 248424 291292 248452
rect 256292 248412 256298 248424
rect 291286 248412 291292 248424
rect 291344 248452 291350 248464
rect 582374 248452 582380 248464
rect 291344 248424 582380 248452
rect 291344 248412 291350 248424
rect 582374 248412 582380 248424
rect 582432 248412 582438 248464
rect 254670 248344 254676 248396
rect 254728 248384 254734 248396
rect 286318 248384 286324 248396
rect 254728 248356 286324 248384
rect 254728 248344 254734 248356
rect 286318 248344 286324 248356
rect 286376 248344 286382 248396
rect 135162 247664 135168 247716
rect 135220 247704 135226 247716
rect 167822 247704 167828 247716
rect 135220 247676 167828 247704
rect 135220 247664 135226 247676
rect 167822 247664 167828 247676
rect 167880 247664 167886 247716
rect 60550 247052 60556 247104
rect 60608 247092 60614 247104
rect 66530 247092 66536 247104
rect 60608 247064 66536 247092
rect 60608 247052 60614 247064
rect 66530 247052 66536 247064
rect 66588 247052 66594 247104
rect 104802 247092 104808 247104
rect 103486 247064 104808 247092
rect 100938 246984 100944 247036
rect 100996 247024 101002 247036
rect 103486 247024 103514 247064
rect 104802 247052 104808 247064
rect 104860 247092 104866 247104
rect 133874 247092 133880 247104
rect 104860 247064 133880 247092
rect 104860 247052 104866 247064
rect 133874 247052 133880 247064
rect 133932 247092 133938 247104
rect 135162 247092 135168 247104
rect 133932 247064 135168 247092
rect 133932 247052 133938 247064
rect 135162 247052 135168 247064
rect 135220 247052 135226 247104
rect 100996 246996 103514 247024
rect 100996 246984 101002 246996
rect 256602 246984 256608 247036
rect 256660 247024 256666 247036
rect 283006 247024 283012 247036
rect 256660 246996 283012 247024
rect 256660 246984 256666 246996
rect 283006 246984 283012 246996
rect 283064 247024 283070 247036
rect 288526 247024 288532 247036
rect 283064 246996 288532 247024
rect 283064 246984 283070 246996
rect 288526 246984 288532 246996
rect 288584 246984 288590 247036
rect 102318 246304 102324 246356
rect 102376 246344 102382 246356
rect 155954 246344 155960 246356
rect 102376 246316 155960 246344
rect 102376 246304 102382 246316
rect 155954 246304 155960 246316
rect 156012 246344 156018 246356
rect 162762 246344 162768 246356
rect 156012 246316 162768 246344
rect 156012 246304 156018 246316
rect 162762 246304 162768 246316
rect 162820 246304 162826 246356
rect 168282 246304 168288 246356
rect 168340 246344 168346 246356
rect 175274 246344 175280 246356
rect 168340 246316 175280 246344
rect 168340 246304 168346 246316
rect 175274 246304 175280 246316
rect 175332 246304 175338 246356
rect 186222 246304 186228 246356
rect 186280 246344 186286 246356
rect 193582 246344 193588 246356
rect 186280 246316 193588 246344
rect 186280 246304 186286 246316
rect 193582 246304 193588 246316
rect 193640 246304 193646 246356
rect 253934 246032 253940 246084
rect 253992 246072 253998 246084
rect 258166 246072 258172 246084
rect 253992 246044 258172 246072
rect 253992 246032 253998 246044
rect 258166 246032 258172 246044
rect 258224 246032 258230 246084
rect 183462 245664 183468 245676
rect 183375 245636 183468 245664
rect 183462 245624 183468 245636
rect 183520 245664 183526 245676
rect 191282 245664 191288 245676
rect 183520 245636 191288 245664
rect 183520 245624 183526 245636
rect 191282 245624 191288 245636
rect 191340 245624 191346 245676
rect 159542 245556 159548 245608
rect 159600 245596 159606 245608
rect 183480 245596 183508 245624
rect 159600 245568 183508 245596
rect 159600 245556 159606 245568
rect 190270 245556 190276 245608
rect 190328 245596 190334 245608
rect 191834 245596 191840 245608
rect 190328 245568 191840 245596
rect 190328 245556 190334 245568
rect 191834 245556 191840 245568
rect 191892 245556 191898 245608
rect 100938 244944 100944 244996
rect 100996 244984 101002 244996
rect 106274 244984 106280 244996
rect 100996 244956 106280 244984
rect 100996 244944 101002 244956
rect 106274 244944 106280 244956
rect 106332 244984 106338 244996
rect 107010 244984 107016 244996
rect 106332 244956 107016 244984
rect 106332 244944 106338 244956
rect 107010 244944 107016 244956
rect 107068 244944 107074 244996
rect 101030 244876 101036 244928
rect 101088 244916 101094 244928
rect 165614 244916 165620 244928
rect 101088 244888 165620 244916
rect 101088 244876 101094 244888
rect 165614 244876 165620 244888
rect 165672 244876 165678 244928
rect 58894 244264 58900 244316
rect 58952 244304 58958 244316
rect 66806 244304 66812 244316
rect 58952 244276 66812 244304
rect 58952 244264 58958 244276
rect 66806 244264 66812 244276
rect 66864 244264 66870 244316
rect 165614 244264 165620 244316
rect 165672 244304 165678 244316
rect 166442 244304 166448 244316
rect 165672 244276 166448 244304
rect 165672 244264 165678 244276
rect 166442 244264 166448 244276
rect 166500 244264 166506 244316
rect 56502 244196 56508 244248
rect 56560 244236 56566 244248
rect 66714 244236 66720 244248
rect 56560 244208 66720 244236
rect 56560 244196 56566 244208
rect 66714 244196 66720 244208
rect 66772 244196 66778 244248
rect 276382 244196 276388 244248
rect 276440 244236 276446 244248
rect 278866 244236 278872 244248
rect 276440 244208 278872 244236
rect 276440 244196 276446 244208
rect 278866 244196 278872 244208
rect 278924 244196 278930 244248
rect 113910 243584 113916 243636
rect 113968 243624 113974 243636
rect 140130 243624 140136 243636
rect 113968 243596 140136 243624
rect 113968 243584 113974 243596
rect 140130 243584 140136 243596
rect 140188 243584 140194 243636
rect 97994 243516 98000 243568
rect 98052 243556 98058 243568
rect 98270 243556 98276 243568
rect 98052 243528 98276 243556
rect 98052 243516 98058 243528
rect 98270 243516 98276 243528
rect 98328 243516 98334 243568
rect 192570 243556 192576 243568
rect 103486 243528 192576 243556
rect 98270 243380 98276 243432
rect 98328 243420 98334 243432
rect 103486 243420 103514 243528
rect 192570 243516 192576 243528
rect 192628 243516 192634 243568
rect 255314 243516 255320 243568
rect 255372 243556 255378 243568
rect 287054 243556 287060 243568
rect 255372 243528 287060 243556
rect 255372 243516 255378 243528
rect 287054 243516 287060 243528
rect 287112 243516 287118 243568
rect 98328 243392 103514 243420
rect 98328 243380 98334 243392
rect 61746 242904 61752 242956
rect 61804 242944 61810 242956
rect 66898 242944 66904 242956
rect 61804 242916 66904 242944
rect 61804 242904 61810 242916
rect 66898 242904 66904 242916
rect 66956 242904 66962 242956
rect 162762 242904 162768 242956
rect 162820 242944 162826 242956
rect 192110 242944 192116 242956
rect 162820 242916 192116 242944
rect 162820 242904 162826 242916
rect 192110 242904 192116 242916
rect 192168 242904 192174 242956
rect 192478 242904 192484 242956
rect 192536 242944 192542 242956
rect 252830 242944 252836 242956
rect 192536 242916 195836 242944
rect 192536 242904 192542 242916
rect 67726 242496 67732 242548
rect 67784 242536 67790 242548
rect 68784 242536 68790 242548
rect 67784 242508 68790 242536
rect 67784 242496 67790 242508
rect 68784 242496 68790 242508
rect 68842 242496 68848 242548
rect 112530 242224 112536 242276
rect 112588 242264 112594 242276
rect 145742 242264 145748 242276
rect 112588 242236 145748 242264
rect 112588 242224 112594 242236
rect 145742 242224 145748 242236
rect 145800 242224 145806 242276
rect 134702 242156 134708 242208
rect 134760 242196 134766 242208
rect 134760 242168 180794 242196
rect 134760 242156 134766 242168
rect 180766 242060 180794 242168
rect 195808 242072 195836 242916
rect 248524 242916 252836 242944
rect 248524 242072 248552 242916
rect 252830 242904 252836 242916
rect 252888 242904 252894 242956
rect 255682 242904 255688 242956
rect 255740 242944 255746 242956
rect 276382 242944 276388 242956
rect 255740 242916 276388 242944
rect 255740 242904 255746 242916
rect 276382 242904 276388 242916
rect 276440 242944 276446 242956
rect 276658 242944 276664 242956
rect 276440 242916 276664 242944
rect 276440 242904 276446 242916
rect 276658 242904 276664 242916
rect 276716 242904 276722 242956
rect 252370 242292 252376 242344
rect 252428 242332 252434 242344
rect 252830 242332 252836 242344
rect 252428 242304 252836 242332
rect 252428 242292 252434 242304
rect 252830 242292 252836 242304
rect 252888 242292 252894 242344
rect 259638 242196 259644 242208
rect 250456 242168 259644 242196
rect 250456 242072 250484 242168
rect 259638 242156 259644 242168
rect 259696 242156 259702 242208
rect 195330 242060 195336 242072
rect 180766 242032 195336 242060
rect 195330 242020 195336 242032
rect 195388 242020 195394 242072
rect 195790 242020 195796 242072
rect 195848 242020 195854 242072
rect 248506 242020 248512 242072
rect 248564 242020 248570 242072
rect 250438 242020 250444 242072
rect 250496 242020 250502 242072
rect 155310 241884 155316 241936
rect 155368 241924 155374 241936
rect 160738 241924 160744 241936
rect 155368 241896 160744 241924
rect 155368 241884 155374 241896
rect 160738 241884 160744 241896
rect 160796 241884 160802 241936
rect 68554 241748 68560 241800
rect 68612 241788 68618 241800
rect 69382 241788 69388 241800
rect 68612 241760 69388 241788
rect 68612 241748 68618 241760
rect 69382 241748 69388 241760
rect 69440 241748 69446 241800
rect 94958 241612 94964 241664
rect 95016 241652 95022 241664
rect 115290 241652 115296 241664
rect 95016 241624 115296 241652
rect 95016 241612 95022 241624
rect 115290 241612 115296 241624
rect 115348 241612 115354 241664
rect 59262 241544 59268 241596
rect 59320 241584 59326 241596
rect 66806 241584 66812 241596
rect 59320 241556 66812 241584
rect 59320 241544 59326 241556
rect 66806 241544 66812 241556
rect 66864 241544 66870 241596
rect 58986 241476 58992 241528
rect 59044 241516 59050 241528
rect 77432 241516 77438 241528
rect 59044 241488 77438 241516
rect 59044 241476 59050 241488
rect 77432 241476 77438 241488
rect 77490 241476 77496 241528
rect 93946 241476 93952 241528
rect 94004 241516 94010 241528
rect 94976 241516 95004 241612
rect 94004 241488 95004 241516
rect 94004 241476 94010 241488
rect 95970 241476 95976 241528
rect 96028 241516 96034 241528
rect 99098 241516 99104 241528
rect 96028 241488 99104 241516
rect 96028 241476 96034 241488
rect 99098 241476 99104 241488
rect 99156 241476 99162 241528
rect 181990 241476 181996 241528
rect 182048 241516 182054 241528
rect 201494 241516 201500 241528
rect 182048 241488 201500 241516
rect 182048 241476 182054 241488
rect 201494 241476 201500 241488
rect 201552 241516 201558 241528
rect 201954 241516 201960 241528
rect 201552 241488 201960 241516
rect 201552 241476 201558 241488
rect 201954 241476 201960 241488
rect 202012 241476 202018 241528
rect 255498 241476 255504 241528
rect 255556 241516 255562 241528
rect 261110 241516 261116 241528
rect 255556 241488 261116 241516
rect 255556 241476 255562 241488
rect 261110 241476 261116 241488
rect 261168 241476 261174 241528
rect 73522 241408 73528 241460
rect 73580 241448 73586 241460
rect 112622 241448 112628 241460
rect 73580 241420 112628 241448
rect 73580 241408 73586 241420
rect 112622 241408 112628 241420
rect 112680 241408 112686 241460
rect 192110 241408 192116 241460
rect 192168 241448 192174 241460
rect 204346 241448 204352 241460
rect 192168 241420 204352 241448
rect 192168 241408 192174 241420
rect 204346 241408 204352 241420
rect 204404 241408 204410 241460
rect 268286 241408 268292 241460
rect 268344 241448 268350 241460
rect 298094 241448 298100 241460
rect 268344 241420 298100 241448
rect 268344 241408 268350 241420
rect 298094 241408 298100 241420
rect 298152 241408 298158 241460
rect 67818 241340 67824 241392
rect 67876 241380 67882 241392
rect 102318 241380 102324 241392
rect 67876 241352 102324 241380
rect 67876 241340 67882 241352
rect 102318 241340 102324 241352
rect 102376 241340 102382 241392
rect 3418 241068 3424 241120
rect 3476 241108 3482 241120
rect 7742 241108 7748 241120
rect 3476 241080 7748 241108
rect 3476 241068 3482 241080
rect 7742 241068 7748 241080
rect 7800 241068 7806 241120
rect 136082 240796 136088 240848
rect 136140 240836 136146 240848
rect 171134 240836 171140 240848
rect 136140 240808 171140 240836
rect 136140 240796 136146 240808
rect 171134 240796 171140 240808
rect 171192 240796 171198 240848
rect 234614 240836 234620 240848
rect 219406 240808 234620 240836
rect 164970 240728 164976 240780
rect 165028 240768 165034 240780
rect 219406 240768 219434 240808
rect 234614 240796 234620 240808
rect 234672 240836 234678 240848
rect 256694 240836 256700 240848
rect 234672 240808 256700 240836
rect 234672 240796 234678 240808
rect 256694 240796 256700 240808
rect 256752 240796 256758 240848
rect 165028 240740 219434 240768
rect 165028 240728 165034 240740
rect 251818 240728 251824 240780
rect 251876 240768 251882 240780
rect 276750 240768 276756 240780
rect 251876 240740 276756 240768
rect 251876 240728 251882 240740
rect 276750 240728 276756 240740
rect 276808 240728 276814 240780
rect 181530 240320 181536 240372
rect 181588 240360 181594 240372
rect 186314 240360 186320 240372
rect 181588 240332 186320 240360
rect 181588 240320 181594 240332
rect 186314 240320 186320 240332
rect 186372 240320 186378 240372
rect 74534 240116 74540 240168
rect 74592 240156 74598 240168
rect 75454 240156 75460 240168
rect 74592 240128 75460 240156
rect 74592 240116 74598 240128
rect 75454 240116 75460 240128
rect 75512 240116 75518 240168
rect 78674 240116 78680 240168
rect 78732 240156 78738 240168
rect 79318 240156 79324 240168
rect 78732 240128 79324 240156
rect 78732 240116 78738 240128
rect 79318 240116 79324 240128
rect 79376 240116 79382 240168
rect 80054 240116 80060 240168
rect 80112 240156 80118 240168
rect 80974 240156 80980 240168
rect 80112 240128 80980 240156
rect 80112 240116 80118 240128
rect 80974 240116 80980 240128
rect 81032 240116 81038 240168
rect 82814 240116 82820 240168
rect 82872 240156 82878 240168
rect 83734 240156 83740 240168
rect 82872 240128 83740 240156
rect 82872 240116 82878 240128
rect 83734 240116 83740 240128
rect 83792 240116 83798 240168
rect 84194 240116 84200 240168
rect 84252 240156 84258 240168
rect 84838 240156 84844 240168
rect 84252 240128 84844 240156
rect 84252 240116 84258 240128
rect 84838 240116 84844 240128
rect 84896 240116 84902 240168
rect 86954 240116 86960 240168
rect 87012 240156 87018 240168
rect 87598 240156 87604 240168
rect 87012 240128 87604 240156
rect 87012 240116 87018 240128
rect 87598 240116 87604 240128
rect 87656 240116 87662 240168
rect 95234 240116 95240 240168
rect 95292 240156 95298 240168
rect 95878 240156 95884 240168
rect 95292 240128 95884 240156
rect 95292 240116 95298 240128
rect 95878 240116 95884 240128
rect 95936 240116 95942 240168
rect 96614 240116 96620 240168
rect 96672 240156 96678 240168
rect 97626 240156 97632 240168
rect 96672 240128 97632 240156
rect 96672 240116 96678 240128
rect 97626 240116 97632 240128
rect 97684 240116 97690 240168
rect 65978 240048 65984 240100
rect 66036 240088 66042 240100
rect 70394 240088 70400 240100
rect 66036 240060 70400 240088
rect 66036 240048 66042 240060
rect 70394 240048 70400 240060
rect 70452 240048 70458 240100
rect 76098 240048 76104 240100
rect 76156 240088 76162 240100
rect 77478 240088 77484 240100
rect 76156 240060 77484 240088
rect 76156 240048 76162 240060
rect 77478 240048 77484 240060
rect 77536 240048 77542 240100
rect 82170 240048 82176 240100
rect 82228 240088 82234 240100
rect 86862 240088 86868 240100
rect 82228 240060 86868 240088
rect 82228 240048 82234 240060
rect 86862 240048 86868 240060
rect 86920 240048 86926 240100
rect 89622 240048 89628 240100
rect 89680 240088 89686 240100
rect 182174 240088 182180 240100
rect 89680 240060 182180 240088
rect 89680 240048 89686 240060
rect 182174 240048 182180 240060
rect 182232 240088 182238 240100
rect 211798 240088 211804 240100
rect 182232 240060 211804 240088
rect 182232 240048 182238 240060
rect 211798 240048 211804 240060
rect 211856 240048 211862 240100
rect 233878 240048 233884 240100
rect 233936 240088 233942 240100
rect 234614 240088 234620 240100
rect 233936 240060 234620 240088
rect 233936 240048 233942 240060
rect 234614 240048 234620 240060
rect 234672 240048 234678 240100
rect 242158 240048 242164 240100
rect 242216 240088 242222 240100
rect 242710 240088 242716 240100
rect 242216 240060 242716 240088
rect 242216 240048 242222 240060
rect 242710 240048 242716 240060
rect 242768 240088 242774 240100
rect 272058 240088 272064 240100
rect 242768 240060 272064 240088
rect 242768 240048 242774 240060
rect 272058 240048 272064 240060
rect 272116 240048 272122 240100
rect 192662 239980 192668 240032
rect 192720 240020 192726 240032
rect 196158 240020 196164 240032
rect 192720 239992 196164 240020
rect 192720 239980 192726 239992
rect 196158 239980 196164 239992
rect 196216 239980 196222 240032
rect 177942 239640 177948 239692
rect 178000 239680 178006 239692
rect 178770 239680 178776 239692
rect 178000 239652 178776 239680
rect 178000 239640 178006 239652
rect 178770 239640 178776 239652
rect 178828 239640 178834 239692
rect 219434 239640 219440 239692
rect 219492 239680 219498 239692
rect 221090 239680 221096 239692
rect 219492 239652 221096 239680
rect 219492 239640 219498 239652
rect 221090 239640 221096 239652
rect 221148 239640 221154 239692
rect 69474 239368 69480 239420
rect 69532 239408 69538 239420
rect 89070 239408 89076 239420
rect 69532 239380 89076 239408
rect 69532 239368 69538 239380
rect 89070 239368 89076 239380
rect 89128 239368 89134 239420
rect 196158 239368 196164 239420
rect 196216 239408 196222 239420
rect 206738 239408 206744 239420
rect 196216 239380 206744 239408
rect 196216 239368 196222 239380
rect 206738 239368 206744 239380
rect 206796 239368 206802 239420
rect 249058 239368 249064 239420
rect 249116 239408 249122 239420
rect 266998 239408 267004 239420
rect 249116 239380 267004 239408
rect 249116 239368 249122 239380
rect 266998 239368 267004 239380
rect 267056 239368 267062 239420
rect 89346 238756 89352 238808
rect 89404 238796 89410 238808
rect 89404 238768 93072 238796
rect 89404 238756 89410 238768
rect 93044 238728 93072 238768
rect 219434 238756 219440 238808
rect 219492 238756 219498 238808
rect 227070 238756 227076 238808
rect 227128 238796 227134 238808
rect 230750 238796 230756 238808
rect 227128 238768 230756 238796
rect 227128 238756 227134 238768
rect 230750 238756 230756 238768
rect 230808 238756 230814 238808
rect 233142 238756 233148 238808
rect 233200 238796 233206 238808
rect 237374 238796 237380 238808
rect 233200 238768 237380 238796
rect 233200 238756 233206 238768
rect 237374 238756 237380 238768
rect 237432 238756 237438 238808
rect 93762 238728 93768 238740
rect 93044 238700 93768 238728
rect 93762 238688 93768 238700
rect 93820 238728 93826 238740
rect 107654 238728 107660 238740
rect 93820 238700 107660 238728
rect 93820 238688 93826 238700
rect 107654 238688 107660 238700
rect 107712 238688 107718 238740
rect 188982 238688 188988 238740
rect 189040 238728 189046 238740
rect 219452 238728 219480 238756
rect 189040 238700 219480 238728
rect 189040 238688 189046 238700
rect 80146 238620 80152 238672
rect 80204 238660 80210 238672
rect 95970 238660 95976 238672
rect 80204 238632 95976 238660
rect 80204 238620 80210 238632
rect 95970 238620 95976 238632
rect 96028 238620 96034 238672
rect 177942 238620 177948 238672
rect 178000 238660 178006 238672
rect 209130 238660 209136 238672
rect 178000 238632 209136 238660
rect 178000 238620 178006 238632
rect 209130 238620 209136 238632
rect 209188 238620 209194 238672
rect 74350 238484 74356 238536
rect 74408 238524 74414 238536
rect 76650 238524 76656 238536
rect 74408 238496 76656 238524
rect 74408 238484 74414 238496
rect 76650 238484 76656 238496
rect 76708 238484 76714 238536
rect 170490 238076 170496 238128
rect 170548 238116 170554 238128
rect 177942 238116 177948 238128
rect 170548 238088 177948 238116
rect 170548 238076 170554 238088
rect 177942 238076 177948 238088
rect 178000 238076 178006 238128
rect 45370 238008 45376 238060
rect 45428 238048 45434 238060
rect 46750 238048 46756 238060
rect 45428 238020 46756 238048
rect 45428 238008 45434 238020
rect 46750 238008 46756 238020
rect 46808 238048 46814 238060
rect 74626 238048 74632 238060
rect 46808 238020 74632 238048
rect 46808 238008 46814 238020
rect 74626 238008 74632 238020
rect 74684 238008 74690 238060
rect 107562 238008 107568 238060
rect 107620 238048 107626 238060
rect 170582 238048 170588 238060
rect 107620 238020 170588 238048
rect 107620 238008 107626 238020
rect 170582 238008 170588 238020
rect 170640 238008 170646 238060
rect 215294 238008 215300 238060
rect 215352 238048 215358 238060
rect 261018 238048 261024 238060
rect 215352 238020 261024 238048
rect 215352 238008 215358 238020
rect 261018 238008 261024 238020
rect 261076 238008 261082 238060
rect 79410 237396 79416 237448
rect 79468 237436 79474 237448
rect 80146 237436 80152 237448
rect 79468 237408 80152 237436
rect 79468 237396 79474 237408
rect 80146 237396 80152 237408
rect 80204 237396 80210 237448
rect 95050 237396 95056 237448
rect 95108 237436 95114 237448
rect 98086 237436 98092 237448
rect 95108 237408 98092 237436
rect 95108 237396 95114 237408
rect 98086 237396 98092 237408
rect 98144 237396 98150 237448
rect 59078 237328 59084 237380
rect 59136 237368 59142 237380
rect 76098 237368 76104 237380
rect 59136 237340 76104 237368
rect 59136 237328 59142 237340
rect 76098 237328 76104 237340
rect 76156 237328 76162 237380
rect 78766 237328 78772 237380
rect 78824 237368 78830 237380
rect 108390 237368 108396 237380
rect 78824 237340 108396 237368
rect 78824 237328 78830 237340
rect 108390 237328 108396 237340
rect 108448 237328 108454 237380
rect 184750 237328 184756 237380
rect 184808 237368 184814 237380
rect 233142 237368 233148 237380
rect 184808 237340 233148 237368
rect 184808 237328 184814 237340
rect 233142 237328 233148 237340
rect 233200 237328 233206 237380
rect 252278 237328 252284 237380
rect 252336 237368 252342 237380
rect 287238 237368 287244 237380
rect 252336 237340 287244 237368
rect 252336 237328 252342 237340
rect 287238 237328 287244 237340
rect 287296 237328 287302 237380
rect 193766 237260 193772 237312
rect 193824 237300 193830 237312
rect 215478 237300 215484 237312
rect 193824 237272 215484 237300
rect 193824 237260 193830 237272
rect 215478 237260 215484 237272
rect 215536 237260 215542 237312
rect 85574 237124 85580 237176
rect 85632 237164 85638 237176
rect 88978 237164 88984 237176
rect 85632 237136 88984 237164
rect 85632 237124 85638 237136
rect 88978 237124 88984 237136
rect 89036 237124 89042 237176
rect 106918 237056 106924 237108
rect 106976 237096 106982 237108
rect 113266 237096 113272 237108
rect 106976 237068 113272 237096
rect 106976 237056 106982 237068
rect 113266 237056 113272 237068
rect 113324 237056 113330 237108
rect 228358 236988 228364 237040
rect 228416 237028 228422 237040
rect 230474 237028 230480 237040
rect 228416 237000 230480 237028
rect 228416 236988 228422 237000
rect 230474 236988 230480 237000
rect 230532 236988 230538 237040
rect 72970 236648 72976 236700
rect 73028 236688 73034 236700
rect 79318 236688 79324 236700
rect 73028 236660 79324 236688
rect 73028 236648 73034 236660
rect 79318 236648 79324 236660
rect 79376 236648 79382 236700
rect 122190 236648 122196 236700
rect 122248 236688 122254 236700
rect 124214 236688 124220 236700
rect 122248 236660 124220 236688
rect 122248 236648 122254 236660
rect 124214 236648 124220 236660
rect 124272 236648 124278 236700
rect 125502 236648 125508 236700
rect 125560 236688 125566 236700
rect 171962 236688 171968 236700
rect 125560 236660 171968 236688
rect 125560 236648 125566 236660
rect 171962 236648 171968 236660
rect 172020 236648 172026 236700
rect 215478 236580 215484 236632
rect 215536 236620 215542 236632
rect 216306 236620 216312 236632
rect 215536 236592 216312 236620
rect 215536 236580 215542 236592
rect 216306 236580 216312 236592
rect 216364 236580 216370 236632
rect 217962 236580 217968 236632
rect 218020 236620 218026 236632
rect 220906 236620 220912 236632
rect 218020 236592 220912 236620
rect 218020 236580 218026 236592
rect 220906 236580 220912 236592
rect 220964 236620 220970 236632
rect 222102 236620 222108 236632
rect 220964 236592 222108 236620
rect 220964 236580 220970 236592
rect 222102 236580 222108 236592
rect 222160 236580 222166 236632
rect 107654 236444 107660 236496
rect 107712 236484 107718 236496
rect 108390 236484 108396 236496
rect 107712 236456 108396 236484
rect 107712 236444 107718 236456
rect 108390 236444 108396 236456
rect 108448 236444 108454 236496
rect 76098 235968 76104 236020
rect 76156 236008 76162 236020
rect 76742 236008 76748 236020
rect 76156 235980 76748 236008
rect 76156 235968 76162 235980
rect 76742 235968 76748 235980
rect 76800 235968 76806 236020
rect 97902 235968 97908 236020
rect 97960 236008 97966 236020
rect 98178 236008 98184 236020
rect 97960 235980 98184 236008
rect 97960 235968 97966 235980
rect 98178 235968 98184 235980
rect 98236 235968 98242 236020
rect 249150 235968 249156 236020
rect 249208 236008 249214 236020
rect 252370 236008 252376 236020
rect 249208 235980 252376 236008
rect 249208 235968 249214 235980
rect 252370 235968 252376 235980
rect 252428 235968 252434 236020
rect 191282 235900 191288 235952
rect 191340 235940 191346 235952
rect 213914 235940 213920 235952
rect 191340 235912 213920 235940
rect 191340 235900 191346 235912
rect 213914 235900 213920 235912
rect 213972 235900 213978 235952
rect 288434 235940 288440 235952
rect 258046 235912 288440 235940
rect 249886 235832 249892 235884
rect 249944 235872 249950 235884
rect 250530 235872 250536 235884
rect 249944 235844 250536 235872
rect 249944 235832 249950 235844
rect 250530 235832 250536 235844
rect 250588 235872 250594 235884
rect 258046 235872 258074 235912
rect 288434 235900 288440 235912
rect 288492 235900 288498 235952
rect 250588 235844 258074 235872
rect 250588 235832 250594 235844
rect 82906 235288 82912 235340
rect 82964 235328 82970 235340
rect 112990 235328 112996 235340
rect 82964 235300 112996 235328
rect 82964 235288 82970 235300
rect 112990 235288 112996 235300
rect 113048 235328 113054 235340
rect 116670 235328 116676 235340
rect 113048 235300 116676 235328
rect 113048 235288 113054 235300
rect 116670 235288 116676 235300
rect 116728 235288 116734 235340
rect 64506 235220 64512 235272
rect 64564 235260 64570 235272
rect 156782 235260 156788 235272
rect 64564 235232 156788 235260
rect 64564 235220 64570 235232
rect 156782 235220 156788 235232
rect 156840 235220 156846 235272
rect 164970 235220 164976 235272
rect 165028 235260 165034 235272
rect 197170 235260 197176 235272
rect 165028 235232 197176 235260
rect 165028 235220 165034 235232
rect 197170 235220 197176 235232
rect 197228 235220 197234 235272
rect 243630 235220 243636 235272
rect 243688 235260 243694 235272
rect 269206 235260 269212 235272
rect 243688 235232 269212 235260
rect 243688 235220 243694 235232
rect 269206 235220 269212 235232
rect 269264 235220 269270 235272
rect 213914 234608 213920 234660
rect 213972 234648 213978 234660
rect 214650 234648 214656 234660
rect 213972 234620 214656 234648
rect 213972 234608 213978 234620
rect 214650 234608 214656 234620
rect 214708 234608 214714 234660
rect 283558 234608 283564 234660
rect 283616 234648 283622 234660
rect 580258 234648 580264 234660
rect 283616 234620 580264 234648
rect 283616 234608 283622 234620
rect 580258 234608 580264 234620
rect 580316 234608 580322 234660
rect 166810 234540 166816 234592
rect 166868 234580 166874 234592
rect 256786 234580 256792 234592
rect 166868 234552 256792 234580
rect 166868 234540 166874 234552
rect 256786 234540 256792 234552
rect 256844 234540 256850 234592
rect 166350 234132 166356 234184
rect 166408 234172 166414 234184
rect 166810 234172 166816 234184
rect 166408 234144 166816 234172
rect 166408 234132 166414 234144
rect 166810 234132 166816 234144
rect 166868 234132 166874 234184
rect 94682 233928 94688 233980
rect 94740 233968 94746 233980
rect 95326 233968 95332 233980
rect 94740 233940 95332 233968
rect 94740 233928 94746 233940
rect 95326 233928 95332 233940
rect 95384 233928 95390 233980
rect 61838 233860 61844 233912
rect 61896 233900 61902 233912
rect 76558 233900 76564 233912
rect 61896 233872 76564 233900
rect 61896 233860 61902 233872
rect 76558 233860 76564 233872
rect 76616 233860 76622 233912
rect 77386 233860 77392 233912
rect 77444 233900 77450 233912
rect 87690 233900 87696 233912
rect 77444 233872 87696 233900
rect 77444 233860 77450 233872
rect 87690 233860 87696 233872
rect 87748 233860 87754 233912
rect 91002 233860 91008 233912
rect 91060 233900 91066 233912
rect 125410 233900 125416 233912
rect 91060 233872 125416 233900
rect 91060 233860 91066 233872
rect 125410 233860 125416 233872
rect 125468 233900 125474 233912
rect 128354 233900 128360 233912
rect 125468 233872 128360 233900
rect 125468 233860 125474 233872
rect 128354 233860 128360 233872
rect 128412 233860 128418 233912
rect 184290 233860 184296 233912
rect 184348 233900 184354 233912
rect 215938 233900 215944 233912
rect 184348 233872 215944 233900
rect 184348 233860 184354 233872
rect 215938 233860 215944 233872
rect 215996 233860 216002 233912
rect 257982 233860 257988 233912
rect 258040 233900 258046 233912
rect 265158 233900 265164 233912
rect 258040 233872 265164 233900
rect 258040 233860 258046 233872
rect 265158 233860 265164 233872
rect 265216 233860 265222 233912
rect 269758 233656 269764 233708
rect 269816 233696 269822 233708
rect 274818 233696 274824 233708
rect 269816 233668 274824 233696
rect 269816 233656 269822 233668
rect 274818 233656 274824 233668
rect 274876 233656 274882 233708
rect 108298 233180 108304 233232
rect 108356 233220 108362 233232
rect 108942 233220 108948 233232
rect 108356 233192 108948 233220
rect 108356 233180 108362 233192
rect 108942 233180 108948 233192
rect 109000 233220 109006 233232
rect 109000 233192 258074 233220
rect 109000 233180 109006 233192
rect 258046 233152 258074 233192
rect 278038 233180 278044 233232
rect 278096 233220 278102 233232
rect 278866 233220 278872 233232
rect 278096 233192 278872 233220
rect 278096 233180 278102 233192
rect 278866 233180 278872 233192
rect 278924 233180 278930 233232
rect 279050 233152 279056 233164
rect 258046 233124 279056 233152
rect 279050 233112 279056 233124
rect 279108 233112 279114 233164
rect 73154 232500 73160 232552
rect 73212 232540 73218 232552
rect 77294 232540 77300 232552
rect 73212 232512 77300 232540
rect 73212 232500 73218 232512
rect 77294 232500 77300 232512
rect 77352 232500 77358 232552
rect 78674 232500 78680 232552
rect 78732 232540 78738 232552
rect 91002 232540 91008 232552
rect 78732 232512 91008 232540
rect 78732 232500 78738 232512
rect 91002 232500 91008 232512
rect 91060 232540 91066 232552
rect 102134 232540 102140 232552
rect 91060 232512 102140 232540
rect 91060 232500 91066 232512
rect 102134 232500 102140 232512
rect 102192 232500 102198 232552
rect 166442 232500 166448 232552
rect 166500 232540 166506 232552
rect 196618 232540 196624 232552
rect 166500 232512 196624 232540
rect 166500 232500 166506 232512
rect 196618 232500 196624 232512
rect 196676 232500 196682 232552
rect 204898 232500 204904 232552
rect 204956 232540 204962 232552
rect 252738 232540 252744 232552
rect 204956 232512 252744 232540
rect 204956 232500 204962 232512
rect 252738 232500 252744 232512
rect 252796 232500 252802 232552
rect 258718 232500 258724 232552
rect 258776 232540 258782 232552
rect 270678 232540 270684 232552
rect 258776 232512 270684 232540
rect 258776 232500 258782 232512
rect 270678 232500 270684 232512
rect 270736 232500 270742 232552
rect 7650 231820 7656 231872
rect 7708 231860 7714 231872
rect 96614 231860 96620 231872
rect 7708 231832 96620 231860
rect 7708 231820 7714 231832
rect 96614 231820 96620 231832
rect 96672 231860 96678 231872
rect 97258 231860 97264 231872
rect 96672 231832 97264 231860
rect 96672 231820 96678 231832
rect 97258 231820 97264 231832
rect 97316 231820 97322 231872
rect 278866 231820 278872 231872
rect 278924 231860 278930 231872
rect 580166 231860 580172 231872
rect 278924 231832 580172 231860
rect 278924 231820 278930 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 89070 231752 89076 231804
rect 89128 231792 89134 231804
rect 170490 231792 170496 231804
rect 89128 231764 170496 231792
rect 89128 231752 89134 231764
rect 170490 231752 170496 231764
rect 170548 231752 170554 231804
rect 215938 231752 215944 231804
rect 215996 231792 216002 231804
rect 266446 231792 266452 231804
rect 215996 231764 266452 231792
rect 215996 231752 216002 231764
rect 266446 231752 266452 231764
rect 266504 231752 266510 231804
rect 67450 231684 67456 231736
rect 67508 231724 67514 231736
rect 112530 231724 112536 231736
rect 67508 231696 112536 231724
rect 67508 231684 67514 231696
rect 112530 231684 112536 231696
rect 112588 231684 112594 231736
rect 63218 231072 63224 231124
rect 63276 231112 63282 231124
rect 73430 231112 73436 231124
rect 63276 231084 73436 231112
rect 63276 231072 63282 231084
rect 73430 231072 73436 231084
rect 73488 231072 73494 231124
rect 138842 231072 138848 231124
rect 138900 231112 138906 231124
rect 213822 231112 213828 231124
rect 138900 231084 213828 231112
rect 138900 231072 138906 231084
rect 213822 231072 213828 231084
rect 213880 231072 213886 231124
rect 224310 231072 224316 231124
rect 224368 231112 224374 231124
rect 280798 231112 280804 231124
rect 224368 231084 280804 231112
rect 224368 231072 224374 231084
rect 280798 231072 280804 231084
rect 280856 231072 280862 231124
rect 80330 230392 80336 230444
rect 80388 230432 80394 230444
rect 156598 230432 156604 230444
rect 80388 230404 156604 230432
rect 80388 230392 80394 230404
rect 156598 230392 156604 230404
rect 156656 230432 156662 230444
rect 164970 230432 164976 230444
rect 156656 230404 164976 230432
rect 156656 230392 156662 230404
rect 164970 230392 164976 230404
rect 165028 230392 165034 230444
rect 185670 230392 185676 230444
rect 185728 230432 185734 230444
rect 262214 230432 262220 230444
rect 185728 230404 262220 230432
rect 185728 230392 185734 230404
rect 262214 230392 262220 230404
rect 262272 230392 262278 230444
rect 77570 229712 77576 229764
rect 77628 229752 77634 229764
rect 105630 229752 105636 229764
rect 77628 229724 105636 229752
rect 77628 229712 77634 229724
rect 105630 229712 105636 229724
rect 105688 229712 105694 229764
rect 120718 229712 120724 229764
rect 120776 229752 120782 229764
rect 160922 229752 160928 229764
rect 120776 229724 160928 229752
rect 120776 229712 120782 229724
rect 160922 229712 160928 229724
rect 160980 229712 160986 229764
rect 161014 229712 161020 229764
rect 161072 229752 161078 229764
rect 204438 229752 204444 229764
rect 161072 229724 204444 229752
rect 161072 229712 161078 229724
rect 204438 229712 204444 229724
rect 204496 229712 204502 229764
rect 235902 229712 235908 229764
rect 235960 229752 235966 229764
rect 255590 229752 255596 229764
rect 235960 229724 255596 229752
rect 235960 229712 235966 229724
rect 255590 229712 255596 229724
rect 255648 229712 255654 229764
rect 89714 229032 89720 229084
rect 89772 229072 89778 229084
rect 105538 229072 105544 229084
rect 89772 229044 105544 229072
rect 89772 229032 89778 229044
rect 105538 229032 105544 229044
rect 105596 229032 105602 229084
rect 156782 229032 156788 229084
rect 156840 229072 156846 229084
rect 273346 229072 273352 229084
rect 156840 229044 273352 229072
rect 156840 229032 156846 229044
rect 273346 229032 273352 229044
rect 273404 229032 273410 229084
rect 65886 228352 65892 228404
rect 65944 228392 65950 228404
rect 76098 228392 76104 228404
rect 65944 228364 76104 228392
rect 65944 228352 65950 228364
rect 76098 228352 76104 228364
rect 76156 228392 76162 228404
rect 77202 228392 77208 228404
rect 76156 228364 77208 228392
rect 76156 228352 76162 228364
rect 77202 228352 77208 228364
rect 77260 228352 77266 228404
rect 156782 227808 156788 227860
rect 156840 227848 156846 227860
rect 157242 227848 157248 227860
rect 156840 227820 157248 227848
rect 156840 227808 156846 227820
rect 157242 227808 157248 227820
rect 157300 227808 157306 227860
rect 77202 227740 77208 227792
rect 77260 227780 77266 227792
rect 187694 227780 187700 227792
rect 77260 227752 187700 227780
rect 77260 227740 77266 227752
rect 187694 227740 187700 227752
rect 187752 227780 187758 227792
rect 188338 227780 188344 227792
rect 187752 227752 188344 227780
rect 187752 227740 187758 227752
rect 188338 227740 188344 227752
rect 188396 227740 188402 227792
rect 155402 227672 155408 227724
rect 155460 227712 155466 227724
rect 277394 227712 277400 227724
rect 155460 227684 277400 227712
rect 155460 227672 155466 227684
rect 277394 227672 277400 227684
rect 277452 227672 277458 227724
rect 105538 227060 105544 227112
rect 105596 227100 105602 227112
rect 118694 227100 118700 227112
rect 105596 227072 118700 227100
rect 105596 227060 105602 227072
rect 118694 227060 118700 227072
rect 118752 227060 118758 227112
rect 84010 226992 84016 227044
rect 84068 227032 84074 227044
rect 84194 227032 84200 227044
rect 84068 227004 84200 227032
rect 84068 226992 84074 227004
rect 84194 226992 84200 227004
rect 84252 226992 84258 227044
rect 87046 226992 87052 227044
rect 87104 227032 87110 227044
rect 104158 227032 104164 227044
rect 87104 227004 104164 227032
rect 87104 226992 87110 227004
rect 104158 226992 104164 227004
rect 104216 227032 104222 227044
rect 110506 227032 110512 227044
rect 104216 227004 110512 227032
rect 104216 226992 104222 227004
rect 110506 226992 110512 227004
rect 110564 226992 110570 227044
rect 195330 226992 195336 227044
rect 195388 227032 195394 227044
rect 224218 227032 224224 227044
rect 195388 227004 224224 227032
rect 195388 226992 195394 227004
rect 224218 226992 224224 227004
rect 224276 227032 224282 227044
rect 254578 227032 254584 227044
rect 224276 227004 254584 227032
rect 224276 226992 224282 227004
rect 254578 226992 254584 227004
rect 254636 226992 254642 227044
rect 95142 226312 95148 226364
rect 95200 226352 95206 226364
rect 100846 226352 100852 226364
rect 95200 226324 100852 226352
rect 95200 226312 95206 226324
rect 100846 226312 100852 226324
rect 100904 226312 100910 226364
rect 80054 226244 80060 226296
rect 80112 226284 80118 226296
rect 113174 226284 113180 226296
rect 80112 226256 113180 226284
rect 80112 226244 80118 226256
rect 113174 226244 113180 226256
rect 113232 226284 113238 226296
rect 113910 226284 113916 226296
rect 113232 226256 113916 226284
rect 113232 226244 113238 226256
rect 113910 226244 113916 226256
rect 113968 226244 113974 226296
rect 245562 225632 245568 225684
rect 245620 225672 245626 225684
rect 257338 225672 257344 225684
rect 245620 225644 257344 225672
rect 245620 225632 245626 225644
rect 257338 225632 257344 225644
rect 257396 225632 257402 225684
rect 242802 225564 242808 225616
rect 242860 225604 242866 225616
rect 289998 225604 290004 225616
rect 242860 225576 290004 225604
rect 242860 225564 242866 225576
rect 289998 225564 290004 225576
rect 290056 225564 290062 225616
rect 100018 224952 100024 225004
rect 100076 224992 100082 225004
rect 242250 224992 242256 225004
rect 100076 224964 242256 224992
rect 100076 224952 100082 224964
rect 242250 224952 242256 224964
rect 242308 224992 242314 225004
rect 242802 224992 242808 225004
rect 242308 224964 242808 224992
rect 242308 224952 242314 224964
rect 242802 224952 242808 224964
rect 242860 224952 242866 225004
rect 176010 224884 176016 224936
rect 176068 224924 176074 224936
rect 259730 224924 259736 224936
rect 176068 224896 259736 224924
rect 176068 224884 176074 224896
rect 259730 224884 259736 224896
rect 259788 224884 259794 224936
rect 76742 224204 76748 224256
rect 76800 224244 76806 224256
rect 108298 224244 108304 224256
rect 76800 224216 108304 224244
rect 76800 224204 76806 224216
rect 108298 224204 108304 224216
rect 108356 224204 108362 224256
rect 121362 224204 121368 224256
rect 121420 224244 121426 224256
rect 187050 224244 187056 224256
rect 121420 224216 187056 224244
rect 121420 224204 121426 224216
rect 187050 224204 187056 224216
rect 187108 224204 187114 224256
rect 234540 223604 235672 223632
rect 196618 223524 196624 223576
rect 196676 223564 196682 223576
rect 234540 223564 234568 223604
rect 196676 223536 234568 223564
rect 196676 223524 196682 223536
rect 234614 223524 234620 223576
rect 234672 223564 234678 223576
rect 235534 223564 235540 223576
rect 234672 223536 235540 223564
rect 234672 223524 234678 223536
rect 235534 223524 235540 223536
rect 235592 223524 235598 223576
rect 235644 223564 235672 223604
rect 237466 223564 237472 223576
rect 235644 223536 237472 223564
rect 237466 223524 237472 223536
rect 237524 223564 237530 223576
rect 237926 223564 237932 223576
rect 237524 223536 237932 223564
rect 237524 223524 237530 223536
rect 237926 223524 237932 223536
rect 237984 223524 237990 223576
rect 204438 223456 204444 223508
rect 204496 223496 204502 223508
rect 234632 223496 234660 223524
rect 204496 223468 234660 223496
rect 204496 223456 204502 223468
rect 80698 222844 80704 222896
rect 80756 222884 80762 222896
rect 104986 222884 104992 222896
rect 80756 222856 104992 222884
rect 80756 222844 80762 222856
rect 104986 222844 104992 222856
rect 105044 222844 105050 222896
rect 111702 222844 111708 222896
rect 111760 222884 111766 222896
rect 188430 222884 188436 222896
rect 111760 222856 188436 222884
rect 111760 222844 111766 222856
rect 188430 222844 188436 222856
rect 188488 222844 188494 222896
rect 255314 222844 255320 222896
rect 255372 222884 255378 222896
rect 287330 222884 287336 222896
rect 255372 222856 287336 222884
rect 255372 222844 255378 222856
rect 287330 222844 287336 222856
rect 287388 222884 287394 222896
rect 580350 222884 580356 222896
rect 287388 222856 580356 222884
rect 287388 222844 287394 222856
rect 580350 222844 580356 222856
rect 580408 222844 580414 222896
rect 153838 222096 153844 222148
rect 153896 222136 153902 222148
rect 252830 222136 252836 222148
rect 153896 222108 252836 222136
rect 153896 222096 153902 222108
rect 252830 222096 252836 222108
rect 252888 222096 252894 222148
rect 133230 221484 133236 221536
rect 133288 221524 133294 221536
rect 148410 221524 148416 221536
rect 133288 221496 148416 221524
rect 133288 221484 133294 221496
rect 148410 221484 148416 221496
rect 148468 221484 148474 221536
rect 82814 221416 82820 221468
rect 82872 221456 82878 221468
rect 204990 221456 204996 221468
rect 82872 221428 204996 221456
rect 82872 221416 82878 221428
rect 204990 221416 204996 221428
rect 205048 221416 205054 221468
rect 227806 221416 227812 221468
rect 227864 221456 227870 221468
rect 255314 221456 255320 221468
rect 227864 221428 255320 221456
rect 227864 221416 227870 221428
rect 255314 221416 255320 221428
rect 255372 221416 255378 221468
rect 88334 220736 88340 220788
rect 88392 220776 88398 220788
rect 121454 220776 121460 220788
rect 88392 220748 121460 220776
rect 88392 220736 88398 220748
rect 121454 220736 121460 220748
rect 121512 220776 121518 220788
rect 122190 220776 122196 220788
rect 121512 220748 122196 220776
rect 121512 220736 121518 220748
rect 122190 220736 122196 220748
rect 122248 220736 122254 220788
rect 163682 220736 163688 220788
rect 163740 220776 163746 220788
rect 164142 220776 164148 220788
rect 163740 220748 164148 220776
rect 163740 220736 163746 220748
rect 164142 220736 164148 220748
rect 164200 220776 164206 220788
rect 227070 220776 227076 220788
rect 164200 220748 227076 220776
rect 164200 220736 164206 220748
rect 227070 220736 227076 220748
rect 227128 220736 227134 220788
rect 118602 220056 118608 220108
rect 118660 220096 118666 220108
rect 182910 220096 182916 220108
rect 118660 220068 182916 220096
rect 118660 220056 118666 220068
rect 182910 220056 182916 220068
rect 182968 220056 182974 220108
rect 226978 220056 226984 220108
rect 227036 220096 227042 220108
rect 251910 220096 251916 220108
rect 227036 220068 251916 220096
rect 227036 220056 227042 220068
rect 251910 220056 251916 220068
rect 251968 220056 251974 220108
rect 232590 218764 232596 218816
rect 232648 218804 232654 218816
rect 283558 218804 283564 218816
rect 232648 218776 283564 218804
rect 232648 218764 232654 218776
rect 283558 218764 283564 218776
rect 283616 218764 283622 218816
rect 147122 218696 147128 218748
rect 147180 218736 147186 218748
rect 235994 218736 236000 218748
rect 147180 218708 236000 218736
rect 147180 218696 147186 218708
rect 235994 218696 236000 218708
rect 236052 218696 236058 218748
rect 101490 217948 101496 218000
rect 101548 217988 101554 218000
rect 103514 217988 103520 218000
rect 101548 217960 103520 217988
rect 101548 217948 101554 217960
rect 103514 217948 103520 217960
rect 103572 217988 103578 218000
rect 284478 217988 284484 218000
rect 103572 217960 284484 217988
rect 103572 217948 103578 217960
rect 284478 217948 284484 217960
rect 284536 217948 284542 218000
rect 104342 217880 104348 217932
rect 104400 217920 104406 217932
rect 245562 217920 245568 217932
rect 104400 217892 245568 217920
rect 104400 217880 104406 217892
rect 245562 217880 245568 217892
rect 245620 217880 245626 217932
rect 256602 217268 256608 217320
rect 256660 217308 256666 217320
rect 273438 217308 273444 217320
rect 256660 217280 273444 217308
rect 256660 217268 256666 217280
rect 273438 217268 273444 217280
rect 273496 217268 273502 217320
rect 245562 216656 245568 216708
rect 245620 216696 245626 216708
rect 246298 216696 246304 216708
rect 245620 216668 246304 216696
rect 245620 216656 245626 216668
rect 246298 216656 246304 216668
rect 246356 216656 246362 216708
rect 160922 216588 160928 216640
rect 160980 216628 160986 216640
rect 161382 216628 161388 216640
rect 160980 216600 161388 216628
rect 160980 216588 160986 216600
rect 161382 216588 161388 216600
rect 161440 216628 161446 216640
rect 278866 216628 278872 216640
rect 161440 216600 278872 216628
rect 161440 216588 161446 216600
rect 278866 216588 278872 216600
rect 278924 216588 278930 216640
rect 49602 215908 49608 215960
rect 49660 215948 49666 215960
rect 162118 215948 162124 215960
rect 49660 215920 162124 215948
rect 49660 215908 49666 215920
rect 162118 215908 162124 215920
rect 162176 215908 162182 215960
rect 3418 214956 3424 215008
rect 3476 214996 3482 215008
rect 7558 214996 7564 215008
rect 3476 214968 7564 214996
rect 3476 214956 3482 214968
rect 7558 214956 7564 214968
rect 7616 214996 7622 215008
rect 8202 214996 8208 215008
rect 7616 214968 8208 214996
rect 7616 214956 7622 214968
rect 8202 214956 8208 214968
rect 8260 214956 8266 215008
rect 86954 214548 86960 214600
rect 87012 214588 87018 214600
rect 111794 214588 111800 214600
rect 87012 214560 111800 214588
rect 87012 214548 87018 214560
rect 111794 214548 111800 214560
rect 111852 214548 111858 214600
rect 218698 214548 218704 214600
rect 218756 214588 218762 214600
rect 237650 214588 237656 214600
rect 218756 214560 237656 214588
rect 218756 214548 218762 214560
rect 237650 214548 237656 214560
rect 237708 214548 237714 214600
rect 111794 213936 111800 213988
rect 111852 213976 111858 213988
rect 196618 213976 196624 213988
rect 111852 213948 196624 213976
rect 111852 213936 111858 213948
rect 196618 213936 196624 213948
rect 196676 213936 196682 213988
rect 100110 213188 100116 213240
rect 100168 213228 100174 213240
rect 266354 213228 266360 213240
rect 100168 213200 266360 213228
rect 100168 213188 100174 213200
rect 266354 213188 266360 213200
rect 266412 213188 266418 213240
rect 181530 212440 181536 212492
rect 181588 212480 181594 212492
rect 182082 212480 182088 212492
rect 181588 212452 182088 212480
rect 181588 212440 181594 212452
rect 182082 212440 182088 212452
rect 182140 212480 182146 212492
rect 249150 212480 249156 212492
rect 182140 212452 249156 212480
rect 182140 212440 182146 212452
rect 249150 212440 249156 212452
rect 249208 212440 249214 212492
rect 236638 212236 236644 212288
rect 236696 212276 236702 212288
rect 237466 212276 237472 212288
rect 236696 212248 237472 212276
rect 236696 212236 236702 212248
rect 237466 212236 237472 212248
rect 237524 212236 237530 212288
rect 58894 211760 58900 211812
rect 58952 211800 58958 211812
rect 159542 211800 159548 211812
rect 58952 211772 159548 211800
rect 58952 211760 58958 211772
rect 159542 211760 159548 211772
rect 159600 211760 159606 211812
rect 259362 211760 259368 211812
rect 259420 211800 259426 211812
rect 582650 211800 582656 211812
rect 259420 211772 582656 211800
rect 259420 211760 259426 211772
rect 582650 211760 582656 211772
rect 582708 211760 582714 211812
rect 253842 211148 253848 211200
rect 253900 211188 253906 211200
rect 258166 211188 258172 211200
rect 253900 211160 258172 211188
rect 253900 211148 253906 211160
rect 258166 211148 258172 211160
rect 258224 211188 258230 211200
rect 259362 211188 259368 211200
rect 258224 211160 259368 211188
rect 258224 211148 258230 211160
rect 259362 211148 259368 211160
rect 259420 211148 259426 211200
rect 56502 211080 56508 211132
rect 56560 211120 56566 211132
rect 167730 211120 167736 211132
rect 56560 211092 167736 211120
rect 56560 211080 56566 211092
rect 167730 211080 167736 211092
rect 167788 211120 167794 211132
rect 287054 211120 287060 211132
rect 167788 211092 287060 211120
rect 167788 211080 167794 211092
rect 287054 211080 287060 211092
rect 287112 211080 287118 211132
rect 161290 209720 161296 209772
rect 161348 209760 161354 209772
rect 232590 209760 232596 209772
rect 161348 209732 232596 209760
rect 161348 209720 161354 209732
rect 232590 209720 232596 209732
rect 232648 209720 232654 209772
rect 160830 209516 160836 209568
rect 160888 209556 160894 209568
rect 161290 209556 161296 209568
rect 160888 209528 161296 209556
rect 160888 209516 160894 209528
rect 161290 209516 161296 209528
rect 161348 209516 161354 209568
rect 97258 209040 97264 209092
rect 97316 209080 97322 209092
rect 129734 209080 129740 209092
rect 97316 209052 129740 209080
rect 97316 209040 97322 209052
rect 129734 209040 129740 209052
rect 129792 209040 129798 209092
rect 129734 208360 129740 208412
rect 129792 208400 129798 208412
rect 273346 208400 273352 208412
rect 129792 208372 273352 208400
rect 129792 208360 129798 208372
rect 273346 208360 273352 208372
rect 273404 208360 273410 208412
rect 102226 208292 102232 208344
rect 102284 208332 102290 208344
rect 262306 208332 262312 208344
rect 102284 208304 262312 208332
rect 102284 208292 102290 208304
rect 262306 208292 262312 208304
rect 262364 208292 262370 208344
rect 93118 207068 93124 207120
rect 93176 207108 93182 207120
rect 96062 207108 96068 207120
rect 93176 207080 96068 207108
rect 93176 207068 93182 207080
rect 96062 207068 96068 207080
rect 96120 207108 96126 207120
rect 96120 207080 103514 207108
rect 96120 207068 96126 207080
rect 98638 207000 98644 207052
rect 98696 207040 98702 207052
rect 102226 207040 102232 207052
rect 98696 207012 102232 207040
rect 98696 207000 98702 207012
rect 102226 207000 102232 207012
rect 102284 207000 102290 207052
rect 103486 207040 103514 207080
rect 263686 207040 263692 207052
rect 103486 207012 263692 207040
rect 263686 207000 263692 207012
rect 263744 207000 263750 207052
rect 196618 206932 196624 206984
rect 196676 206972 196682 206984
rect 197262 206972 197268 206984
rect 196676 206944 197268 206972
rect 196676 206932 196682 206944
rect 197262 206932 197268 206944
rect 197320 206972 197326 206984
rect 269298 206972 269304 206984
rect 197320 206944 269304 206972
rect 197320 206932 197326 206944
rect 269298 206932 269304 206944
rect 269356 206932 269362 206984
rect 95234 206252 95240 206304
rect 95292 206292 95298 206304
rect 122834 206292 122840 206304
rect 95292 206264 122840 206292
rect 95292 206252 95298 206264
rect 122834 206252 122840 206264
rect 122892 206292 122898 206304
rect 123754 206292 123760 206304
rect 122892 206264 123760 206292
rect 122892 206252 122898 206264
rect 123754 206252 123760 206264
rect 123812 206252 123818 206304
rect 123754 205640 123760 205692
rect 123812 205680 123818 205692
rect 280154 205680 280160 205692
rect 123812 205652 280160 205680
rect 123812 205640 123818 205652
rect 280154 205640 280160 205652
rect 280212 205680 280218 205692
rect 280430 205680 280436 205692
rect 280212 205652 280436 205680
rect 280212 205640 280218 205652
rect 280430 205640 280436 205652
rect 280488 205640 280494 205692
rect 93854 204960 93860 205012
rect 93912 205000 93918 205012
rect 103514 205000 103520 205012
rect 93912 204972 103520 205000
rect 93912 204960 93918 204972
rect 103514 204960 103520 204972
rect 103572 205000 103578 205012
rect 104710 205000 104716 205012
rect 103572 204972 104716 205000
rect 103572 204960 103578 204972
rect 104710 204960 104716 204972
rect 104768 204960 104774 205012
rect 84010 204892 84016 204944
rect 84068 204932 84074 204944
rect 115198 204932 115204 204944
rect 84068 204904 115204 204932
rect 84068 204892 84074 204904
rect 115198 204892 115204 204904
rect 115256 204892 115262 204944
rect 225782 204892 225788 204944
rect 225840 204932 225846 204944
rect 266538 204932 266544 204944
rect 225840 204904 266544 204932
rect 225840 204892 225846 204904
rect 266538 204892 266544 204904
rect 266596 204892 266602 204944
rect 104710 204348 104716 204400
rect 104768 204388 104774 204400
rect 225138 204388 225144 204400
rect 104768 204360 225144 204388
rect 104768 204348 104774 204360
rect 225138 204348 225144 204360
rect 225196 204388 225202 204400
rect 225782 204388 225788 204400
rect 225196 204360 225788 204388
rect 225196 204348 225202 204360
rect 225782 204348 225788 204360
rect 225840 204348 225846 204400
rect 114646 204280 114652 204332
rect 114704 204320 114710 204332
rect 115198 204320 115204 204332
rect 114704 204292 115204 204320
rect 114704 204280 114710 204292
rect 115198 204280 115204 204292
rect 115256 204320 115262 204332
rect 258074 204320 258080 204332
rect 115256 204292 258080 204320
rect 115256 204280 115262 204292
rect 258074 204280 258080 204292
rect 258132 204280 258138 204332
rect 266998 203600 267004 203652
rect 267056 203640 267062 203652
rect 284478 203640 284484 203652
rect 267056 203612 284484 203640
rect 267056 203600 267062 203612
rect 284478 203600 284484 203612
rect 284536 203600 284542 203652
rect 200022 203532 200028 203584
rect 200080 203572 200086 203584
rect 582466 203572 582472 203584
rect 200080 203544 582472 203572
rect 200080 203532 200086 203544
rect 582466 203532 582472 203544
rect 582524 203532 582530 203584
rect 99466 202784 99472 202836
rect 99524 202824 99530 202836
rect 100110 202824 100116 202836
rect 99524 202796 100116 202824
rect 99524 202784 99530 202796
rect 100110 202784 100116 202796
rect 100168 202784 100174 202836
rect 111242 202784 111248 202836
rect 111300 202824 111306 202836
rect 201586 202824 201592 202836
rect 111300 202796 201592 202824
rect 111300 202784 111306 202796
rect 201586 202784 201592 202796
rect 201644 202824 201650 202836
rect 202230 202824 202236 202836
rect 201644 202796 202236 202824
rect 201644 202784 201650 202796
rect 202230 202784 202236 202796
rect 202288 202784 202294 202836
rect 201402 202716 201408 202768
rect 201460 202756 201466 202768
rect 224310 202756 224316 202768
rect 201460 202728 224316 202756
rect 201460 202716 201466 202728
rect 224310 202716 224316 202728
rect 224368 202716 224374 202768
rect 3234 202104 3240 202156
rect 3292 202144 3298 202156
rect 99466 202144 99472 202156
rect 3292 202116 99472 202144
rect 3292 202104 3298 202116
rect 99466 202104 99472 202116
rect 99524 202104 99530 202156
rect 214650 202104 214656 202156
rect 214708 202144 214714 202156
rect 222286 202144 222292 202156
rect 214708 202116 222292 202144
rect 214708 202104 214714 202116
rect 222286 202104 222292 202116
rect 222344 202104 222350 202156
rect 243538 202104 243544 202156
rect 243596 202144 243602 202156
rect 280338 202144 280344 202156
rect 243596 202116 280344 202144
rect 243596 202104 243602 202116
rect 280338 202104 280344 202116
rect 280396 202104 280402 202156
rect 148410 201492 148416 201544
rect 148468 201532 148474 201544
rect 152642 201532 152648 201544
rect 148468 201504 152648 201532
rect 148468 201492 148474 201504
rect 152642 201492 152648 201504
rect 152700 201492 152706 201544
rect 54846 201424 54852 201476
rect 54904 201464 54910 201476
rect 55030 201464 55036 201476
rect 54904 201436 55036 201464
rect 54904 201424 54910 201436
rect 55030 201424 55036 201436
rect 55088 201464 55094 201476
rect 247678 201464 247684 201476
rect 55088 201436 247684 201464
rect 55088 201424 55094 201436
rect 247678 201424 247684 201436
rect 247736 201424 247742 201476
rect 96522 200744 96528 200796
rect 96580 200784 96586 200796
rect 109678 200784 109684 200796
rect 96580 200756 109684 200784
rect 96580 200744 96586 200756
rect 109678 200744 109684 200756
rect 109736 200744 109742 200796
rect 244918 200744 244924 200796
rect 244976 200784 244982 200796
rect 277578 200784 277584 200796
rect 244976 200756 277584 200784
rect 244976 200744 244982 200756
rect 277578 200744 277584 200756
rect 277636 200744 277642 200796
rect 74534 199452 74540 199504
rect 74592 199492 74598 199504
rect 95878 199492 95884 199504
rect 74592 199464 95884 199492
rect 74592 199452 74598 199464
rect 95878 199452 95884 199464
rect 95936 199452 95942 199504
rect 52270 199384 52276 199436
rect 52328 199424 52334 199436
rect 79410 199424 79416 199436
rect 52328 199396 79416 199424
rect 52328 199384 52334 199396
rect 79410 199384 79416 199396
rect 79468 199384 79474 199436
rect 117222 199384 117228 199436
rect 117280 199424 117286 199436
rect 126330 199424 126336 199436
rect 117280 199396 126336 199424
rect 117280 199384 117286 199396
rect 126330 199384 126336 199396
rect 126388 199384 126394 199436
rect 153838 199384 153844 199436
rect 153896 199424 153902 199436
rect 173342 199424 173348 199436
rect 153896 199396 173348 199424
rect 153896 199384 153902 199396
rect 173342 199384 173348 199396
rect 173400 199384 173406 199436
rect 193122 199384 193128 199436
rect 193180 199424 193186 199436
rect 226426 199424 226432 199436
rect 193180 199396 226432 199424
rect 193180 199384 193186 199396
rect 226426 199384 226432 199396
rect 226484 199384 226490 199436
rect 256050 199384 256056 199436
rect 256108 199424 256114 199436
rect 267918 199424 267924 199436
rect 256108 199396 267924 199424
rect 256108 199384 256114 199396
rect 267918 199384 267924 199396
rect 267976 199384 267982 199436
rect 162578 198636 162584 198688
rect 162636 198676 162642 198688
rect 291286 198676 291292 198688
rect 162636 198648 291292 198676
rect 162636 198636 162642 198648
rect 291286 198636 291292 198648
rect 291344 198636 291350 198688
rect 53466 198568 53472 198620
rect 53524 198608 53530 198620
rect 169754 198608 169760 198620
rect 53524 198580 169760 198608
rect 53524 198568 53530 198580
rect 169754 198568 169760 198580
rect 169812 198568 169818 198620
rect 162118 198228 162124 198280
rect 162176 198268 162182 198280
rect 162578 198268 162584 198280
rect 162176 198240 162584 198268
rect 162176 198228 162182 198240
rect 162578 198228 162584 198240
rect 162636 198228 162642 198280
rect 92382 197956 92388 198008
rect 92440 197996 92446 198008
rect 125594 197996 125600 198008
rect 92440 197968 125600 197996
rect 92440 197956 92446 197968
rect 125594 197956 125600 197968
rect 125652 197956 125658 198008
rect 176102 197956 176108 198008
rect 176160 197996 176166 198008
rect 196618 197996 196624 198008
rect 176160 197968 196624 197996
rect 176160 197956 176166 197968
rect 196618 197956 196624 197968
rect 196676 197956 196682 198008
rect 169754 197888 169760 197940
rect 169812 197928 169818 197940
rect 171042 197928 171048 197940
rect 169812 197900 171048 197928
rect 169812 197888 169818 197900
rect 171042 197888 171048 197900
rect 171100 197928 171106 197940
rect 171870 197928 171876 197940
rect 171100 197900 171876 197928
rect 171100 197888 171106 197900
rect 171870 197888 171876 197900
rect 171928 197888 171934 197940
rect 195238 196596 195244 196648
rect 195296 196636 195302 196648
rect 226334 196636 226340 196648
rect 195296 196608 226340 196636
rect 195296 196596 195302 196608
rect 226334 196596 226340 196608
rect 226392 196596 226398 196648
rect 49602 195236 49608 195288
rect 49660 195276 49666 195288
rect 130470 195276 130476 195288
rect 49660 195248 130476 195276
rect 49660 195236 49666 195248
rect 130470 195236 130476 195248
rect 130528 195236 130534 195288
rect 204990 195236 204996 195288
rect 205048 195276 205054 195288
rect 260834 195276 260840 195288
rect 205048 195248 260840 195276
rect 205048 195236 205054 195248
rect 260834 195236 260840 195248
rect 260892 195236 260898 195288
rect 87690 193808 87696 193860
rect 87748 193848 87754 193860
rect 102778 193848 102784 193860
rect 87748 193820 102784 193848
rect 87748 193808 87754 193820
rect 102778 193808 102784 193820
rect 102836 193808 102842 193860
rect 111150 193808 111156 193860
rect 111208 193848 111214 193860
rect 151262 193848 151268 193860
rect 111208 193820 151268 193848
rect 111208 193808 111214 193820
rect 151262 193808 151268 193820
rect 151320 193808 151326 193860
rect 195238 193808 195244 193860
rect 195296 193848 195302 193860
rect 287146 193848 287152 193860
rect 195296 193820 287152 193848
rect 195296 193808 195302 193820
rect 287146 193808 287152 193820
rect 287204 193808 287210 193860
rect 27522 192448 27528 192500
rect 27580 192488 27586 192500
rect 138750 192488 138756 192500
rect 27580 192460 138756 192488
rect 27580 192448 27586 192460
rect 138750 192448 138756 192460
rect 138808 192448 138814 192500
rect 195330 192448 195336 192500
rect 195388 192488 195394 192500
rect 243630 192488 243636 192500
rect 195388 192460 243636 192488
rect 195388 192448 195394 192460
rect 243630 192448 243636 192460
rect 243688 192448 243694 192500
rect 246298 192448 246304 192500
rect 246356 192488 246362 192500
rect 580166 192488 580172 192500
rect 246356 192460 580172 192488
rect 246356 192448 246362 192460
rect 580166 192448 580172 192460
rect 580224 192448 580230 192500
rect 184750 191088 184756 191140
rect 184808 191128 184814 191140
rect 226978 191128 226984 191140
rect 184808 191100 226984 191128
rect 184808 191088 184814 191100
rect 226978 191088 226984 191100
rect 227036 191088 227042 191140
rect 213178 189728 213184 189780
rect 213236 189768 213242 189780
rect 265066 189768 265072 189780
rect 213236 189740 265072 189768
rect 213236 189728 213242 189740
rect 265066 189728 265072 189740
rect 265124 189728 265130 189780
rect 3418 188844 3424 188896
rect 3476 188884 3482 188896
rect 7650 188884 7656 188896
rect 3476 188856 7656 188884
rect 3476 188844 3482 188856
rect 7650 188844 7656 188856
rect 7708 188844 7714 188896
rect 194502 188300 194508 188352
rect 194560 188340 194566 188352
rect 223574 188340 223580 188352
rect 194560 188312 223580 188340
rect 194560 188300 194566 188312
rect 223574 188300 223580 188312
rect 223632 188300 223638 188352
rect 231118 188300 231124 188352
rect 231176 188340 231182 188352
rect 263778 188340 263784 188352
rect 231176 188312 263784 188340
rect 231176 188300 231182 188312
rect 263778 188300 263784 188312
rect 263836 188300 263842 188352
rect 60550 187688 60556 187740
rect 60608 187728 60614 187740
rect 60608 187700 185808 187728
rect 60608 187688 60614 187700
rect 185780 187660 185808 187700
rect 186222 187660 186228 187672
rect 185780 187632 186228 187660
rect 186222 187620 186228 187632
rect 186280 187660 186286 187672
rect 232498 187660 232504 187672
rect 186280 187632 232504 187660
rect 186280 187620 186286 187632
rect 232498 187620 232504 187632
rect 232556 187620 232562 187672
rect 44082 186260 44088 186312
rect 44140 186300 44146 186312
rect 292574 186300 292580 186312
rect 44140 186272 292580 186300
rect 44140 186260 44146 186272
rect 292574 186260 292580 186272
rect 292632 186260 292638 186312
rect 90910 184152 90916 184204
rect 90968 184192 90974 184204
rect 121546 184192 121552 184204
rect 90968 184164 121552 184192
rect 90968 184152 90974 184164
rect 121546 184152 121552 184164
rect 121604 184152 121610 184204
rect 193490 184152 193496 184204
rect 193548 184192 193554 184204
rect 225966 184192 225972 184204
rect 193548 184164 225972 184192
rect 193548 184152 193554 184164
rect 225966 184152 225972 184164
rect 226024 184152 226030 184204
rect 183462 182792 183468 182844
rect 183520 182832 183526 182844
rect 295334 182832 295340 182844
rect 183520 182804 295340 182832
rect 183520 182792 183526 182804
rect 295334 182792 295340 182804
rect 295392 182792 295398 182844
rect 181530 181500 181536 181552
rect 181588 181540 181594 181552
rect 201494 181540 201500 181552
rect 181588 181512 201500 181540
rect 181588 181500 181594 181512
rect 201494 181500 201500 181512
rect 201552 181500 201558 181552
rect 84102 181432 84108 181484
rect 84160 181472 84166 181484
rect 106458 181472 106464 181484
rect 84160 181444 106464 181472
rect 84160 181432 84166 181444
rect 106458 181432 106464 181444
rect 106516 181432 106522 181484
rect 198090 181432 198096 181484
rect 198148 181472 198154 181484
rect 244918 181472 244924 181484
rect 198148 181444 244924 181472
rect 198148 181432 198154 181444
rect 244918 181432 244924 181444
rect 244976 181432 244982 181484
rect 12342 180072 12348 180124
rect 12400 180112 12406 180124
rect 153930 180112 153936 180124
rect 12400 180084 153936 180112
rect 12400 180072 12406 180084
rect 153930 180072 153936 180084
rect 153988 180072 153994 180124
rect 206278 180072 206284 180124
rect 206336 180112 206342 180124
rect 226518 180112 226524 180124
rect 206336 180084 226524 180112
rect 206336 180072 206342 180084
rect 226518 180072 226524 180084
rect 226576 180072 226582 180124
rect 87598 178644 87604 178696
rect 87656 178684 87662 178696
rect 120074 178684 120080 178696
rect 87656 178656 120080 178684
rect 87656 178644 87662 178656
rect 120074 178644 120080 178656
rect 120132 178644 120138 178696
rect 236730 178644 236736 178696
rect 236788 178684 236794 178696
rect 237282 178684 237288 178696
rect 236788 178656 237288 178684
rect 236788 178644 236794 178656
rect 237282 178644 237288 178656
rect 237340 178684 237346 178696
rect 580166 178684 580172 178696
rect 237340 178656 580172 178684
rect 237340 178644 237346 178656
rect 580166 178644 580172 178656
rect 580224 178644 580230 178696
rect 95970 178032 95976 178084
rect 96028 178072 96034 178084
rect 101490 178072 101496 178084
rect 96028 178044 101496 178072
rect 96028 178032 96034 178044
rect 101490 178032 101496 178044
rect 101548 178032 101554 178084
rect 88242 177284 88248 177336
rect 88300 177324 88306 177336
rect 204898 177324 204904 177336
rect 88300 177296 204904 177324
rect 88300 177284 88306 177296
rect 204898 177284 204904 177296
rect 204956 177284 204962 177336
rect 209958 177284 209964 177336
rect 210016 177324 210022 177336
rect 274726 177324 274732 177336
rect 210016 177296 274732 177324
rect 210016 177284 210022 177296
rect 274726 177284 274732 177296
rect 274784 177284 274790 177336
rect 87598 176672 87604 176724
rect 87656 176712 87662 176724
rect 88242 176712 88248 176724
rect 87656 176684 88248 176712
rect 87656 176672 87662 176684
rect 88242 176672 88248 176684
rect 88300 176672 88306 176724
rect 91186 176672 91192 176724
rect 91244 176712 91250 176724
rect 220814 176712 220820 176724
rect 91244 176684 220820 176712
rect 91244 176672 91250 176684
rect 220814 176672 220820 176684
rect 220872 176712 220878 176724
rect 221458 176712 221464 176724
rect 220872 176684 221464 176712
rect 220872 176672 220878 176684
rect 221458 176672 221464 176684
rect 221516 176672 221522 176724
rect 222838 176332 222844 176384
rect 222896 176372 222902 176384
rect 224954 176372 224960 176384
rect 222896 176344 224960 176372
rect 222896 176332 222902 176344
rect 224954 176332 224960 176344
rect 225012 176332 225018 176384
rect 88978 175924 88984 175976
rect 89036 175964 89042 175976
rect 105538 175964 105544 175976
rect 89036 175936 105544 175964
rect 89036 175924 89042 175936
rect 105538 175924 105544 175936
rect 105596 175924 105602 175976
rect 117958 175244 117964 175296
rect 118016 175284 118022 175296
rect 213270 175284 213276 175296
rect 118016 175256 213276 175284
rect 118016 175244 118022 175256
rect 213270 175244 213276 175256
rect 213328 175244 213334 175296
rect 203518 174496 203524 174548
rect 203576 174536 203582 174548
rect 281626 174536 281632 174548
rect 203576 174508 281632 174536
rect 203576 174496 203582 174508
rect 281626 174496 281632 174508
rect 281684 174536 281690 174548
rect 306374 174536 306380 174548
rect 281684 174508 306380 174536
rect 281684 174496 281690 174508
rect 306374 174496 306380 174508
rect 306432 174496 306438 174548
rect 89714 173884 89720 173936
rect 89772 173924 89778 173936
rect 90818 173924 90824 173936
rect 89772 173896 90824 173924
rect 89772 173884 89778 173896
rect 90818 173884 90824 173896
rect 90876 173924 90882 173936
rect 220078 173924 220084 173936
rect 90876 173896 220084 173924
rect 90876 173884 90882 173896
rect 220078 173884 220084 173896
rect 220136 173884 220142 173936
rect 223574 173000 223580 173052
rect 223632 173040 223638 173052
rect 224310 173040 224316 173052
rect 223632 173012 224316 173040
rect 223632 173000 223638 173012
rect 224310 173000 224316 173012
rect 224368 173000 224374 173052
rect 145650 172592 145656 172644
rect 145708 172632 145714 172644
rect 223574 172632 223580 172644
rect 145708 172604 223580 172632
rect 145708 172592 145714 172604
rect 223574 172592 223580 172604
rect 223632 172592 223638 172644
rect 89162 172524 89168 172576
rect 89220 172564 89226 172576
rect 201494 172564 201500 172576
rect 89220 172536 201500 172564
rect 89220 172524 89226 172536
rect 201494 172524 201500 172536
rect 201552 172524 201558 172576
rect 253198 172524 253204 172576
rect 253256 172564 253262 172576
rect 583018 172564 583024 172576
rect 253256 172536 583024 172564
rect 253256 172524 253262 172536
rect 583018 172524 583024 172536
rect 583076 172524 583082 172576
rect 194778 172456 194784 172508
rect 194836 172496 194842 172508
rect 195330 172496 195336 172508
rect 194836 172468 195336 172496
rect 194836 172456 194842 172468
rect 195330 172456 195336 172468
rect 195388 172456 195394 172508
rect 189718 171844 189724 171896
rect 189776 171884 189782 171896
rect 288710 171884 288716 171896
rect 189776 171856 288716 171884
rect 189776 171844 189782 171856
rect 288710 171844 288716 171856
rect 288768 171844 288774 171896
rect 56410 171776 56416 171828
rect 56468 171816 56474 171828
rect 194778 171816 194784 171828
rect 56468 171788 194784 171816
rect 56468 171776 56474 171788
rect 194778 171776 194784 171788
rect 194836 171776 194842 171828
rect 201494 171028 201500 171080
rect 201552 171068 201558 171080
rect 269114 171068 269120 171080
rect 201552 171040 269120 171068
rect 201552 171028 201558 171040
rect 269114 171028 269120 171040
rect 269172 171028 269178 171080
rect 76650 170348 76656 170400
rect 76708 170388 76714 170400
rect 202966 170388 202972 170400
rect 76708 170360 202972 170388
rect 76708 170348 76714 170360
rect 202966 170348 202972 170360
rect 203024 170388 203030 170400
rect 203518 170388 203524 170400
rect 203024 170360 203524 170388
rect 203024 170348 203030 170360
rect 203518 170348 203524 170360
rect 203576 170348 203582 170400
rect 75914 169736 75920 169788
rect 75972 169776 75978 169788
rect 76650 169776 76656 169788
rect 75972 169748 76656 169776
rect 75972 169736 75978 169748
rect 76650 169736 76656 169748
rect 76708 169736 76714 169788
rect 195974 168376 195980 168428
rect 196032 168416 196038 168428
rect 196618 168416 196624 168428
rect 196032 168388 196624 168416
rect 196032 168376 196038 168388
rect 196618 168376 196624 168388
rect 196676 168416 196682 168428
rect 300118 168416 300124 168428
rect 196676 168388 300124 168416
rect 196676 168376 196682 168388
rect 300118 168376 300124 168388
rect 300176 168376 300182 168428
rect 177942 167628 177948 167680
rect 178000 167668 178006 167680
rect 191190 167668 191196 167680
rect 178000 167640 191196 167668
rect 178000 167628 178006 167640
rect 191190 167628 191196 167640
rect 191248 167628 191254 167680
rect 215386 167628 215392 167680
rect 215444 167668 215450 167680
rect 259546 167668 259552 167680
rect 215444 167640 259552 167668
rect 215444 167628 215450 167640
rect 259546 167628 259552 167640
rect 259604 167628 259610 167680
rect 135990 167016 135996 167068
rect 136048 167056 136054 167068
rect 215294 167056 215300 167068
rect 136048 167028 215300 167056
rect 136048 167016 136054 167028
rect 215294 167016 215300 167028
rect 215352 167016 215358 167068
rect 186314 166336 186320 166388
rect 186372 166376 186378 166388
rect 187602 166376 187608 166388
rect 186372 166348 187608 166376
rect 186372 166336 186378 166348
rect 187602 166336 187608 166348
rect 187660 166376 187666 166388
rect 198090 166376 198096 166388
rect 187660 166348 198096 166376
rect 187660 166336 187666 166348
rect 198090 166336 198096 166348
rect 198148 166336 198154 166388
rect 82906 166268 82912 166320
rect 82964 166308 82970 166320
rect 177850 166308 177856 166320
rect 82964 166280 177856 166308
rect 82964 166268 82970 166280
rect 177850 166268 177856 166280
rect 177908 166308 177914 166320
rect 207658 166308 207664 166320
rect 177908 166280 207664 166308
rect 177908 166268 177914 166280
rect 207658 166268 207664 166280
rect 207716 166268 207722 166320
rect 63310 165588 63316 165640
rect 63368 165628 63374 165640
rect 186314 165628 186320 165640
rect 63368 165600 186320 165628
rect 63368 165588 63374 165600
rect 186314 165588 186320 165600
rect 186372 165588 186378 165640
rect 215294 164840 215300 164892
rect 215352 164880 215358 164892
rect 231854 164880 231860 164892
rect 215352 164852 231860 164880
rect 215352 164840 215358 164852
rect 231854 164840 231860 164852
rect 231912 164840 231918 164892
rect 123478 164296 123484 164348
rect 123536 164336 123542 164348
rect 233234 164336 233240 164348
rect 123536 164308 233240 164336
rect 123536 164296 123542 164308
rect 233234 164296 233240 164308
rect 233292 164296 233298 164348
rect 86954 164228 86960 164280
rect 87012 164268 87018 164280
rect 215938 164268 215944 164280
rect 87012 164240 215944 164268
rect 87012 164228 87018 164240
rect 215938 164228 215944 164240
rect 215996 164228 216002 164280
rect 60458 164160 60464 164212
rect 60516 164200 60522 164212
rect 60642 164200 60648 164212
rect 60516 164172 60648 164200
rect 60516 164160 60522 164172
rect 60642 164160 60648 164172
rect 60700 164160 60706 164212
rect 189074 164160 189080 164212
rect 189132 164200 189138 164212
rect 189718 164200 189724 164212
rect 189132 164172 189724 164200
rect 189132 164160 189138 164172
rect 189718 164160 189724 164172
rect 189776 164160 189782 164212
rect 200114 163888 200120 163940
rect 200172 163928 200178 163940
rect 204990 163928 204996 163940
rect 200172 163900 204996 163928
rect 200172 163888 200178 163900
rect 204990 163888 204996 163900
rect 205048 163888 205054 163940
rect 60458 163480 60464 163532
rect 60516 163520 60522 163532
rect 189074 163520 189080 163532
rect 60516 163492 189080 163520
rect 60516 163480 60522 163492
rect 189074 163480 189080 163492
rect 189132 163480 189138 163532
rect 222194 163480 222200 163532
rect 222252 163520 222258 163532
rect 276014 163520 276020 163532
rect 222252 163492 276020 163520
rect 222252 163480 222258 163492
rect 276014 163480 276020 163492
rect 276072 163480 276078 163532
rect 87138 162868 87144 162920
rect 87196 162908 87202 162920
rect 215386 162908 215392 162920
rect 87196 162880 215392 162908
rect 87196 162868 87202 162880
rect 215386 162868 215392 162880
rect 215444 162868 215450 162920
rect 235994 162800 236000 162852
rect 236052 162840 236058 162852
rect 236730 162840 236736 162852
rect 236052 162812 236736 162840
rect 236052 162800 236058 162812
rect 236730 162800 236736 162812
rect 236788 162800 236794 162852
rect 247126 162120 247132 162172
rect 247184 162160 247190 162172
rect 280522 162160 280528 162172
rect 247184 162132 280528 162160
rect 247184 162120 247190 162132
rect 280522 162120 280528 162132
rect 280580 162160 280586 162172
rect 340138 162160 340144 162172
rect 280580 162132 340144 162160
rect 280580 162120 280586 162132
rect 340138 162120 340144 162132
rect 340196 162120 340202 162172
rect 183002 161508 183008 161560
rect 183060 161548 183066 161560
rect 235994 161548 236000 161560
rect 183060 161520 236000 161548
rect 183060 161508 183066 161520
rect 235994 161508 236000 161520
rect 236052 161508 236058 161560
rect 147030 161440 147036 161492
rect 147088 161480 147094 161492
rect 224954 161480 224960 161492
rect 147088 161452 224960 161480
rect 147088 161440 147094 161452
rect 224954 161440 224960 161452
rect 225012 161440 225018 161492
rect 191926 161372 191932 161424
rect 191984 161412 191990 161424
rect 247126 161412 247132 161424
rect 191984 161384 247132 161412
rect 191984 161372 191990 161384
rect 247126 161372 247132 161384
rect 247184 161372 247190 161424
rect 91002 160692 91008 160744
rect 91060 160732 91066 160744
rect 109034 160732 109040 160744
rect 91060 160704 109040 160732
rect 91060 160692 91066 160704
rect 109034 160692 109040 160704
rect 109092 160732 109098 160744
rect 220170 160732 220176 160744
rect 109092 160704 220176 160732
rect 109092 160692 109098 160704
rect 220170 160692 220176 160704
rect 220228 160692 220234 160744
rect 183462 160080 183468 160132
rect 183520 160120 183526 160132
rect 184198 160120 184204 160132
rect 183520 160092 184204 160120
rect 183520 160080 183526 160092
rect 184198 160080 184204 160092
rect 184256 160080 184262 160132
rect 191650 160080 191656 160132
rect 191708 160120 191714 160132
rect 191926 160120 191932 160132
rect 191708 160092 191932 160120
rect 191708 160080 191714 160092
rect 191926 160080 191932 160092
rect 191984 160080 191990 160132
rect 220354 160080 220360 160132
rect 220412 160120 220418 160132
rect 302234 160120 302240 160132
rect 220412 160092 302240 160120
rect 220412 160080 220418 160092
rect 302234 160080 302240 160092
rect 302292 160080 302298 160132
rect 208578 159332 208584 159384
rect 208636 159372 208642 159384
rect 270586 159372 270592 159384
rect 208636 159344 270592 159372
rect 208636 159332 208642 159344
rect 270586 159332 270592 159344
rect 270644 159332 270650 159384
rect 255406 158924 255412 158976
rect 255464 158964 255470 158976
rect 255958 158964 255964 158976
rect 255464 158936 255964 158964
rect 255464 158924 255470 158936
rect 255958 158924 255964 158936
rect 256016 158924 256022 158976
rect 88978 158788 88984 158840
rect 89036 158828 89042 158840
rect 127710 158828 127716 158840
rect 89036 158800 127716 158828
rect 89036 158788 89042 158800
rect 127710 158788 127716 158800
rect 127768 158788 127774 158840
rect 153930 158788 153936 158840
rect 153988 158828 153994 158840
rect 255406 158828 255412 158840
rect 153988 158800 255412 158828
rect 153988 158788 153994 158800
rect 255406 158788 255412 158800
rect 255464 158788 255470 158840
rect 64690 158720 64696 158772
rect 64748 158760 64754 158772
rect 193122 158760 193128 158772
rect 64748 158732 193128 158760
rect 64748 158720 64754 158732
rect 193122 158720 193128 158732
rect 193180 158720 193186 158772
rect 75270 157972 75276 158024
rect 75328 158012 75334 158024
rect 89162 158012 89168 158024
rect 75328 157984 89168 158012
rect 75328 157972 75334 157984
rect 89162 157972 89168 157984
rect 89220 157972 89226 158024
rect 127710 157972 127716 158024
rect 127768 158012 127774 158024
rect 220814 158012 220820 158024
rect 127768 157984 220820 158012
rect 127768 157972 127774 157984
rect 220814 157972 220820 157984
rect 220872 157972 220878 158024
rect 61930 157360 61936 157412
rect 61988 157400 61994 157412
rect 191742 157400 191748 157412
rect 61988 157372 191748 157400
rect 61988 157360 61994 157372
rect 191742 157360 191748 157372
rect 191800 157360 191806 157412
rect 214558 157360 214564 157412
rect 214616 157400 214622 157412
rect 215110 157400 215116 157412
rect 214616 157372 215116 157400
rect 214616 157360 214622 157372
rect 215110 157360 215116 157372
rect 215168 157400 215174 157412
rect 582742 157400 582748 157412
rect 215168 157372 582748 157400
rect 215168 157360 215174 157372
rect 582742 157360 582748 157372
rect 582800 157360 582806 157412
rect 65978 156612 65984 156664
rect 66036 156652 66042 156664
rect 163590 156652 163596 156664
rect 66036 156624 163596 156652
rect 66036 156612 66042 156624
rect 163590 156612 163596 156624
rect 163648 156612 163654 156664
rect 209866 156408 209872 156460
rect 209924 156448 209930 156460
rect 210418 156448 210424 156460
rect 209924 156420 210424 156448
rect 209924 156408 209930 156420
rect 210418 156408 210424 156420
rect 210476 156408 210482 156460
rect 152642 156000 152648 156052
rect 152700 156040 152706 156052
rect 256970 156040 256976 156052
rect 152700 156012 256976 156040
rect 152700 156000 152706 156012
rect 256970 156000 256976 156012
rect 257028 156000 257034 156052
rect 210418 155932 210424 155984
rect 210476 155972 210482 155984
rect 582374 155972 582380 155984
rect 210476 155944 582380 155972
rect 210476 155932 210482 155944
rect 582374 155932 582380 155944
rect 582432 155932 582438 155984
rect 191558 155864 191564 155916
rect 191616 155904 191622 155916
rect 191742 155904 191748 155916
rect 191616 155876 191748 155904
rect 191616 155864 191622 155876
rect 191742 155864 191748 155876
rect 191800 155904 191806 155916
rect 230474 155904 230480 155916
rect 191800 155876 230480 155904
rect 191800 155864 191806 155876
rect 230474 155864 230480 155876
rect 230532 155904 230538 155916
rect 231762 155904 231768 155916
rect 230532 155876 231768 155904
rect 230532 155864 230538 155876
rect 231762 155864 231768 155876
rect 231820 155864 231826 155916
rect 231762 155252 231768 155304
rect 231820 155292 231826 155304
rect 243630 155292 243636 155304
rect 231820 155264 243636 155292
rect 231820 155252 231826 155264
rect 243630 155252 243636 155264
rect 243688 155252 243694 155304
rect 37090 155184 37096 155236
rect 37148 155224 37154 155236
rect 48130 155224 48136 155236
rect 37148 155196 48136 155224
rect 37148 155184 37154 155196
rect 48130 155184 48136 155196
rect 48188 155184 48194 155236
rect 249794 155224 249800 155236
rect 103486 155196 249800 155224
rect 97258 155116 97264 155168
rect 97316 155156 97322 155168
rect 97810 155156 97816 155168
rect 97316 155128 97816 155156
rect 97316 155116 97322 155128
rect 97810 155116 97816 155128
rect 97868 155156 97874 155168
rect 103486 155156 103514 155196
rect 249794 155184 249800 155196
rect 249852 155224 249858 155236
rect 250530 155224 250536 155236
rect 249852 155196 250536 155224
rect 249852 155184 249858 155196
rect 250530 155184 250536 155196
rect 250588 155184 250594 155236
rect 97868 155128 103514 155156
rect 97868 155116 97874 155128
rect 48130 154572 48136 154624
rect 48188 154612 48194 154624
rect 186958 154612 186964 154624
rect 48188 154584 186964 154612
rect 48188 154572 48194 154584
rect 186958 154572 186964 154584
rect 187016 154572 187022 154624
rect 164234 154504 164240 154556
rect 164292 154544 164298 154556
rect 165062 154544 165068 154556
rect 164292 154516 165068 154544
rect 164292 154504 164298 154516
rect 165062 154504 165068 154516
rect 165120 154504 165126 154556
rect 193122 154504 193128 154556
rect 193180 154544 193186 154556
rect 218054 154544 218060 154556
rect 193180 154516 218060 154544
rect 193180 154504 193186 154516
rect 218054 154504 218060 154516
rect 218112 154504 218118 154556
rect 61654 153824 61660 153876
rect 61712 153864 61718 153876
rect 75178 153864 75184 153876
rect 61712 153836 75184 153864
rect 61712 153824 61718 153836
rect 75178 153824 75184 153836
rect 75236 153824 75242 153876
rect 65886 153280 65892 153332
rect 65944 153320 65950 153332
rect 165062 153320 165068 153332
rect 65944 153292 165068 153320
rect 65944 153280 65950 153292
rect 165062 153280 165068 153292
rect 165120 153280 165126 153332
rect 93854 153212 93860 153264
rect 93912 153252 93918 153264
rect 95050 153252 95056 153264
rect 93912 153224 95056 153252
rect 93912 153212 93918 153224
rect 95050 153212 95056 153224
rect 95108 153252 95114 153264
rect 223574 153252 223580 153264
rect 95108 153224 223580 153252
rect 95108 153212 95114 153224
rect 223574 153212 223580 153224
rect 223632 153212 223638 153264
rect 239950 153212 239956 153264
rect 240008 153252 240014 153264
rect 333974 153252 333980 153264
rect 240008 153224 333980 153252
rect 240008 153212 240014 153224
rect 333974 153212 333980 153224
rect 334032 153212 334038 153264
rect 60642 152532 60648 152584
rect 60700 152572 60706 152584
rect 82078 152572 82084 152584
rect 60700 152544 82084 152572
rect 60700 152532 60706 152544
rect 82078 152532 82084 152544
rect 82136 152532 82142 152584
rect 207014 152532 207020 152584
rect 207072 152572 207078 152584
rect 220354 152572 220360 152584
rect 207072 152544 220360 152572
rect 207072 152532 207078 152544
rect 220354 152532 220360 152544
rect 220412 152532 220418 152584
rect 64598 152464 64604 152516
rect 64656 152504 64662 152516
rect 64782 152504 64788 152516
rect 64656 152476 64788 152504
rect 64656 152464 64662 152476
rect 64782 152464 64788 152476
rect 64840 152504 64846 152516
rect 190454 152504 190460 152516
rect 64840 152476 190460 152504
rect 64840 152464 64846 152476
rect 190454 152464 190460 152476
rect 190512 152504 190518 152516
rect 191098 152504 191104 152516
rect 190512 152476 191104 152504
rect 190512 152464 190518 152476
rect 191098 152464 191104 152476
rect 191156 152464 191162 152516
rect 191190 152464 191196 152516
rect 191248 152504 191254 152516
rect 239950 152504 239956 152516
rect 191248 152476 239956 152504
rect 191248 152464 191254 152476
rect 239950 152464 239956 152476
rect 240008 152464 240014 152516
rect 161474 151784 161480 151836
rect 161532 151824 161538 151836
rect 162578 151824 162584 151836
rect 161532 151796 162584 151824
rect 161532 151784 161538 151796
rect 162578 151784 162584 151796
rect 162636 151824 162642 151836
rect 185762 151824 185768 151836
rect 162636 151796 185768 151824
rect 162636 151784 162642 151796
rect 185762 151784 185768 151796
rect 185820 151784 185826 151836
rect 281442 151716 281448 151768
rect 281500 151756 281506 151768
rect 291470 151756 291476 151768
rect 281500 151728 291476 151756
rect 281500 151716 281506 151728
rect 291470 151716 291476 151728
rect 291528 151716 291534 151768
rect 81986 151036 81992 151088
rect 82044 151076 82050 151088
rect 104894 151076 104900 151088
rect 82044 151048 104900 151076
rect 82044 151036 82050 151048
rect 104894 151036 104900 151048
rect 104952 151036 104958 151088
rect 199286 151036 199292 151088
rect 199344 151076 199350 151088
rect 263962 151076 263968 151088
rect 199344 151048 263968 151076
rect 199344 151036 199350 151048
rect 263962 151036 263968 151048
rect 264020 151036 264026 151088
rect 131850 150532 131856 150544
rect 64846 150504 131856 150532
rect 61746 150424 61752 150476
rect 61804 150464 61810 150476
rect 62022 150464 62028 150476
rect 61804 150436 62028 150464
rect 61804 150424 61810 150436
rect 62022 150424 62028 150436
rect 62080 150464 62086 150476
rect 64846 150464 64874 150504
rect 131850 150492 131856 150504
rect 131908 150492 131914 150544
rect 62080 150436 64874 150464
rect 62080 150424 62086 150436
rect 126882 150424 126888 150476
rect 126940 150464 126946 150476
rect 216674 150464 216680 150476
rect 126940 150436 216680 150464
rect 126940 150424 126946 150436
rect 216674 150424 216680 150436
rect 216732 150424 216738 150476
rect 201402 149676 201408 149728
rect 201460 149716 201466 149728
rect 271874 149716 271880 149728
rect 201460 149688 271880 149716
rect 201460 149676 201466 149688
rect 271874 149676 271880 149688
rect 271932 149676 271938 149728
rect 218054 149268 218060 149320
rect 218112 149308 218118 149320
rect 218606 149308 218612 149320
rect 218112 149280 218612 149308
rect 218112 149268 218118 149280
rect 218606 149268 218612 149280
rect 218664 149268 218670 149320
rect 73062 149132 73068 149184
rect 73120 149172 73126 149184
rect 199286 149172 199292 149184
rect 73120 149144 199292 149172
rect 73120 149132 73126 149144
rect 199286 149132 199292 149144
rect 199344 149132 199350 149184
rect 55030 149064 55036 149116
rect 55088 149104 55094 149116
rect 181438 149104 181444 149116
rect 55088 149076 181444 149104
rect 55088 149064 55094 149076
rect 181438 149064 181444 149076
rect 181496 149064 181502 149116
rect 204530 149064 204536 149116
rect 204588 149104 204594 149116
rect 244918 149104 244924 149116
rect 204588 149076 244924 149104
rect 204588 149064 204594 149076
rect 244918 149064 244924 149076
rect 244976 149064 244982 149116
rect 53742 148316 53748 148368
rect 53800 148356 53806 148368
rect 182818 148356 182824 148368
rect 53800 148328 182824 148356
rect 53800 148316 53806 148328
rect 182818 148316 182824 148328
rect 182876 148316 182882 148368
rect 184658 148316 184664 148368
rect 184716 148356 184722 148368
rect 191834 148356 191840 148368
rect 184716 148328 191840 148356
rect 184716 148316 184722 148328
rect 191834 148316 191840 148328
rect 191892 148316 191898 148368
rect 206922 147704 206928 147756
rect 206980 147744 206986 147756
rect 232498 147744 232504 147756
rect 206980 147716 232504 147744
rect 206980 147704 206986 147716
rect 232498 147704 232504 147716
rect 232556 147704 232562 147756
rect 98730 147636 98736 147688
rect 98788 147676 98794 147688
rect 99282 147676 99288 147688
rect 98788 147648 99288 147676
rect 98788 147636 98794 147648
rect 99282 147636 99288 147648
rect 99340 147676 99346 147688
rect 224954 147676 224960 147688
rect 99340 147648 224960 147676
rect 99340 147636 99346 147648
rect 224954 147636 224960 147648
rect 225012 147636 225018 147688
rect 207658 147568 207664 147620
rect 207716 147608 207722 147620
rect 211154 147608 211160 147620
rect 207716 147580 211160 147608
rect 207716 147568 207722 147580
rect 211154 147568 211160 147580
rect 211212 147568 211218 147620
rect 227806 147160 227812 147212
rect 227864 147160 227870 147212
rect 192478 147024 192484 147076
rect 192536 147064 192542 147076
rect 215478 147064 215484 147076
rect 192536 147036 215484 147064
rect 192536 147024 192542 147036
rect 215478 147024 215484 147036
rect 215536 147024 215542 147076
rect 3418 146956 3424 147008
rect 3476 146996 3482 147008
rect 88242 146996 88248 147008
rect 3476 146968 88248 146996
rect 3476 146956 3482 146968
rect 88242 146956 88248 146968
rect 88300 146956 88306 147008
rect 108482 146956 108488 147008
rect 108540 146996 108546 147008
rect 108942 146996 108948 147008
rect 108540 146968 108948 146996
rect 108540 146956 108546 146968
rect 108942 146956 108948 146968
rect 109000 146996 109006 147008
rect 197906 146996 197912 147008
rect 109000 146968 197912 146996
rect 109000 146956 109006 146968
rect 197906 146956 197912 146968
rect 197964 146956 197970 147008
rect 208394 146956 208400 147008
rect 208452 146996 208458 147008
rect 208854 146996 208860 147008
rect 208452 146968 208860 146996
rect 208452 146956 208458 146968
rect 208854 146956 208860 146968
rect 208912 146956 208918 147008
rect 209866 146956 209872 147008
rect 209924 146996 209930 147008
rect 210694 146996 210700 147008
rect 209924 146968 210700 146996
rect 209924 146956 209930 146968
rect 210694 146956 210700 146968
rect 210752 146956 210758 147008
rect 215386 146956 215392 147008
rect 215444 146996 215450 147008
rect 216214 146996 216220 147008
rect 215444 146968 216220 146996
rect 215444 146956 215450 146968
rect 216214 146956 216220 146968
rect 216272 146956 216278 147008
rect 223574 146956 223580 147008
rect 223632 146996 223638 147008
rect 224494 146996 224500 147008
rect 223632 146968 224500 146996
rect 223632 146956 223638 146968
rect 224494 146956 224500 146968
rect 224552 146956 224558 147008
rect 227714 146956 227720 147008
rect 227772 146996 227778 147008
rect 227824 146996 227852 147160
rect 227772 146968 227852 146996
rect 227772 146956 227778 146968
rect 57790 146888 57796 146940
rect 57848 146928 57854 146940
rect 181530 146928 181536 146940
rect 57848 146900 181536 146928
rect 57848 146888 57854 146900
rect 181530 146888 181536 146900
rect 181588 146888 181594 146940
rect 213454 146888 213460 146940
rect 213512 146928 213518 146940
rect 257982 146928 257988 146940
rect 213512 146900 257988 146928
rect 213512 146888 213518 146900
rect 257982 146888 257988 146900
rect 258040 146928 258046 146940
rect 258810 146928 258816 146940
rect 258040 146900 258816 146928
rect 258040 146888 258046 146900
rect 258810 146888 258816 146900
rect 258868 146888 258874 146940
rect 252462 146276 252468 146328
rect 252520 146316 252526 146328
rect 341518 146316 341524 146328
rect 252520 146288 341524 146316
rect 252520 146276 252526 146288
rect 341518 146276 341524 146288
rect 341576 146276 341582 146328
rect 87506 146208 87512 146260
rect 87564 146248 87570 146260
rect 88242 146248 88248 146260
rect 87564 146220 88248 146248
rect 87564 146208 87570 146220
rect 88242 146208 88248 146220
rect 88300 146248 88306 146260
rect 126882 146248 126888 146260
rect 88300 146220 126888 146248
rect 88300 146208 88306 146220
rect 126882 146208 126888 146220
rect 126940 146208 126946 146260
rect 184290 146208 184296 146260
rect 184348 146248 184354 146260
rect 184842 146248 184848 146260
rect 184348 146220 184848 146248
rect 184348 146208 184354 146220
rect 184842 146208 184848 146220
rect 184900 146208 184906 146260
rect 220170 146208 220176 146260
rect 220228 146248 220234 146260
rect 220906 146248 220912 146260
rect 220228 146220 220912 146248
rect 220228 146208 220234 146220
rect 220906 146208 220912 146220
rect 220964 146208 220970 146260
rect 192570 145528 192576 145580
rect 192628 145568 192634 145580
rect 245102 145568 245108 145580
rect 192628 145540 245108 145568
rect 192628 145528 192634 145540
rect 245102 145528 245108 145540
rect 245160 145568 245166 145580
rect 338114 145568 338120 145580
rect 245160 145540 338120 145568
rect 245160 145528 245166 145540
rect 338114 145528 338120 145540
rect 338172 145528 338178 145580
rect 67358 144916 67364 144968
rect 67416 144956 67422 144968
rect 109770 144956 109776 144968
rect 67416 144928 109776 144956
rect 67416 144916 67422 144928
rect 109770 144916 109776 144928
rect 109828 144916 109834 144968
rect 184290 144916 184296 144968
rect 184348 144956 184354 144968
rect 217226 144956 217232 144968
rect 184348 144928 217232 144956
rect 184348 144916 184354 144928
rect 217226 144916 217232 144928
rect 217284 144916 217290 144968
rect 80146 144780 80152 144832
rect 80204 144820 80210 144832
rect 83458 144820 83464 144832
rect 80204 144792 83464 144820
rect 80204 144780 80210 144792
rect 83458 144780 83464 144792
rect 83516 144780 83522 144832
rect 85574 144440 85580 144492
rect 85632 144480 85638 144492
rect 89070 144480 89076 144492
rect 85632 144452 89076 144480
rect 85632 144440 85638 144452
rect 89070 144440 89076 144452
rect 89128 144440 89134 144492
rect 240778 144168 240784 144220
rect 240836 144208 240842 144220
rect 258718 144208 258724 144220
rect 240836 144180 258724 144208
rect 240836 144168 240842 144180
rect 258718 144168 258724 144180
rect 258776 144168 258782 144220
rect 286778 144168 286784 144220
rect 286836 144208 286842 144220
rect 295334 144208 295340 144220
rect 286836 144180 295340 144208
rect 286836 144168 286842 144180
rect 295334 144168 295340 144180
rect 295392 144168 295398 144220
rect 97350 144032 97356 144084
rect 97408 144072 97414 144084
rect 99374 144072 99380 144084
rect 97408 144044 99380 144072
rect 97408 144032 97414 144044
rect 99374 144032 99380 144044
rect 99432 144032 99438 144084
rect 82814 143692 82820 143744
rect 82872 143732 82878 143744
rect 86310 143732 86316 143744
rect 82872 143704 86316 143732
rect 82872 143692 82878 143704
rect 86310 143692 86316 143704
rect 86368 143692 86374 143744
rect 161474 143624 161480 143676
rect 161532 143664 161538 143676
rect 162670 143664 162676 143676
rect 161532 143636 162676 143664
rect 161532 143624 161538 143636
rect 162670 143624 162676 143636
rect 162728 143664 162734 143676
rect 194134 143664 194140 143676
rect 162728 143636 194140 143664
rect 162728 143624 162734 143636
rect 194134 143624 194140 143636
rect 194192 143624 194198 143676
rect 204990 143624 204996 143676
rect 205048 143664 205054 143676
rect 209774 143664 209780 143676
rect 205048 143636 209780 143664
rect 205048 143624 205054 143636
rect 209774 143624 209780 143636
rect 209832 143624 209838 143676
rect 63126 143556 63132 143608
rect 63184 143596 63190 143608
rect 182910 143596 182916 143608
rect 63184 143568 182916 143596
rect 63184 143556 63190 143568
rect 182910 143556 182916 143568
rect 182968 143556 182974 143608
rect 187142 143556 187148 143608
rect 187200 143596 187206 143608
rect 225230 143596 225236 143608
rect 187200 143568 225236 143596
rect 187200 143556 187206 143568
rect 225230 143556 225236 143568
rect 225288 143556 225294 143608
rect 219526 143488 219532 143540
rect 219584 143528 219590 143540
rect 220262 143528 220268 143540
rect 219584 143500 220268 143528
rect 219584 143488 219590 143500
rect 220262 143488 220268 143500
rect 220320 143488 220326 143540
rect 240778 143528 240784 143540
rect 229066 143500 240784 143528
rect 220078 143420 220084 143472
rect 220136 143460 220142 143472
rect 229066 143460 229094 143500
rect 240778 143488 240784 143500
rect 240836 143488 240842 143540
rect 220136 143432 229094 143460
rect 220136 143420 220142 143432
rect 214006 143216 214012 143268
rect 214064 143256 214070 143268
rect 215110 143256 215116 143268
rect 214064 143228 215116 143256
rect 214064 143216 214070 143228
rect 215110 143216 215116 143228
rect 215168 143216 215174 143268
rect 53558 142808 53564 142860
rect 53616 142848 53622 142860
rect 53616 142820 64874 142848
rect 53616 142808 53622 142820
rect 64846 142780 64874 142820
rect 223666 142808 223672 142860
rect 223724 142848 223730 142860
rect 245010 142848 245016 142860
rect 223724 142820 245016 142848
rect 223724 142808 223730 142820
rect 245010 142808 245016 142820
rect 245068 142808 245074 142860
rect 69014 142780 69020 142792
rect 64846 142752 69020 142780
rect 69014 142740 69020 142752
rect 69072 142780 69078 142792
rect 70578 142780 70584 142792
rect 69072 142752 70584 142780
rect 69072 142740 69078 142752
rect 70578 142740 70584 142752
rect 70636 142740 70642 142792
rect 223206 142536 223212 142588
rect 223264 142576 223270 142588
rect 223666 142576 223672 142588
rect 223264 142548 223672 142576
rect 223264 142536 223270 142548
rect 223666 142536 223672 142548
rect 223724 142536 223730 142588
rect 57698 142332 57704 142384
rect 57756 142372 57762 142384
rect 89898 142372 89904 142384
rect 57756 142344 89904 142372
rect 57756 142332 57762 142344
rect 89898 142332 89904 142344
rect 89956 142332 89962 142384
rect 88610 142264 88616 142316
rect 88668 142304 88674 142316
rect 218238 142304 218244 142316
rect 88668 142276 218244 142304
rect 88668 142264 88674 142276
rect 218238 142264 218244 142276
rect 218296 142264 218302 142316
rect 90910 142196 90916 142248
rect 90968 142236 90974 142248
rect 213454 142236 213460 142248
rect 90968 142208 213460 142236
rect 90968 142196 90974 142208
rect 213454 142196 213460 142208
rect 213512 142196 213518 142248
rect 215294 142128 215300 142180
rect 215352 142168 215358 142180
rect 223482 142168 223488 142180
rect 215352 142140 223488 142168
rect 215352 142128 215358 142140
rect 223482 142128 223488 142140
rect 223540 142128 223546 142180
rect 63402 141380 63408 141432
rect 63460 141420 63466 141432
rect 77294 141420 77300 141432
rect 63460 141392 77300 141420
rect 63460 141380 63466 141392
rect 77294 141380 77300 141392
rect 77352 141380 77358 141432
rect 88518 141380 88524 141432
rect 88576 141420 88582 141432
rect 184290 141420 184296 141432
rect 88576 141392 184296 141420
rect 88576 141380 88582 141392
rect 184290 141380 184296 141392
rect 184348 141380 184354 141432
rect 223022 140972 223028 141024
rect 223080 141012 223086 141024
rect 227990 141012 227996 141024
rect 223080 140984 227996 141012
rect 223080 140972 223086 140984
rect 227990 140972 227996 140984
rect 228048 140972 228054 141024
rect 21358 140768 21364 140820
rect 21416 140808 21422 140820
rect 88978 140808 88984 140820
rect 21416 140780 88984 140808
rect 21416 140768 21422 140780
rect 88978 140768 88984 140780
rect 89036 140768 89042 140820
rect 193306 140768 193312 140820
rect 193364 140808 193370 140820
rect 196618 140808 196624 140820
rect 193364 140780 196624 140808
rect 193364 140768 193370 140780
rect 196618 140768 196624 140780
rect 196676 140768 196682 140820
rect 203426 140768 203432 140820
rect 203484 140808 203490 140820
rect 289078 140808 289084 140820
rect 203484 140780 289084 140808
rect 203484 140768 203490 140780
rect 289078 140768 289084 140780
rect 289136 140768 289142 140820
rect 223482 140700 223488 140752
rect 223540 140740 223546 140752
rect 251818 140740 251824 140752
rect 223540 140712 251824 140740
rect 223540 140700 223546 140712
rect 251818 140700 251824 140712
rect 251876 140700 251882 140752
rect 200086 140576 209774 140604
rect 193030 140428 193036 140480
rect 193088 140468 193094 140480
rect 194778 140468 194784 140480
rect 193088 140440 194784 140468
rect 193088 140428 193094 140440
rect 194778 140428 194784 140440
rect 194836 140428 194842 140480
rect 78030 140020 78036 140072
rect 78088 140060 78094 140072
rect 87598 140060 87604 140072
rect 78088 140032 87604 140060
rect 78088 140020 78094 140032
rect 87598 140020 87604 140032
rect 87656 140020 87662 140072
rect 89898 139476 89904 139528
rect 89956 139516 89962 139528
rect 96154 139516 96160 139528
rect 89956 139488 96160 139516
rect 89956 139476 89962 139488
rect 96154 139476 96160 139488
rect 96212 139476 96218 139528
rect 86862 139408 86868 139460
rect 86920 139448 86926 139460
rect 200086 139448 200114 140576
rect 205174 140536 205180 140548
rect 86920 139420 200114 139448
rect 204180 140508 205180 140536
rect 86920 139408 86926 139420
rect 84746 139340 84752 139392
rect 84804 139380 84810 139392
rect 90910 139380 90916 139392
rect 84804 139352 90916 139380
rect 84804 139340 84810 139352
rect 90910 139340 90916 139352
rect 90968 139340 90974 139392
rect 204180 139380 204208 140508
rect 205174 140496 205180 140508
rect 205232 140496 205238 140548
rect 209746 140468 209774 140576
rect 210050 140496 210056 140548
rect 210108 140536 210114 140548
rect 210108 140508 219434 140536
rect 210108 140496 210114 140508
rect 215386 140468 215392 140480
rect 209746 140440 215392 140468
rect 215386 140428 215392 140440
rect 215444 140428 215450 140480
rect 219406 140060 219434 140508
rect 287698 140060 287704 140072
rect 219406 140032 287704 140060
rect 287698 140020 287704 140032
rect 287756 140020 287762 140072
rect 251266 139748 251272 139800
rect 251324 139788 251330 139800
rect 251818 139788 251824 139800
rect 251324 139760 251824 139788
rect 251324 139748 251330 139760
rect 251818 139748 251824 139760
rect 251876 139748 251882 139800
rect 200086 139352 204208 139380
rect 193398 138660 193404 138712
rect 193456 138700 193462 138712
rect 200086 138700 200114 139352
rect 225322 138932 225328 138984
rect 225380 138972 225386 138984
rect 227714 138972 227720 138984
rect 225380 138944 227720 138972
rect 225380 138932 225386 138944
rect 227714 138932 227720 138944
rect 227772 138932 227778 138984
rect 193456 138672 200114 138700
rect 193456 138660 193462 138672
rect 70210 138116 70216 138168
rect 70268 138156 70274 138168
rect 71866 138156 71872 138168
rect 70268 138128 71872 138156
rect 70268 138116 70274 138128
rect 71866 138116 71872 138128
rect 71924 138116 71930 138168
rect 70394 138048 70400 138100
rect 70452 138088 70458 138100
rect 71222 138088 71228 138100
rect 70452 138060 71228 138088
rect 70452 138048 70458 138060
rect 71222 138048 71228 138060
rect 71280 138048 71286 138100
rect 73338 138048 73344 138100
rect 73396 138088 73402 138100
rect 73798 138088 73804 138100
rect 73396 138060 73804 138088
rect 73396 138048 73402 138060
rect 73798 138048 73804 138060
rect 73856 138048 73862 138100
rect 88334 138048 88340 138100
rect 88392 138088 88398 138100
rect 89254 138088 89260 138100
rect 88392 138060 89260 138088
rect 88392 138048 88398 138060
rect 89254 138048 89260 138060
rect 89312 138048 89318 138100
rect 67910 137980 67916 138032
rect 67968 138020 67974 138032
rect 159450 138020 159456 138032
rect 67968 137992 159456 138020
rect 67968 137980 67974 137992
rect 159450 137980 159456 137992
rect 159508 137980 159514 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 3292 137924 70394 137952
rect 3292 137912 3298 137924
rect 70366 137884 70394 137924
rect 73062 137884 73068 137896
rect 70366 137856 73068 137884
rect 73062 137844 73068 137856
rect 73120 137844 73126 137896
rect 88978 137708 88984 137760
rect 89036 137748 89042 137760
rect 91186 137748 91192 137760
rect 89036 137720 91192 137748
rect 89036 137708 89042 137720
rect 91186 137708 91192 137720
rect 91244 137708 91250 137760
rect 173342 137232 173348 137284
rect 173400 137272 173406 137284
rect 183002 137272 183008 137284
rect 173400 137244 183008 137272
rect 173400 137232 173406 137244
rect 183002 137232 183008 137244
rect 183060 137232 183066 137284
rect 79962 136824 79968 136876
rect 80020 136864 80026 136876
rect 80974 136864 80980 136876
rect 80020 136836 80980 136864
rect 80020 136824 80026 136836
rect 80974 136824 80980 136836
rect 81032 136824 81038 136876
rect 76558 136688 76564 136740
rect 76616 136728 76622 136740
rect 77386 136728 77392 136740
rect 76616 136700 77392 136728
rect 76616 136688 76622 136700
rect 77386 136688 77392 136700
rect 77444 136688 77450 136740
rect 85482 136688 85488 136740
rect 85540 136728 85546 136740
rect 86218 136728 86224 136740
rect 85540 136700 86224 136728
rect 85540 136688 85546 136700
rect 86218 136688 86224 136700
rect 86276 136688 86282 136740
rect 66070 136620 66076 136672
rect 66128 136660 66134 136672
rect 94498 136660 94504 136672
rect 66128 136632 94504 136660
rect 66128 136620 66134 136632
rect 94498 136620 94504 136632
rect 94556 136620 94562 136672
rect 182818 136620 182824 136672
rect 182876 136660 182882 136672
rect 191650 136660 191656 136672
rect 182876 136632 191656 136660
rect 182876 136620 182882 136632
rect 191650 136620 191656 136632
rect 191708 136620 191714 136672
rect 173802 136552 173808 136604
rect 173860 136592 173866 136604
rect 191742 136592 191748 136604
rect 173860 136564 191748 136592
rect 173860 136552 173866 136564
rect 191742 136552 191748 136564
rect 191800 136552 191806 136604
rect 54478 135940 54484 135992
rect 54536 135980 54542 135992
rect 90818 135980 90824 135992
rect 54536 135952 90824 135980
rect 54536 135940 54542 135952
rect 90818 135940 90824 135952
rect 90876 135980 90882 135992
rect 91278 135980 91284 135992
rect 90876 135952 91284 135980
rect 90876 135940 90882 135952
rect 91278 135940 91284 135952
rect 91336 135940 91342 135992
rect 64782 135872 64788 135924
rect 64840 135912 64846 135924
rect 69658 135912 69664 135924
rect 64840 135884 69664 135912
rect 64840 135872 64846 135884
rect 69658 135872 69664 135884
rect 69716 135872 69722 135924
rect 70302 135872 70308 135924
rect 70360 135912 70366 135924
rect 161474 135912 161480 135924
rect 70360 135884 161480 135912
rect 70360 135872 70366 135884
rect 161474 135872 161480 135884
rect 161532 135872 161538 135924
rect 226518 135872 226524 135924
rect 226576 135912 226582 135924
rect 239398 135912 239404 135924
rect 226576 135884 239404 135912
rect 226576 135872 226582 135884
rect 239398 135872 239404 135884
rect 239456 135872 239462 135924
rect 243630 135872 243636 135924
rect 243688 135912 243694 135924
rect 304258 135912 304264 135924
rect 243688 135884 304264 135912
rect 243688 135872 243694 135884
rect 304258 135872 304264 135884
rect 304316 135872 304322 135924
rect 226518 135600 226524 135652
rect 226576 135640 226582 135652
rect 230474 135640 230480 135652
rect 226576 135612 230480 135640
rect 226576 135600 226582 135612
rect 230474 135600 230480 135612
rect 230532 135600 230538 135652
rect 160738 135260 160744 135312
rect 160796 135300 160802 135312
rect 191742 135300 191748 135312
rect 160796 135272 191748 135300
rect 160796 135260 160802 135272
rect 191742 135260 191748 135272
rect 191800 135260 191806 135312
rect 94498 135192 94504 135244
rect 94556 135232 94562 135244
rect 192478 135232 192484 135244
rect 94556 135204 192484 135232
rect 94556 135192 94562 135204
rect 192478 135192 192484 135204
rect 192536 135192 192542 135244
rect 232498 135192 232504 135244
rect 232556 135232 232562 135244
rect 249058 135232 249064 135244
rect 232556 135204 249064 135232
rect 232556 135192 232562 135204
rect 249058 135192 249064 135204
rect 249116 135192 249122 135244
rect 96798 135124 96804 135176
rect 96856 135164 96862 135176
rect 188522 135164 188528 135176
rect 96856 135136 188528 135164
rect 96856 135124 96862 135136
rect 188522 135124 188528 135136
rect 188580 135124 188586 135176
rect 93762 134580 93768 134632
rect 93820 134620 93826 134632
rect 95234 134620 95240 134632
rect 93820 134592 95240 134620
rect 93820 134580 93826 134592
rect 95234 134580 95240 134592
rect 95292 134580 95298 134632
rect 247678 134512 247684 134564
rect 247736 134552 247742 134564
rect 298738 134552 298744 134564
rect 247736 134524 298744 134552
rect 247736 134512 247742 134524
rect 298738 134512 298744 134524
rect 298796 134512 298802 134564
rect 96614 133832 96620 133884
rect 96672 133872 96678 133884
rect 102870 133872 102876 133884
rect 96672 133844 102876 133872
rect 96672 133832 96678 133844
rect 102870 133832 102876 133844
rect 102928 133832 102934 133884
rect 188430 133832 188436 133884
rect 188488 133872 188494 133884
rect 191742 133872 191748 133884
rect 188488 133844 191748 133872
rect 188488 133832 188494 133844
rect 191742 133832 191748 133844
rect 191800 133832 191806 133884
rect 226702 133832 226708 133884
rect 226760 133872 226766 133884
rect 229278 133872 229284 133884
rect 226760 133844 229284 133872
rect 226760 133832 226766 133844
rect 229278 133832 229284 133844
rect 229336 133832 229342 133884
rect 268010 133872 268016 133884
rect 238726 133844 268016 133872
rect 226886 133764 226892 133816
rect 226944 133804 226950 133816
rect 227898 133804 227904 133816
rect 226944 133776 227904 133804
rect 226944 133764 226950 133776
rect 227898 133764 227904 133776
rect 227956 133804 227962 133816
rect 238726 133804 238754 133844
rect 268010 133832 268016 133844
rect 268068 133832 268074 133884
rect 227956 133776 238754 133804
rect 227956 133764 227962 133776
rect 103054 133220 103060 133272
rect 103112 133260 103118 133272
rect 160830 133260 160836 133272
rect 103112 133232 160836 133260
rect 103112 133220 103118 133232
rect 160830 133220 160836 133232
rect 160888 133220 160894 133272
rect 56410 133152 56416 133204
rect 56468 133192 56474 133204
rect 66346 133192 66352 133204
rect 56468 133164 66352 133192
rect 56468 133152 56474 133164
rect 66346 133152 66352 133164
rect 66404 133152 66410 133204
rect 110874 133152 110880 133204
rect 110932 133192 110938 133204
rect 187142 133192 187148 133204
rect 110932 133164 187148 133192
rect 110932 133152 110938 133164
rect 187142 133152 187148 133164
rect 187200 133152 187206 133204
rect 50982 132404 50988 132456
rect 51040 132444 51046 132456
rect 66898 132444 66904 132456
rect 51040 132416 66904 132444
rect 51040 132404 51046 132416
rect 66898 132404 66904 132416
rect 66956 132404 66962 132456
rect 96154 132404 96160 132456
rect 96212 132444 96218 132456
rect 191190 132444 191196 132456
rect 96212 132416 191196 132444
rect 96212 132404 96218 132416
rect 191190 132404 191196 132416
rect 191248 132404 191254 132456
rect 226702 132404 226708 132456
rect 226760 132444 226766 132456
rect 229094 132444 229100 132456
rect 226760 132416 229100 132444
rect 226760 132404 226766 132416
rect 229094 132404 229100 132416
rect 229152 132404 229158 132456
rect 96614 132336 96620 132388
rect 96672 132376 96678 132388
rect 148502 132376 148508 132388
rect 96672 132348 148508 132376
rect 96672 132336 96678 132348
rect 148502 132336 148508 132348
rect 148560 132336 148566 132388
rect 187602 131452 187608 131504
rect 187660 131492 187666 131504
rect 192938 131492 192944 131504
rect 187660 131464 192944 131492
rect 187660 131452 187666 131464
rect 192938 131452 192944 131464
rect 192996 131452 193002 131504
rect 165062 131044 165068 131096
rect 165120 131084 165126 131096
rect 182818 131084 182824 131096
rect 165120 131056 182824 131084
rect 165120 131044 165126 131056
rect 182818 131044 182824 131056
rect 182876 131044 182882 131096
rect 225414 131044 225420 131096
rect 225472 131084 225478 131096
rect 273254 131084 273260 131096
rect 225472 131056 273260 131084
rect 225472 131044 225478 131056
rect 273254 131044 273260 131056
rect 273312 131044 273318 131096
rect 226610 130976 226616 131028
rect 226668 131016 226674 131028
rect 256694 131016 256700 131028
rect 226668 130988 256700 131016
rect 226668 130976 226674 130988
rect 256694 130976 256700 130988
rect 256752 130976 256758 131028
rect 96614 130364 96620 130416
rect 96672 130404 96678 130416
rect 170582 130404 170588 130416
rect 96672 130376 170588 130404
rect 96672 130364 96678 130376
rect 170582 130364 170588 130376
rect 170640 130364 170646 130416
rect 96614 130160 96620 130212
rect 96672 130200 96678 130212
rect 102962 130200 102968 130212
rect 96672 130172 102968 130200
rect 96672 130160 96678 130172
rect 102962 130160 102968 130172
rect 103020 130160 103026 130212
rect 127710 129888 127716 129940
rect 127768 129928 127774 129940
rect 133138 129928 133144 129940
rect 127768 129900 133144 129928
rect 127768 129888 127774 129900
rect 133138 129888 133144 129900
rect 133196 129888 133202 129940
rect 186314 129752 186320 129804
rect 186372 129792 186378 129804
rect 191006 129792 191012 129804
rect 186372 129764 191012 129792
rect 186372 129752 186378 129764
rect 191006 129752 191012 129764
rect 191064 129752 191070 129804
rect 159450 129684 159456 129736
rect 159508 129724 159514 129736
rect 185486 129724 185492 129736
rect 159508 129696 185492 129724
rect 159508 129684 159514 129696
rect 185486 129684 185492 129696
rect 185544 129724 185550 129736
rect 185670 129724 185676 129736
rect 185544 129696 185676 129724
rect 185544 129684 185550 129696
rect 185670 129684 185676 129696
rect 185728 129684 185734 129736
rect 227162 129276 227168 129328
rect 227220 129316 227226 129328
rect 227990 129316 227996 129328
rect 227220 129288 227996 129316
rect 227220 129276 227226 129288
rect 227990 129276 227996 129288
rect 228048 129276 228054 129328
rect 104342 129004 104348 129056
rect 104400 129044 104406 129056
rect 191466 129044 191472 129056
rect 104400 129016 191472 129044
rect 104400 129004 104406 129016
rect 191466 129004 191472 129016
rect 191524 129044 191530 129056
rect 192570 129044 192576 129056
rect 191524 129016 192576 129044
rect 191524 129004 191530 129016
rect 192570 129004 192576 129016
rect 192628 129004 192634 129056
rect 230382 129004 230388 129056
rect 230440 129044 230446 129056
rect 249794 129044 249800 129056
rect 230440 129016 249800 129044
rect 230440 129004 230446 129016
rect 249794 129004 249800 129016
rect 249852 129004 249858 129056
rect 187602 128392 187608 128444
rect 187660 128432 187666 128444
rect 189074 128432 189080 128444
rect 187660 128404 189080 128432
rect 187660 128392 187666 128404
rect 189074 128392 189080 128404
rect 189132 128432 189138 128444
rect 191190 128432 191196 128444
rect 189132 128404 191196 128432
rect 189132 128392 189138 128404
rect 191190 128392 191196 128404
rect 191248 128392 191254 128444
rect 226150 128324 226156 128376
rect 226208 128364 226214 128376
rect 299474 128364 299480 128376
rect 226208 128336 299480 128364
rect 226208 128324 226214 128336
rect 299474 128324 299480 128336
rect 299532 128324 299538 128376
rect 48130 128256 48136 128308
rect 48188 128296 48194 128308
rect 66898 128296 66904 128308
rect 48188 128268 66904 128296
rect 48188 128256 48194 128268
rect 66898 128256 66904 128268
rect 66956 128256 66962 128308
rect 97534 128256 97540 128308
rect 97592 128296 97598 128308
rect 127802 128296 127808 128308
rect 97592 128268 127808 128296
rect 97592 128256 97598 128268
rect 127802 128256 127808 128268
rect 127860 128256 127866 128308
rect 163590 128256 163596 128308
rect 163648 128296 163654 128308
rect 191742 128296 191748 128308
rect 163648 128268 191748 128296
rect 163648 128256 163654 128268
rect 191742 128256 191748 128268
rect 191800 128256 191806 128308
rect 226610 128256 226616 128308
rect 226668 128296 226674 128308
rect 231854 128296 231860 128308
rect 226668 128268 231860 128296
rect 226668 128256 226674 128268
rect 231854 128256 231860 128268
rect 231912 128296 231918 128308
rect 233142 128296 233148 128308
rect 231912 128268 233148 128296
rect 231912 128256 231918 128268
rect 233142 128256 233148 128268
rect 233200 128256 233206 128308
rect 227990 127644 227996 127696
rect 228048 127684 228054 127696
rect 267826 127684 267832 127696
rect 228048 127656 267832 127684
rect 228048 127644 228054 127656
rect 267826 127644 267832 127656
rect 267884 127644 267890 127696
rect 97074 127576 97080 127628
rect 97132 127616 97138 127628
rect 183094 127616 183100 127628
rect 97132 127588 183100 127616
rect 97132 127576 97138 127588
rect 183094 127576 183100 127588
rect 183152 127576 183158 127628
rect 233142 127576 233148 127628
rect 233200 127616 233206 127628
rect 331858 127616 331864 127628
rect 233200 127588 331864 127616
rect 233200 127576 233206 127588
rect 331858 127576 331864 127588
rect 331916 127576 331922 127628
rect 57606 126896 57612 126948
rect 57664 126936 57670 126948
rect 66806 126936 66812 126948
rect 57664 126908 66812 126936
rect 57664 126896 57670 126908
rect 66806 126896 66812 126908
rect 66864 126896 66870 126948
rect 97810 126896 97816 126948
rect 97868 126936 97874 126948
rect 110874 126936 110880 126948
rect 97868 126908 110880 126936
rect 97868 126896 97874 126908
rect 110874 126896 110880 126908
rect 110932 126896 110938 126948
rect 226426 126896 226432 126948
rect 226484 126936 226490 126948
rect 255406 126936 255412 126948
rect 226484 126908 255412 126936
rect 226484 126896 226490 126908
rect 255406 126896 255412 126908
rect 255464 126896 255470 126948
rect 63310 126828 63316 126880
rect 63368 126868 63374 126880
rect 66714 126868 66720 126880
rect 63368 126840 66720 126868
rect 63368 126828 63374 126840
rect 66714 126828 66720 126840
rect 66772 126828 66778 126880
rect 226886 126828 226892 126880
rect 226944 126868 226950 126880
rect 227530 126868 227536 126880
rect 226944 126840 227536 126868
rect 226944 126828 226950 126840
rect 227530 126828 227536 126840
rect 227588 126868 227594 126880
rect 230382 126868 230388 126880
rect 227588 126840 230388 126868
rect 227588 126828 227594 126840
rect 230382 126828 230388 126840
rect 230440 126828 230446 126880
rect 126330 126284 126336 126336
rect 126388 126324 126394 126336
rect 141602 126324 141608 126336
rect 126388 126296 141608 126324
rect 126388 126284 126394 126296
rect 141602 126284 141608 126296
rect 141660 126284 141666 126336
rect 108390 126216 108396 126268
rect 108448 126256 108454 126268
rect 191650 126256 191656 126268
rect 108448 126228 191656 126256
rect 108448 126216 108454 126228
rect 191650 126216 191656 126228
rect 191708 126256 191714 126268
rect 193398 126256 193404 126268
rect 191708 126228 193404 126256
rect 191708 126216 191714 126228
rect 193398 126216 193404 126228
rect 193456 126216 193462 126268
rect 98454 125536 98460 125588
rect 98512 125576 98518 125588
rect 152642 125576 152648 125588
rect 98512 125548 152648 125576
rect 98512 125536 98518 125548
rect 152642 125536 152648 125548
rect 152700 125536 152706 125588
rect 166350 125536 166356 125588
rect 166408 125576 166414 125588
rect 186314 125576 186320 125588
rect 166408 125548 186320 125576
rect 166408 125536 166414 125548
rect 186314 125536 186320 125548
rect 186372 125536 186378 125588
rect 226610 125536 226616 125588
rect 226668 125576 226674 125588
rect 259454 125576 259460 125588
rect 226668 125548 259460 125576
rect 226668 125536 226674 125548
rect 259454 125536 259460 125548
rect 259512 125536 259518 125588
rect 115198 124856 115204 124908
rect 115256 124896 115262 124908
rect 127618 124896 127624 124908
rect 115256 124868 127624 124896
rect 115256 124856 115262 124868
rect 127618 124856 127624 124868
rect 127676 124856 127682 124908
rect 60458 124788 60464 124840
rect 60516 124828 60522 124840
rect 66622 124828 66628 124840
rect 60516 124800 66628 124828
rect 60516 124788 60522 124800
rect 66622 124788 66628 124800
rect 66680 124788 66686 124840
rect 57698 124108 57704 124160
rect 57756 124148 57762 124160
rect 66254 124148 66260 124160
rect 57756 124120 66260 124148
rect 57756 124108 57762 124120
rect 66254 124108 66260 124120
rect 66312 124108 66318 124160
rect 97810 124108 97816 124160
rect 97868 124148 97874 124160
rect 147030 124148 147036 124160
rect 97868 124120 147036 124148
rect 97868 124108 97874 124120
rect 147030 124108 147036 124120
rect 147088 124108 147094 124160
rect 180058 124108 180064 124160
rect 180116 124148 180122 124160
rect 191006 124148 191012 124160
rect 180116 124120 191012 124148
rect 180116 124108 180122 124120
rect 191006 124108 191012 124120
rect 191064 124108 191070 124160
rect 226702 124108 226708 124160
rect 226760 124148 226766 124160
rect 233234 124148 233240 124160
rect 226760 124120 233240 124148
rect 226760 124108 226766 124120
rect 233234 124108 233240 124120
rect 233292 124148 233298 124160
rect 288526 124148 288532 124160
rect 233292 124120 288532 124148
rect 233292 124108 233298 124120
rect 288526 124108 288532 124120
rect 288584 124148 288590 124160
rect 582926 124148 582932 124160
rect 288584 124120 582932 124148
rect 288584 124108 288590 124120
rect 582926 124108 582932 124120
rect 582984 124108 582990 124160
rect 97166 124040 97172 124092
rect 97224 124080 97230 124092
rect 135990 124080 135996 124092
rect 97224 124052 135996 124080
rect 97224 124040 97230 124052
rect 135990 124040 135996 124052
rect 136048 124040 136054 124092
rect 226518 123836 226524 123888
rect 226576 123876 226582 123888
rect 229186 123876 229192 123888
rect 226576 123848 229192 123876
rect 226576 123836 226582 123848
rect 229186 123836 229192 123848
rect 229244 123836 229250 123888
rect 162118 123428 162124 123480
rect 162176 123468 162182 123480
rect 173250 123468 173256 123480
rect 162176 123440 173256 123468
rect 162176 123428 162182 123440
rect 173250 123428 173256 123440
rect 173308 123428 173314 123480
rect 97534 122748 97540 122800
rect 97592 122788 97598 122800
rect 153930 122788 153936 122800
rect 97592 122760 153936 122788
rect 97592 122748 97598 122760
rect 153930 122748 153936 122760
rect 153988 122748 153994 122800
rect 226518 122748 226524 122800
rect 226576 122788 226582 122800
rect 235994 122788 236000 122800
rect 226576 122760 236000 122788
rect 226576 122748 226582 122760
rect 235994 122748 236000 122760
rect 236052 122748 236058 122800
rect 181530 122068 181536 122120
rect 181588 122108 181594 122120
rect 181990 122108 181996 122120
rect 181588 122080 181996 122108
rect 181588 122068 181594 122080
rect 181990 122068 181996 122080
rect 182048 122108 182054 122120
rect 191742 122108 191748 122120
rect 182048 122080 191748 122108
rect 182048 122068 182054 122080
rect 191742 122068 191748 122080
rect 191800 122068 191806 122120
rect 226978 122068 226984 122120
rect 227036 122108 227042 122120
rect 309778 122108 309784 122120
rect 227036 122080 309784 122108
rect 227036 122068 227042 122080
rect 309778 122068 309784 122080
rect 309836 122068 309842 122120
rect 54938 121388 54944 121440
rect 54996 121428 55002 121440
rect 66898 121428 66904 121440
rect 54996 121400 66904 121428
rect 54996 121388 55002 121400
rect 66898 121388 66904 121400
rect 66956 121388 66962 121440
rect 96982 121388 96988 121440
rect 97040 121428 97046 121440
rect 103054 121428 103060 121440
rect 97040 121400 103060 121428
rect 97040 121388 97046 121400
rect 103054 121388 103060 121400
rect 103112 121388 103118 121440
rect 185762 121388 185768 121440
rect 185820 121428 185826 121440
rect 191742 121428 191748 121440
rect 185820 121400 191748 121428
rect 185820 121388 185826 121400
rect 191742 121388 191748 121400
rect 191800 121388 191806 121440
rect 226702 121388 226708 121440
rect 226760 121428 226766 121440
rect 240134 121428 240140 121440
rect 226760 121400 240140 121428
rect 226760 121388 226766 121400
rect 240134 121388 240140 121400
rect 240192 121388 240198 121440
rect 61930 121320 61936 121372
rect 61988 121360 61994 121372
rect 66806 121360 66812 121372
rect 61988 121332 66812 121360
rect 61988 121320 61994 121332
rect 66806 121320 66812 121332
rect 66864 121320 66870 121372
rect 110322 120776 110328 120828
rect 110380 120816 110386 120828
rect 142982 120816 142988 120828
rect 110380 120788 142988 120816
rect 110380 120776 110386 120788
rect 142982 120776 142988 120788
rect 143040 120776 143046 120828
rect 108390 120708 108396 120760
rect 108448 120748 108454 120760
rect 124858 120748 124864 120760
rect 108448 120720 124864 120748
rect 108448 120708 108454 120720
rect 124858 120708 124864 120720
rect 124916 120708 124922 120760
rect 131850 120708 131856 120760
rect 131908 120748 131914 120760
rect 187694 120748 187700 120760
rect 131908 120720 187700 120748
rect 131908 120708 131914 120720
rect 187694 120708 187700 120720
rect 187752 120708 187758 120760
rect 239398 120708 239404 120760
rect 239456 120748 239462 120760
rect 282178 120748 282184 120760
rect 239456 120720 282184 120748
rect 239456 120708 239462 120720
rect 282178 120708 282184 120720
rect 282236 120708 282242 120760
rect 96062 120300 96068 120352
rect 96120 120340 96126 120352
rect 98822 120340 98828 120352
rect 96120 120312 98828 120340
rect 96120 120300 96126 120312
rect 98822 120300 98828 120312
rect 98880 120300 98886 120352
rect 187694 120164 187700 120216
rect 187752 120204 187758 120216
rect 188982 120204 188988 120216
rect 187752 120176 188988 120204
rect 187752 120164 187758 120176
rect 188982 120164 188988 120176
rect 189040 120204 189046 120216
rect 191742 120204 191748 120216
rect 189040 120176 191748 120204
rect 189040 120164 189046 120176
rect 191742 120164 191748 120176
rect 191800 120164 191806 120216
rect 53650 120028 53656 120080
rect 53708 120068 53714 120080
rect 66898 120068 66904 120080
rect 53708 120040 66904 120068
rect 53708 120028 53714 120040
rect 66898 120028 66904 120040
rect 66956 120028 66962 120080
rect 97902 120028 97908 120080
rect 97960 120068 97966 120080
rect 123478 120068 123484 120080
rect 97960 120040 123484 120068
rect 97960 120028 97966 120040
rect 123478 120028 123484 120040
rect 123536 120028 123542 120080
rect 181438 120028 181444 120080
rect 181496 120068 181502 120080
rect 191742 120068 191748 120080
rect 181496 120040 191748 120068
rect 181496 120028 181502 120040
rect 191742 120028 191748 120040
rect 191800 120028 191806 120080
rect 64690 119960 64696 120012
rect 64748 120000 64754 120012
rect 66806 120000 66812 120012
rect 64748 119972 66812 120000
rect 64748 119960 64754 119972
rect 66806 119960 66812 119972
rect 66864 119960 66870 120012
rect 109678 118668 109684 118720
rect 109736 118708 109742 118720
rect 173802 118708 173808 118720
rect 109736 118680 173808 118708
rect 109736 118668 109742 118680
rect 173802 118668 173808 118680
rect 173860 118708 173866 118720
rect 174630 118708 174636 118720
rect 173860 118680 174636 118708
rect 173860 118668 173866 118680
rect 174630 118668 174636 118680
rect 174688 118668 174694 118720
rect 57790 118600 57796 118652
rect 57848 118640 57854 118652
rect 66714 118640 66720 118652
rect 57848 118612 66720 118640
rect 57848 118600 57854 118612
rect 66714 118600 66720 118612
rect 66772 118600 66778 118652
rect 97902 118600 97908 118652
rect 97960 118640 97966 118652
rect 173342 118640 173348 118652
rect 97960 118612 173348 118640
rect 97960 118600 97966 118612
rect 173342 118600 173348 118612
rect 173400 118600 173406 118652
rect 181990 118600 181996 118652
rect 182048 118640 182054 118652
rect 184198 118640 184204 118652
rect 182048 118612 184204 118640
rect 182048 118600 182054 118612
rect 184198 118600 184204 118612
rect 184256 118600 184262 118652
rect 181990 117920 181996 117972
rect 182048 117960 182054 117972
rect 191006 117960 191012 117972
rect 182048 117932 191012 117960
rect 182048 117920 182054 117932
rect 191006 117920 191012 117932
rect 191064 117920 191070 117972
rect 227530 117920 227536 117972
rect 227588 117960 227594 117972
rect 353294 117960 353300 117972
rect 227588 117932 353300 117960
rect 227588 117920 227594 117932
rect 353294 117920 353300 117932
rect 353352 117920 353358 117972
rect 99374 117308 99380 117360
rect 99432 117348 99438 117360
rect 100662 117348 100668 117360
rect 99432 117320 100668 117348
rect 99432 117308 99438 117320
rect 100662 117308 100668 117320
rect 100720 117348 100726 117360
rect 108482 117348 108488 117360
rect 100720 117320 108488 117348
rect 100720 117308 100726 117320
rect 108482 117308 108488 117320
rect 108540 117308 108546 117360
rect 226610 117308 226616 117360
rect 226668 117348 226674 117360
rect 252738 117348 252744 117360
rect 226668 117320 252744 117348
rect 226668 117308 226674 117320
rect 252738 117308 252744 117320
rect 252796 117308 252802 117360
rect 64506 117240 64512 117292
rect 64564 117280 64570 117292
rect 66806 117280 66812 117292
rect 64564 117252 66812 117280
rect 64564 117240 64570 117252
rect 66806 117240 66812 117252
rect 66864 117240 66870 117292
rect 97902 117240 97908 117292
rect 97960 117280 97966 117292
rect 177390 117280 177396 117292
rect 97960 117252 177396 117280
rect 97960 117240 97966 117252
rect 177390 117240 177396 117252
rect 177448 117240 177454 117292
rect 182910 117240 182916 117292
rect 182968 117280 182974 117292
rect 191742 117280 191748 117292
rect 182968 117252 191748 117280
rect 182968 117240 182974 117252
rect 191742 117240 191748 117252
rect 191800 117240 191806 117292
rect 61746 117172 61752 117224
rect 61804 117212 61810 117224
rect 66254 117212 66260 117224
rect 61804 117184 66260 117212
rect 61804 117172 61810 117184
rect 66254 117172 66260 117184
rect 66312 117172 66318 117224
rect 97350 117172 97356 117224
rect 97408 117212 97414 117224
rect 155402 117212 155408 117224
rect 97408 117184 155408 117212
rect 97408 117172 97414 117184
rect 155402 117172 155408 117184
rect 155460 117172 155466 117224
rect 188338 117172 188344 117224
rect 188396 117212 188402 117224
rect 191006 117212 191012 117224
rect 188396 117184 191012 117212
rect 188396 117172 188402 117184
rect 191006 117172 191012 117184
rect 191064 117172 191070 117224
rect 226702 116968 226708 117020
rect 226760 117008 226766 117020
rect 230474 117008 230480 117020
rect 226760 116980 230480 117008
rect 226760 116968 226766 116980
rect 230474 116968 230480 116980
rect 230532 117008 230538 117020
rect 231118 117008 231124 117020
rect 230532 116980 231124 117008
rect 230532 116968 230538 116980
rect 231118 116968 231124 116980
rect 231176 116968 231182 117020
rect 230382 116628 230388 116680
rect 230440 116668 230446 116680
rect 262214 116668 262220 116680
rect 230440 116640 262220 116668
rect 230440 116628 230446 116640
rect 262214 116628 262220 116640
rect 262272 116628 262278 116680
rect 231118 116560 231124 116612
rect 231176 116600 231182 116612
rect 281534 116600 281540 116612
rect 231176 116572 281540 116600
rect 231176 116560 231182 116572
rect 281534 116560 281540 116572
rect 281592 116600 281598 116612
rect 304350 116600 304356 116612
rect 281592 116572 304356 116600
rect 281592 116560 281598 116572
rect 304350 116560 304356 116572
rect 304408 116560 304414 116612
rect 226702 115948 226708 116000
rect 226760 115988 226766 116000
rect 229094 115988 229100 116000
rect 226760 115960 229100 115988
rect 226760 115948 226766 115960
rect 229094 115948 229100 115960
rect 229152 115988 229158 116000
rect 230382 115988 230388 116000
rect 229152 115960 230388 115988
rect 229152 115948 229158 115960
rect 230382 115948 230388 115960
rect 230440 115948 230446 116000
rect 55030 115880 55036 115932
rect 55088 115920 55094 115932
rect 66898 115920 66904 115932
rect 55088 115892 66904 115920
rect 55088 115880 55094 115892
rect 66898 115880 66904 115892
rect 66956 115880 66962 115932
rect 97810 115880 97816 115932
rect 97868 115920 97874 115932
rect 99374 115920 99380 115932
rect 97868 115892 99380 115920
rect 97868 115880 97874 115892
rect 99374 115880 99380 115892
rect 99432 115880 99438 115932
rect 180702 115880 180708 115932
rect 180760 115920 180766 115932
rect 190822 115920 190828 115932
rect 180760 115892 190828 115920
rect 180760 115880 180766 115892
rect 190822 115880 190828 115892
rect 190880 115880 190886 115932
rect 64598 115268 64604 115320
rect 64656 115308 64662 115320
rect 66806 115308 66812 115320
rect 64656 115280 66812 115308
rect 64656 115268 64662 115280
rect 66806 115268 66812 115280
rect 66864 115268 66870 115320
rect 233234 115200 233240 115252
rect 233292 115240 233298 115252
rect 277394 115240 277400 115252
rect 233292 115212 277400 115240
rect 233292 115200 233298 115212
rect 277394 115200 277400 115212
rect 277452 115200 277458 115252
rect 97902 114520 97908 114572
rect 97960 114560 97966 114572
rect 169110 114560 169116 114572
rect 97960 114532 169116 114560
rect 97960 114520 97966 114532
rect 169110 114520 169116 114532
rect 169168 114520 169174 114572
rect 226702 114520 226708 114572
rect 226760 114560 226766 114572
rect 233234 114560 233240 114572
rect 226760 114532 233240 114560
rect 226760 114520 226766 114532
rect 233234 114520 233240 114532
rect 233292 114520 233298 114572
rect 8202 114452 8208 114504
rect 8260 114492 8266 114504
rect 8260 114464 45554 114492
rect 8260 114452 8266 114464
rect 45526 114424 45554 114464
rect 59170 114452 59176 114504
rect 59228 114492 59234 114504
rect 66806 114492 66812 114504
rect 59228 114464 66812 114492
rect 59228 114452 59234 114464
rect 66806 114452 66812 114464
rect 66864 114452 66870 114504
rect 226610 114452 226616 114504
rect 226668 114492 226674 114504
rect 242250 114492 242256 114504
rect 226668 114464 242256 114492
rect 226668 114452 226674 114464
rect 242250 114452 242256 114464
rect 242308 114492 242314 114504
rect 250530 114492 250536 114504
rect 242308 114464 250536 114492
rect 242308 114452 242314 114464
rect 250530 114452 250536 114464
rect 250588 114452 250594 114504
rect 63126 114424 63132 114436
rect 45526 114396 63132 114424
rect 63126 114384 63132 114396
rect 63184 114424 63190 114436
rect 66898 114424 66904 114436
rect 63184 114396 66904 114424
rect 63184 114384 63190 114396
rect 66898 114384 66904 114396
rect 66956 114384 66962 114436
rect 97810 113976 97816 114028
rect 97868 114016 97874 114028
rect 101490 114016 101496 114028
rect 97868 113988 101496 114016
rect 97868 113976 97874 113988
rect 101490 113976 101496 113988
rect 101548 113976 101554 114028
rect 235258 113772 235264 113824
rect 235316 113812 235322 113824
rect 242158 113812 242164 113824
rect 235316 113784 242164 113812
rect 235316 113772 235322 113784
rect 242158 113772 242164 113784
rect 242216 113772 242222 113824
rect 97902 113160 97908 113212
rect 97960 113200 97966 113212
rect 173250 113200 173256 113212
rect 97960 113172 173256 113200
rect 97960 113160 97966 113172
rect 173250 113160 173256 113172
rect 173308 113160 173314 113212
rect 188246 113160 188252 113212
rect 188304 113200 188310 113212
rect 191742 113200 191748 113212
rect 188304 113172 191748 113200
rect 188304 113160 188310 113172
rect 191742 113160 191748 113172
rect 191800 113160 191806 113212
rect 52362 112412 52368 112464
rect 52420 112452 52426 112464
rect 66806 112452 66812 112464
rect 52420 112424 66812 112452
rect 52420 112412 52426 112424
rect 66806 112412 66812 112424
rect 66864 112412 66870 112464
rect 157242 112412 157248 112464
rect 157300 112452 157306 112464
rect 191742 112452 191748 112464
rect 157300 112424 191748 112452
rect 157300 112412 157306 112424
rect 191742 112412 191748 112424
rect 191800 112412 191806 112464
rect 97074 111868 97080 111920
rect 97132 111908 97138 111920
rect 100018 111908 100024 111920
rect 97132 111880 100024 111908
rect 97132 111868 97138 111880
rect 100018 111868 100024 111880
rect 100076 111868 100082 111920
rect 98086 111800 98092 111852
rect 98144 111840 98150 111852
rect 100754 111840 100760 111852
rect 98144 111812 100760 111840
rect 98144 111800 98150 111812
rect 100754 111800 100760 111812
rect 100812 111800 100818 111852
rect 156690 111800 156696 111852
rect 156748 111840 156754 111852
rect 157242 111840 157248 111852
rect 156748 111812 157248 111840
rect 156748 111800 156754 111812
rect 157242 111800 157248 111812
rect 157300 111800 157306 111852
rect 226702 111800 226708 111852
rect 226760 111840 226766 111852
rect 231946 111840 231952 111852
rect 226760 111812 231952 111840
rect 226760 111800 226766 111812
rect 231946 111800 231952 111812
rect 232004 111840 232010 111852
rect 324314 111840 324320 111852
rect 232004 111812 324320 111840
rect 232004 111800 232010 111812
rect 324314 111800 324320 111812
rect 324372 111800 324378 111852
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 21358 111772 21364 111784
rect 3476 111744 21364 111772
rect 3476 111732 3482 111744
rect 21358 111732 21364 111744
rect 21416 111732 21422 111784
rect 96706 111664 96712 111716
rect 96764 111704 96770 111716
rect 98730 111704 98736 111716
rect 96764 111676 98736 111704
rect 96764 111664 96770 111676
rect 98730 111664 98736 111676
rect 98788 111664 98794 111716
rect 239398 111120 239404 111172
rect 239456 111160 239462 111172
rect 252646 111160 252652 111172
rect 239456 111132 252652 111160
rect 239456 111120 239462 111132
rect 252646 111120 252652 111132
rect 252704 111120 252710 111172
rect 41138 111052 41144 111104
rect 41196 111092 41202 111104
rect 57146 111092 57152 111104
rect 41196 111064 57152 111092
rect 41196 111052 41202 111064
rect 57146 111052 57152 111064
rect 57204 111052 57210 111104
rect 101582 111052 101588 111104
rect 101640 111092 101646 111104
rect 114646 111092 114652 111104
rect 101640 111064 114652 111092
rect 101640 111052 101646 111064
rect 114646 111052 114652 111064
rect 114704 111052 114710 111104
rect 227070 111052 227076 111104
rect 227128 111092 227134 111104
rect 227714 111092 227720 111104
rect 227128 111064 227720 111092
rect 227128 111052 227134 111064
rect 227714 111052 227720 111064
rect 227772 111092 227778 111104
rect 242158 111092 242164 111104
rect 227772 111064 242164 111092
rect 227772 111052 227778 111064
rect 242158 111052 242164 111064
rect 242216 111052 242222 111104
rect 188890 110508 188896 110560
rect 188948 110548 188954 110560
rect 191834 110548 191840 110560
rect 188948 110520 191840 110548
rect 188948 110508 188954 110520
rect 191834 110508 191840 110520
rect 191892 110508 191898 110560
rect 57146 110440 57152 110492
rect 57204 110480 57210 110492
rect 57790 110480 57796 110492
rect 57204 110452 57796 110480
rect 57204 110440 57210 110452
rect 57790 110440 57796 110452
rect 57848 110480 57854 110492
rect 66806 110480 66812 110492
rect 57848 110452 66812 110480
rect 57848 110440 57854 110452
rect 66806 110440 66812 110452
rect 66864 110440 66870 110492
rect 102042 110480 102048 110492
rect 100772 110452 102048 110480
rect 97902 110372 97908 110424
rect 97960 110412 97966 110424
rect 100772 110412 100800 110452
rect 102042 110440 102048 110452
rect 102100 110480 102106 110492
rect 186958 110480 186964 110492
rect 102100 110452 186964 110480
rect 102100 110440 102106 110452
rect 186958 110440 186964 110452
rect 187016 110440 187022 110492
rect 187694 110440 187700 110492
rect 187752 110480 187758 110492
rect 191742 110480 191748 110492
rect 187752 110452 191748 110480
rect 187752 110440 187758 110452
rect 191742 110440 191748 110452
rect 191800 110440 191806 110492
rect 97960 110384 100800 110412
rect 97960 110372 97966 110384
rect 227714 110372 227720 110424
rect 227772 110412 227778 110424
rect 228358 110412 228364 110424
rect 227772 110384 228364 110412
rect 227772 110372 227778 110384
rect 228358 110372 228364 110384
rect 228416 110412 228422 110424
rect 233878 110412 233884 110424
rect 228416 110384 233884 110412
rect 228416 110372 228422 110384
rect 233878 110372 233884 110384
rect 233936 110372 233942 110424
rect 100110 109692 100116 109744
rect 100168 109732 100174 109744
rect 111794 109732 111800 109744
rect 100168 109704 111800 109732
rect 100168 109692 100174 109704
rect 111794 109692 111800 109704
rect 111852 109692 111858 109744
rect 160830 109692 160836 109744
rect 160888 109732 160894 109744
rect 188246 109732 188252 109744
rect 160888 109704 188252 109732
rect 160888 109692 160894 109704
rect 188246 109692 188252 109704
rect 188304 109692 188310 109744
rect 236730 109692 236736 109744
rect 236788 109732 236794 109744
rect 258074 109732 258080 109744
rect 236788 109704 258080 109732
rect 236788 109692 236794 109704
rect 258074 109692 258080 109704
rect 258132 109692 258138 109744
rect 50890 109012 50896 109064
rect 50948 109052 50954 109064
rect 57238 109052 57244 109064
rect 50948 109024 57244 109052
rect 50948 109012 50954 109024
rect 57238 109012 57244 109024
rect 57296 109052 57302 109064
rect 66806 109052 66812 109064
rect 57296 109024 66812 109052
rect 57296 109012 57302 109024
rect 66806 109012 66812 109024
rect 66864 109012 66870 109064
rect 123478 109012 123484 109064
rect 123536 109052 123542 109064
rect 123536 109024 156644 109052
rect 123536 109012 123542 109024
rect 156616 108996 156644 109024
rect 156598 108944 156604 108996
rect 156656 108984 156662 108996
rect 189074 108984 189080 108996
rect 156656 108956 189080 108984
rect 156656 108944 156662 108956
rect 189074 108944 189080 108956
rect 189132 108944 189138 108996
rect 226426 108944 226432 108996
rect 226484 108984 226490 108996
rect 245654 108984 245660 108996
rect 226484 108956 245660 108984
rect 226484 108944 226490 108956
rect 245654 108944 245660 108956
rect 245712 108944 245718 108996
rect 97902 108332 97908 108384
rect 97960 108372 97966 108384
rect 107470 108372 107476 108384
rect 97960 108344 107476 108372
rect 97960 108332 97966 108344
rect 107470 108332 107476 108344
rect 107528 108332 107534 108384
rect 108482 108332 108488 108384
rect 108540 108372 108546 108384
rect 155402 108372 155408 108384
rect 108540 108344 155408 108372
rect 108540 108332 108546 108344
rect 155402 108332 155408 108344
rect 155460 108332 155466 108384
rect 44082 108264 44088 108316
rect 44140 108304 44146 108316
rect 63494 108304 63500 108316
rect 44140 108276 63500 108304
rect 44140 108264 44146 108276
rect 63494 108264 63500 108276
rect 63552 108264 63558 108316
rect 101674 108264 101680 108316
rect 101732 108304 101738 108316
rect 187694 108304 187700 108316
rect 101732 108276 187700 108304
rect 101732 108264 101738 108276
rect 187694 108264 187700 108276
rect 187752 108264 187758 108316
rect 231762 108264 231768 108316
rect 231820 108304 231826 108316
rect 269206 108304 269212 108316
rect 231820 108276 269212 108304
rect 231820 108264 231826 108276
rect 269206 108264 269212 108276
rect 269264 108264 269270 108316
rect 63494 107652 63500 107704
rect 63552 107692 63558 107704
rect 64598 107692 64604 107704
rect 63552 107664 64604 107692
rect 63552 107652 63558 107664
rect 64598 107652 64604 107664
rect 64656 107692 64662 107704
rect 66806 107692 66812 107704
rect 64656 107664 66812 107692
rect 64656 107652 64662 107664
rect 66806 107652 66812 107664
rect 66864 107652 66870 107704
rect 226702 107652 226708 107704
rect 226760 107692 226766 107704
rect 230566 107692 230572 107704
rect 226760 107664 230572 107692
rect 226760 107652 226766 107664
rect 230566 107652 230572 107664
rect 230624 107692 230630 107704
rect 231762 107692 231768 107704
rect 230624 107664 231768 107692
rect 230624 107652 230630 107664
rect 231762 107652 231768 107664
rect 231820 107652 231826 107704
rect 171870 107584 171876 107636
rect 171928 107624 171934 107636
rect 191742 107624 191748 107636
rect 171928 107596 191748 107624
rect 171928 107584 171934 107596
rect 191742 107584 191748 107596
rect 191800 107584 191806 107636
rect 226794 107584 226800 107636
rect 226852 107624 226858 107636
rect 282914 107624 282920 107636
rect 226852 107596 282920 107624
rect 226852 107584 226858 107596
rect 282914 107584 282920 107596
rect 282972 107584 282978 107636
rect 7558 106904 7564 106956
rect 7616 106944 7622 106956
rect 34330 106944 34336 106956
rect 7616 106916 34336 106944
rect 7616 106904 7622 106916
rect 34330 106904 34336 106916
rect 34388 106944 34394 106956
rect 60734 106944 60740 106956
rect 34388 106916 60740 106944
rect 34388 106904 34394 106916
rect 60734 106904 60740 106916
rect 60792 106904 60798 106956
rect 97810 106904 97816 106956
rect 97868 106944 97874 106956
rect 180058 106944 180064 106956
rect 97868 106916 180064 106944
rect 97868 106904 97874 106916
rect 180058 106904 180064 106916
rect 180116 106904 180122 106956
rect 282914 106904 282920 106956
rect 282972 106944 282978 106956
rect 342898 106944 342904 106956
rect 282972 106916 342904 106944
rect 282972 106904 282978 106916
rect 342898 106904 342904 106916
rect 342956 106904 342962 106956
rect 96706 106360 96712 106412
rect 96764 106400 96770 106412
rect 98730 106400 98736 106412
rect 96764 106372 98736 106400
rect 96764 106360 96770 106372
rect 98730 106360 98736 106372
rect 98788 106360 98794 106412
rect 60734 106292 60740 106344
rect 60792 106332 60798 106344
rect 61930 106332 61936 106344
rect 60792 106304 61936 106332
rect 60792 106292 60798 106304
rect 61930 106292 61936 106304
rect 61988 106332 61994 106344
rect 66806 106332 66812 106344
rect 61988 106304 66812 106332
rect 61988 106292 61994 106304
rect 66806 106292 66812 106304
rect 66864 106292 66870 106344
rect 109770 106224 109776 106276
rect 109828 106264 109834 106276
rect 191190 106264 191196 106276
rect 109828 106236 191196 106264
rect 109828 106224 109834 106236
rect 191190 106224 191196 106236
rect 191248 106224 191254 106276
rect 46842 105544 46848 105596
rect 46900 105584 46906 105596
rect 65886 105584 65892 105596
rect 46900 105556 65892 105584
rect 46900 105544 46906 105556
rect 65886 105544 65892 105556
rect 65944 105584 65950 105596
rect 66530 105584 66536 105596
rect 65944 105556 66536 105584
rect 65944 105544 65950 105556
rect 66530 105544 66536 105556
rect 66588 105544 66594 105596
rect 158070 105544 158076 105596
rect 158128 105584 158134 105596
rect 190270 105584 190276 105596
rect 158128 105556 190276 105584
rect 158128 105544 158134 105556
rect 190270 105544 190276 105556
rect 190328 105584 190334 105596
rect 191742 105584 191748 105596
rect 190328 105556 191748 105584
rect 190328 105544 190334 105556
rect 191742 105544 191748 105556
rect 191800 105544 191806 105596
rect 226702 105544 226708 105596
rect 226760 105584 226766 105596
rect 266998 105584 267004 105596
rect 226760 105556 267004 105584
rect 226760 105544 226766 105556
rect 266998 105544 267004 105556
rect 267056 105544 267062 105596
rect 112438 105340 112444 105392
rect 112496 105380 112502 105392
rect 113266 105380 113272 105392
rect 112496 105352 113272 105380
rect 112496 105340 112502 105352
rect 113266 105340 113272 105352
rect 113324 105340 113330 105392
rect 53466 104796 53472 104848
rect 53524 104836 53530 104848
rect 66806 104836 66812 104848
rect 53524 104808 66812 104836
rect 53524 104796 53530 104808
rect 66806 104796 66812 104808
rect 66864 104796 66870 104848
rect 96798 104116 96804 104168
rect 96856 104156 96862 104168
rect 112438 104156 112444 104168
rect 96856 104128 112444 104156
rect 96856 104116 96862 104128
rect 112438 104116 112444 104128
rect 112496 104116 112502 104168
rect 130470 104116 130476 104168
rect 130528 104156 130534 104168
rect 152550 104156 152556 104168
rect 130528 104128 152556 104156
rect 130528 104116 130534 104128
rect 152550 104116 152556 104128
rect 152608 104116 152614 104168
rect 233326 104116 233332 104168
rect 233384 104156 233390 104168
rect 235902 104156 235908 104168
rect 233384 104128 235908 104156
rect 233384 104116 233390 104128
rect 235902 104116 235908 104128
rect 235960 104156 235966 104168
rect 305638 104156 305644 104168
rect 235960 104128 305644 104156
rect 235960 104116 235966 104128
rect 305638 104116 305644 104128
rect 305696 104116 305702 104168
rect 96522 103504 96528 103556
rect 96580 103544 96586 103556
rect 183002 103544 183008 103556
rect 96580 103516 183008 103544
rect 96580 103504 96586 103516
rect 183002 103504 183008 103516
rect 183060 103504 183066 103556
rect 226702 103504 226708 103556
rect 226760 103544 226766 103556
rect 233326 103544 233332 103556
rect 226760 103516 233332 103544
rect 226760 103504 226766 103516
rect 233326 103504 233332 103516
rect 233384 103504 233390 103556
rect 63218 103436 63224 103488
rect 63276 103476 63282 103488
rect 66806 103476 66812 103488
rect 63276 103448 66812 103476
rect 63276 103436 63282 103448
rect 66806 103436 66812 103448
rect 66864 103436 66870 103488
rect 164142 103436 164148 103488
rect 164200 103476 164206 103488
rect 193030 103476 193036 103488
rect 164200 103448 193036 103476
rect 164200 103436 164206 103448
rect 193030 103436 193036 103448
rect 193088 103436 193094 103488
rect 97994 102824 98000 102876
rect 98052 102864 98058 102876
rect 166350 102864 166356 102876
rect 98052 102836 166356 102864
rect 98052 102824 98058 102836
rect 166350 102824 166356 102836
rect 166408 102824 166414 102876
rect 94590 102756 94596 102808
rect 94648 102796 94654 102808
rect 164142 102796 164148 102808
rect 94648 102768 164148 102796
rect 94648 102756 94654 102768
rect 164142 102756 164148 102768
rect 164200 102756 164206 102808
rect 233142 102756 233148 102808
rect 233200 102796 233206 102808
rect 278774 102796 278780 102808
rect 233200 102768 278780 102796
rect 233200 102756 233206 102768
rect 278774 102756 278780 102768
rect 278832 102796 278838 102808
rect 321646 102796 321652 102808
rect 278832 102768 321652 102796
rect 278832 102756 278838 102768
rect 321646 102756 321652 102768
rect 321704 102756 321710 102808
rect 182910 102212 182916 102264
rect 182968 102252 182974 102264
rect 191742 102252 191748 102264
rect 182968 102224 191748 102252
rect 182968 102212 182974 102224
rect 191742 102212 191748 102224
rect 191800 102212 191806 102264
rect 226610 102212 226616 102264
rect 226668 102252 226674 102264
rect 231854 102252 231860 102264
rect 226668 102224 231860 102252
rect 226668 102212 226674 102224
rect 231854 102212 231860 102224
rect 231912 102252 231918 102264
rect 233142 102252 233148 102264
rect 231912 102224 233148 102252
rect 231912 102212 231918 102224
rect 233142 102212 233148 102224
rect 233200 102212 233206 102264
rect 226702 102144 226708 102196
rect 226760 102184 226766 102196
rect 237558 102184 237564 102196
rect 226760 102156 237564 102184
rect 226760 102144 226766 102156
rect 237558 102144 237564 102156
rect 237616 102144 237622 102196
rect 97902 102076 97908 102128
rect 97960 102116 97966 102128
rect 129090 102116 129096 102128
rect 97960 102088 129096 102116
rect 97960 102076 97966 102088
rect 129090 102076 129096 102088
rect 129148 102076 129154 102128
rect 226518 102076 226524 102128
rect 226576 102116 226582 102128
rect 266354 102116 266360 102128
rect 226576 102088 266360 102116
rect 226576 102076 226582 102088
rect 266354 102076 266360 102088
rect 266412 102076 266418 102128
rect 129090 101464 129096 101516
rect 129148 101504 129154 101516
rect 162210 101504 162216 101516
rect 129148 101476 162216 101504
rect 129148 101464 129154 101476
rect 162210 101464 162216 101476
rect 162268 101464 162274 101516
rect 55122 101396 55128 101448
rect 55180 101436 55186 101448
rect 66070 101436 66076 101448
rect 55180 101408 66076 101436
rect 55180 101396 55186 101408
rect 66070 101396 66076 101408
rect 66128 101436 66134 101448
rect 66622 101436 66628 101448
rect 66128 101408 66628 101436
rect 66128 101396 66134 101408
rect 66622 101396 66628 101408
rect 66680 101396 66686 101448
rect 98822 101396 98828 101448
rect 98880 101436 98886 101448
rect 162762 101436 162768 101448
rect 98880 101408 162768 101436
rect 98880 101396 98886 101408
rect 162762 101396 162768 101408
rect 162820 101436 162826 101448
rect 191466 101436 191472 101448
rect 162820 101408 191472 101436
rect 162820 101396 162826 101408
rect 191466 101396 191472 101408
rect 191524 101436 191530 101448
rect 191742 101436 191748 101448
rect 191524 101408 191748 101436
rect 191524 101396 191530 101408
rect 191742 101396 191748 101408
rect 191800 101396 191806 101448
rect 186222 100648 186228 100700
rect 186280 100688 186286 100700
rect 191742 100688 191748 100700
rect 186280 100660 191748 100688
rect 186280 100648 186286 100660
rect 191742 100648 191748 100660
rect 191800 100648 191806 100700
rect 178862 100036 178868 100088
rect 178920 100076 178926 100088
rect 191098 100076 191104 100088
rect 178920 100048 191104 100076
rect 178920 100036 178926 100048
rect 191098 100036 191104 100048
rect 191156 100036 191162 100088
rect 57882 99968 57888 100020
rect 57940 100008 57946 100020
rect 64690 100008 64696 100020
rect 57940 99980 64696 100008
rect 57940 99968 57946 99980
rect 64690 99968 64696 99980
rect 64748 100008 64754 100020
rect 66806 100008 66812 100020
rect 64748 99980 66812 100008
rect 64748 99968 64754 99980
rect 66806 99968 66812 99980
rect 66864 99968 66870 100020
rect 97902 99968 97908 100020
rect 97960 100008 97966 100020
rect 101398 100008 101404 100020
rect 97960 99980 101404 100008
rect 97960 99968 97966 99980
rect 101398 99968 101404 99980
rect 101456 100008 101462 100020
rect 184290 100008 184296 100020
rect 101456 99980 184296 100008
rect 101456 99968 101462 99980
rect 184290 99968 184296 99980
rect 184348 99968 184354 100020
rect 226702 99424 226708 99476
rect 226760 99464 226766 99476
rect 229186 99464 229192 99476
rect 226760 99436 229192 99464
rect 226760 99424 226766 99436
rect 229186 99424 229192 99436
rect 229244 99464 229250 99476
rect 245654 99464 245660 99476
rect 229244 99436 245660 99464
rect 229244 99424 229250 99436
rect 245654 99424 245660 99436
rect 245712 99424 245718 99476
rect 97534 99356 97540 99408
rect 97592 99396 97598 99408
rect 133782 99396 133788 99408
rect 97592 99368 133788 99396
rect 97592 99356 97598 99368
rect 133782 99356 133788 99368
rect 133840 99356 133846 99408
rect 226610 99356 226616 99408
rect 226668 99396 226674 99408
rect 320818 99396 320824 99408
rect 226668 99368 320824 99396
rect 226668 99356 226674 99368
rect 320818 99356 320824 99368
rect 320876 99356 320882 99408
rect 60550 99288 60556 99340
rect 60608 99328 60614 99340
rect 66806 99328 66812 99340
rect 60608 99300 66812 99328
rect 60608 99288 60614 99300
rect 66806 99288 66812 99300
rect 66864 99288 66870 99340
rect 227346 98608 227352 98660
rect 227404 98648 227410 98660
rect 236638 98648 236644 98660
rect 227404 98620 236644 98648
rect 227404 98608 227410 98620
rect 236638 98608 236644 98620
rect 236696 98608 236702 98660
rect 245654 98608 245660 98660
rect 245712 98648 245718 98660
rect 277394 98648 277400 98660
rect 245712 98620 277400 98648
rect 245712 98608 245718 98620
rect 277394 98608 277400 98620
rect 277452 98608 277458 98660
rect 97810 98064 97816 98116
rect 97868 98104 97874 98116
rect 106274 98104 106280 98116
rect 97868 98076 106280 98104
rect 97868 98064 97874 98076
rect 106274 98064 106280 98076
rect 106332 98064 106338 98116
rect 97902 97996 97908 98048
rect 97960 98036 97966 98048
rect 152550 98036 152556 98048
rect 97960 98008 152556 98036
rect 97960 97996 97966 98008
rect 152550 97996 152556 98008
rect 152608 97996 152614 98048
rect 187510 97996 187516 98048
rect 187568 98036 187574 98048
rect 190546 98036 190552 98048
rect 187568 98008 190552 98036
rect 187568 97996 187574 98008
rect 190546 97996 190552 98008
rect 190604 97996 190610 98048
rect 159542 97928 159548 97980
rect 159600 97968 159606 97980
rect 190454 97968 190460 97980
rect 159600 97940 190460 97968
rect 159600 97928 159606 97940
rect 190454 97928 190460 97940
rect 190512 97928 190518 97980
rect 226242 97928 226248 97980
rect 226300 97968 226306 97980
rect 237650 97968 237656 97980
rect 226300 97940 237656 97968
rect 226300 97928 226306 97940
rect 237650 97928 237656 97940
rect 237708 97928 237714 97980
rect 96706 97724 96712 97776
rect 96764 97764 96770 97776
rect 98638 97764 98644 97776
rect 96764 97736 98644 97764
rect 96764 97724 96770 97736
rect 98638 97724 98644 97736
rect 98696 97724 98702 97776
rect 97810 97248 97816 97300
rect 97868 97288 97874 97300
rect 129734 97288 129740 97300
rect 97868 97260 129740 97288
rect 97868 97248 97874 97260
rect 129734 97248 129740 97260
rect 129792 97248 129798 97300
rect 3418 96636 3424 96688
rect 3476 96676 3482 96688
rect 61378 96676 61384 96688
rect 3476 96648 61384 96676
rect 3476 96636 3482 96648
rect 61378 96636 61384 96648
rect 61436 96636 61442 96688
rect 226702 96568 226708 96620
rect 226760 96608 226766 96620
rect 262306 96608 262312 96620
rect 226760 96580 262312 96608
rect 226760 96568 226766 96580
rect 262306 96568 262312 96580
rect 262364 96568 262370 96620
rect 59078 95888 59084 95940
rect 59136 95928 59142 95940
rect 66438 95928 66444 95940
rect 59136 95900 66444 95928
rect 59136 95888 59142 95900
rect 66438 95888 66444 95900
rect 66496 95888 66502 95940
rect 226886 95888 226892 95940
rect 226944 95928 226950 95940
rect 273346 95928 273352 95940
rect 226944 95900 273352 95928
rect 226944 95888 226950 95900
rect 273346 95888 273352 95900
rect 273404 95888 273410 95940
rect 97074 95276 97080 95328
rect 97132 95316 97138 95328
rect 100018 95316 100024 95328
rect 97132 95288 100024 95316
rect 97132 95276 97138 95288
rect 100018 95276 100024 95288
rect 100076 95276 100082 95328
rect 97902 95208 97908 95260
rect 97960 95248 97966 95260
rect 188338 95248 188344 95260
rect 97960 95220 188344 95248
rect 97960 95208 97966 95220
rect 188338 95208 188344 95220
rect 188396 95208 188402 95260
rect 61838 95140 61844 95192
rect 61896 95180 61902 95192
rect 66806 95180 66812 95192
rect 61896 95152 66812 95180
rect 61896 95140 61902 95152
rect 66806 95140 66812 95152
rect 66864 95140 66870 95192
rect 67542 95140 67548 95192
rect 67600 95180 67606 95192
rect 68278 95180 68284 95192
rect 67600 95152 68284 95180
rect 67600 95140 67606 95152
rect 68278 95140 68284 95152
rect 68336 95140 68342 95192
rect 99006 94528 99012 94580
rect 99064 94568 99070 94580
rect 166442 94568 166448 94580
rect 99064 94540 166448 94568
rect 99064 94528 99070 94540
rect 166442 94528 166448 94540
rect 166500 94528 166506 94580
rect 191466 94528 191472 94580
rect 191524 94568 191530 94580
rect 191742 94568 191748 94580
rect 191524 94540 191748 94568
rect 191524 94528 191530 94540
rect 191742 94528 191748 94540
rect 191800 94528 191806 94580
rect 95510 94460 95516 94512
rect 95568 94500 95574 94512
rect 177942 94500 177948 94512
rect 95568 94472 177948 94500
rect 95568 94460 95574 94472
rect 177942 94460 177948 94472
rect 178000 94500 178006 94512
rect 191834 94500 191840 94512
rect 178000 94472 191840 94500
rect 178000 94460 178006 94472
rect 191834 94460 191840 94472
rect 191892 94460 191898 94512
rect 170490 93848 170496 93900
rect 170548 93888 170554 93900
rect 193398 93888 193404 93900
rect 170548 93860 193404 93888
rect 170548 93848 170554 93860
rect 193398 93848 193404 93860
rect 193456 93848 193462 93900
rect 67542 93780 67548 93832
rect 67600 93820 67606 93832
rect 67910 93820 67916 93832
rect 67600 93792 67916 93820
rect 67600 93780 67606 93792
rect 67910 93780 67916 93792
rect 67968 93780 67974 93832
rect 97902 93780 97908 93832
rect 97960 93820 97966 93832
rect 106366 93820 106372 93832
rect 97960 93792 106372 93820
rect 97960 93780 97966 93792
rect 106366 93780 106372 93792
rect 106424 93780 106430 93832
rect 186958 93780 186964 93832
rect 187016 93820 187022 93832
rect 193214 93820 193220 93832
rect 187016 93792 193220 93820
rect 187016 93780 187022 93792
rect 193214 93780 193220 93792
rect 193272 93780 193278 93832
rect 191834 93372 191840 93424
rect 191892 93412 191898 93424
rect 199102 93412 199108 93424
rect 191892 93384 199108 93412
rect 191892 93372 191898 93384
rect 199102 93372 199108 93384
rect 199160 93372 199166 93424
rect 221642 93372 221648 93424
rect 221700 93412 221706 93424
rect 225138 93412 225144 93424
rect 221700 93384 225144 93412
rect 221700 93372 221706 93384
rect 225138 93372 225144 93384
rect 225196 93372 225202 93424
rect 193398 93304 193404 93356
rect 193456 93344 193462 93356
rect 193766 93344 193772 93356
rect 193456 93316 193772 93344
rect 193456 93304 193462 93316
rect 193766 93304 193772 93316
rect 193824 93304 193830 93356
rect 168282 93168 168288 93220
rect 168340 93208 168346 93220
rect 183554 93208 183560 93220
rect 168340 93180 183560 93208
rect 168340 93168 168346 93180
rect 183554 93168 183560 93180
rect 183612 93208 183618 93220
rect 190454 93208 190460 93220
rect 183612 93180 190460 93208
rect 183612 93168 183618 93180
rect 190454 93168 190460 93180
rect 190512 93168 190518 93220
rect 249150 93168 249156 93220
rect 249208 93208 249214 93220
rect 264974 93208 264980 93220
rect 249208 93180 264980 93208
rect 249208 93168 249214 93180
rect 264974 93168 264980 93180
rect 265032 93168 265038 93220
rect 107470 93100 107476 93152
rect 107528 93140 107534 93152
rect 170490 93140 170496 93152
rect 107528 93112 170496 93140
rect 107528 93100 107534 93112
rect 170490 93100 170496 93112
rect 170548 93100 170554 93152
rect 207658 93100 207664 93152
rect 207716 93140 207722 93152
rect 225046 93140 225052 93152
rect 207716 93112 225052 93140
rect 207716 93100 207722 93112
rect 225046 93100 225052 93112
rect 225104 93100 225110 93152
rect 258810 93100 258816 93152
rect 258868 93140 258874 93152
rect 316034 93140 316040 93152
rect 258868 93112 316040 93140
rect 258868 93100 258874 93112
rect 316034 93100 316040 93112
rect 316092 93100 316098 93152
rect 67634 92828 67640 92880
rect 67692 92868 67698 92880
rect 68462 92868 68468 92880
rect 67692 92840 68468 92868
rect 67692 92828 67698 92840
rect 68462 92828 68468 92840
rect 68520 92828 68526 92880
rect 95234 92800 95240 92812
rect 87570 92772 95240 92800
rect 87570 92744 87598 92772
rect 95234 92760 95240 92772
rect 95292 92760 95298 92812
rect 71728 92692 71734 92744
rect 71786 92692 71792 92744
rect 87552 92692 87558 92744
rect 87610 92692 87616 92744
rect 93808 92692 93814 92744
rect 93866 92732 93872 92744
rect 94682 92732 94688 92744
rect 93866 92704 94688 92732
rect 93866 92692 93872 92704
rect 94682 92692 94688 92704
rect 94740 92692 94746 92744
rect 71746 92608 71774 92692
rect 59262 92556 59268 92608
rect 59320 92596 59326 92608
rect 66990 92596 66996 92608
rect 59320 92568 66996 92596
rect 59320 92556 59326 92568
rect 66990 92556 66996 92568
rect 67048 92596 67054 92608
rect 67266 92596 67272 92608
rect 67048 92568 67272 92596
rect 67048 92556 67054 92568
rect 67266 92556 67272 92568
rect 67324 92556 67330 92608
rect 71746 92568 71780 92608
rect 71774 92556 71780 92568
rect 71832 92556 71838 92608
rect 74534 92556 74540 92608
rect 74592 92596 74598 92608
rect 75776 92596 75782 92608
rect 74592 92568 75782 92596
rect 74592 92556 74598 92568
rect 75776 92556 75782 92568
rect 75834 92556 75840 92608
rect 81618 92556 81624 92608
rect 81676 92596 81682 92608
rect 82584 92596 82590 92608
rect 81676 92568 82590 92596
rect 81676 92556 81682 92568
rect 82584 92556 82590 92568
rect 82642 92556 82648 92608
rect 86954 92556 86960 92608
rect 87012 92596 87018 92608
rect 88104 92596 88110 92608
rect 87012 92568 88110 92596
rect 87012 92556 87018 92568
rect 88104 92556 88110 92568
rect 88162 92556 88168 92608
rect 89898 92556 89904 92608
rect 89956 92596 89962 92608
rect 90680 92596 90686 92608
rect 89956 92568 90686 92596
rect 89956 92556 89962 92568
rect 90680 92556 90686 92568
rect 90738 92556 90744 92608
rect 94498 92488 94504 92540
rect 94556 92528 94562 92540
rect 122834 92528 122840 92540
rect 94556 92500 122840 92528
rect 94556 92488 94562 92500
rect 122834 92488 122840 92500
rect 122892 92488 122898 92540
rect 56502 92420 56508 92472
rect 56560 92460 56566 92472
rect 72786 92460 72792 92472
rect 56560 92432 72792 92460
rect 56560 92420 56566 92432
rect 72786 92420 72792 92432
rect 72844 92420 72850 92472
rect 75454 92420 75460 92472
rect 75512 92460 75518 92472
rect 95878 92460 95884 92472
rect 75512 92432 95884 92460
rect 75512 92420 75518 92432
rect 95878 92420 95884 92432
rect 95936 92420 95942 92472
rect 184290 92420 184296 92472
rect 184348 92460 184354 92472
rect 226610 92460 226616 92472
rect 184348 92432 226616 92460
rect 184348 92420 184354 92432
rect 226610 92420 226616 92432
rect 226668 92420 226674 92472
rect 60642 92352 60648 92404
rect 60700 92392 60706 92404
rect 81434 92392 81440 92404
rect 60700 92364 81440 92392
rect 60700 92352 60706 92364
rect 81434 92352 81440 92364
rect 81492 92352 81498 92404
rect 92382 92352 92388 92404
rect 92440 92392 92446 92404
rect 103514 92392 103520 92404
rect 92440 92364 103520 92392
rect 92440 92352 92446 92364
rect 103514 92352 103520 92364
rect 103572 92352 103578 92404
rect 205634 92352 205640 92404
rect 205692 92392 205698 92404
rect 225230 92392 225236 92404
rect 205692 92364 225236 92392
rect 205692 92352 205698 92364
rect 225230 92352 225236 92364
rect 225288 92352 225294 92404
rect 193214 92080 193220 92132
rect 193272 92120 193278 92132
rect 193766 92120 193772 92132
rect 193272 92092 193772 92120
rect 193272 92080 193278 92092
rect 193766 92080 193772 92092
rect 193824 92080 193830 92132
rect 112438 91740 112444 91792
rect 112496 91780 112502 91792
rect 205634 91780 205640 91792
rect 112496 91752 205640 91780
rect 112496 91740 112502 91752
rect 205634 91740 205640 91752
rect 205692 91740 205698 91792
rect 245010 91740 245016 91792
rect 245068 91780 245074 91792
rect 258718 91780 258724 91792
rect 245068 91752 258724 91780
rect 245068 91740 245074 91752
rect 258718 91740 258724 91752
rect 258776 91740 258782 91792
rect 104342 91060 104348 91112
rect 104400 91100 104406 91112
rect 111058 91100 111064 91112
rect 104400 91072 111064 91100
rect 104400 91060 104406 91072
rect 111058 91060 111064 91072
rect 111116 91060 111122 91112
rect 63402 90992 63408 91044
rect 63460 91032 63466 91044
rect 73706 91032 73712 91044
rect 63460 91004 73712 91032
rect 63460 90992 63466 91004
rect 73706 90992 73712 91004
rect 73764 90992 73770 91044
rect 112438 90992 112444 91044
rect 112496 91032 112502 91044
rect 113174 91032 113180 91044
rect 112496 91004 113180 91032
rect 112496 90992 112502 91004
rect 113174 90992 113180 91004
rect 113232 90992 113238 91044
rect 179322 90992 179328 91044
rect 179380 91032 179386 91044
rect 194686 91032 194692 91044
rect 179380 91004 194692 91032
rect 179380 90992 179386 91004
rect 194686 90992 194692 91004
rect 194744 91032 194750 91044
rect 195238 91032 195244 91044
rect 194744 91004 195244 91032
rect 194744 90992 194750 91004
rect 195238 90992 195244 91004
rect 195296 90992 195302 91044
rect 217318 90992 217324 91044
rect 217376 91032 217382 91044
rect 296714 91032 296720 91044
rect 217376 91004 296720 91032
rect 217376 90992 217382 91004
rect 296714 90992 296720 91004
rect 296772 90992 296778 91044
rect 66162 90924 66168 90976
rect 66220 90964 66226 90976
rect 70302 90964 70308 90976
rect 66220 90936 70308 90964
rect 66220 90924 66226 90936
rect 70302 90924 70308 90936
rect 70360 90924 70366 90976
rect 78950 90312 78956 90364
rect 79008 90352 79014 90364
rect 96706 90352 96712 90364
rect 79008 90324 96712 90352
rect 79008 90312 79014 90324
rect 96706 90312 96712 90324
rect 96764 90352 96770 90364
rect 97258 90352 97264 90364
rect 96764 90324 97264 90352
rect 96764 90312 96770 90324
rect 97258 90312 97264 90324
rect 97316 90312 97322 90364
rect 105538 90312 105544 90364
rect 105596 90352 105602 90364
rect 212902 90352 212908 90364
rect 105596 90324 212908 90352
rect 105596 90312 105602 90324
rect 212902 90312 212908 90324
rect 212960 90312 212966 90364
rect 242158 90312 242164 90364
rect 242216 90352 242222 90364
rect 271138 90352 271144 90364
rect 242216 90324 271144 90352
rect 242216 90312 242222 90324
rect 271138 90312 271144 90324
rect 271196 90312 271202 90364
rect 70302 90244 70308 90296
rect 70360 90284 70366 90296
rect 71038 90284 71044 90296
rect 70360 90256 71044 90284
rect 70360 90244 70366 90256
rect 71038 90244 71044 90256
rect 71096 90244 71102 90296
rect 223758 90244 223764 90296
rect 223816 90284 223822 90296
rect 224862 90284 224868 90296
rect 223816 90256 224868 90284
rect 223816 90244 223822 90256
rect 224862 90244 224868 90256
rect 224920 90244 224926 90296
rect 204346 89768 204352 89820
rect 204404 89808 204410 89820
rect 205542 89808 205548 89820
rect 204404 89780 205548 89808
rect 204404 89768 204410 89780
rect 205542 89768 205548 89780
rect 205600 89768 205606 89820
rect 124858 89700 124864 89752
rect 124916 89740 124922 89752
rect 125594 89740 125600 89752
rect 124916 89712 125600 89740
rect 124916 89700 124922 89712
rect 125594 89700 125600 89712
rect 125652 89700 125658 89752
rect 204898 89700 204904 89752
rect 204956 89740 204962 89752
rect 207934 89740 207940 89752
rect 204956 89712 207940 89740
rect 204956 89700 204962 89712
rect 207934 89700 207940 89712
rect 207992 89700 207998 89752
rect 67542 89632 67548 89684
rect 67600 89672 67606 89684
rect 99006 89672 99012 89684
rect 67600 89644 99012 89672
rect 67600 89632 67606 89644
rect 99006 89632 99012 89644
rect 99064 89632 99070 89684
rect 217686 89672 217692 89684
rect 122806 89644 217692 89672
rect 61654 89564 61660 89616
rect 61712 89604 61718 89616
rect 74810 89604 74816 89616
rect 61712 89576 74816 89604
rect 61712 89564 61718 89576
rect 74810 89564 74816 89576
rect 74868 89564 74874 89616
rect 89254 89564 89260 89616
rect 89312 89604 89318 89616
rect 118694 89604 118700 89616
rect 89312 89576 118700 89604
rect 89312 89564 89318 89576
rect 118694 89564 118700 89576
rect 118752 89604 118758 89616
rect 122806 89604 122834 89644
rect 217686 89632 217692 89644
rect 217744 89632 217750 89684
rect 219986 89632 219992 89684
rect 220044 89672 220050 89684
rect 277486 89672 277492 89684
rect 220044 89644 277492 89672
rect 220044 89632 220050 89644
rect 277486 89632 277492 89644
rect 277544 89672 277550 89684
rect 278682 89672 278688 89684
rect 277544 89644 278688 89672
rect 277544 89632 277550 89644
rect 278682 89632 278688 89644
rect 278740 89632 278746 89684
rect 118752 89576 122834 89604
rect 118752 89564 118758 89576
rect 125410 89564 125416 89616
rect 125468 89604 125474 89616
rect 218238 89604 218244 89616
rect 125468 89576 218244 89604
rect 125468 89564 125474 89576
rect 218238 89564 218244 89576
rect 218296 89564 218302 89616
rect 278682 88952 278688 89004
rect 278740 88992 278746 89004
rect 582374 88992 582380 89004
rect 278740 88964 582380 88992
rect 278740 88952 278746 88964
rect 582374 88952 582380 88964
rect 582432 88952 582438 89004
rect 52270 88272 52276 88324
rect 52328 88312 52334 88324
rect 79410 88312 79416 88324
rect 52328 88284 79416 88312
rect 52328 88272 52334 88284
rect 79410 88272 79416 88284
rect 79468 88272 79474 88324
rect 87598 88272 87604 88324
rect 87656 88312 87662 88324
rect 88150 88312 88156 88324
rect 87656 88284 88156 88312
rect 87656 88272 87662 88284
rect 88150 88272 88156 88284
rect 88208 88272 88214 88324
rect 121454 88272 121460 88324
rect 121512 88312 121518 88324
rect 215386 88312 215392 88324
rect 121512 88284 215392 88312
rect 121512 88272 121518 88284
rect 215386 88272 215392 88284
rect 215444 88272 215450 88324
rect 73706 88204 73712 88256
rect 73764 88244 73770 88256
rect 95510 88244 95516 88256
rect 73764 88216 95516 88244
rect 73764 88204 73770 88216
rect 95510 88204 95516 88216
rect 95568 88204 95574 88256
rect 205634 88204 205640 88256
rect 205692 88244 205698 88256
rect 226426 88244 226432 88256
rect 205692 88216 226432 88244
rect 205692 88204 205698 88216
rect 226426 88204 226432 88216
rect 226484 88204 226490 88256
rect 100110 87592 100116 87644
rect 100168 87632 100174 87644
rect 125410 87632 125416 87644
rect 100168 87604 125416 87632
rect 100168 87592 100174 87604
rect 125410 87592 125416 87604
rect 125468 87592 125474 87644
rect 164970 87592 164976 87644
rect 165028 87632 165034 87644
rect 165522 87632 165528 87644
rect 165028 87604 165528 87632
rect 165028 87592 165034 87604
rect 165522 87592 165528 87604
rect 165580 87632 165586 87644
rect 206830 87632 206836 87644
rect 165580 87604 206836 87632
rect 165580 87592 165586 87604
rect 206830 87592 206836 87604
rect 206888 87592 206894 87644
rect 227530 87592 227536 87644
rect 227588 87632 227594 87644
rect 241514 87632 241520 87644
rect 227588 87604 241520 87632
rect 227588 87592 227594 87604
rect 241514 87592 241520 87604
rect 241572 87592 241578 87644
rect 80054 86912 80060 86964
rect 80112 86952 80118 86964
rect 165522 86952 165528 86964
rect 80112 86924 165528 86952
rect 80112 86912 80118 86924
rect 165522 86912 165528 86924
rect 165580 86912 165586 86964
rect 184658 86912 184664 86964
rect 184716 86952 184722 86964
rect 199378 86952 199384 86964
rect 184716 86924 199384 86952
rect 184716 86912 184722 86924
rect 199378 86912 199384 86924
rect 199436 86912 199442 86964
rect 212902 86912 212908 86964
rect 212960 86952 212966 86964
rect 213822 86952 213828 86964
rect 212960 86924 213828 86952
rect 212960 86912 212966 86924
rect 213822 86912 213828 86924
rect 213880 86952 213886 86964
rect 235258 86952 235264 86964
rect 213880 86924 235264 86952
rect 213880 86912 213886 86924
rect 235258 86912 235264 86924
rect 235316 86912 235322 86964
rect 259362 86912 259368 86964
rect 259420 86952 259426 86964
rect 276658 86952 276664 86964
rect 259420 86924 276664 86952
rect 259420 86912 259426 86924
rect 276658 86912 276664 86924
rect 276716 86952 276722 86964
rect 580166 86952 580172 86964
rect 276716 86924 580172 86952
rect 276716 86912 276722 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 67358 86844 67364 86896
rect 67416 86884 67422 86896
rect 98822 86884 98828 86896
rect 67416 86856 98828 86884
rect 67416 86844 67422 86856
rect 98822 86844 98828 86856
rect 98880 86844 98886 86896
rect 199470 86232 199476 86284
rect 199528 86272 199534 86284
rect 244274 86272 244280 86284
rect 199528 86244 244280 86272
rect 199528 86232 199534 86244
rect 244274 86232 244280 86244
rect 244332 86232 244338 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 57238 85524 57244 85536
rect 3200 85496 57244 85524
rect 3200 85484 3206 85496
rect 57238 85484 57244 85496
rect 57296 85524 57302 85536
rect 160830 85524 160836 85536
rect 57296 85496 160836 85524
rect 57296 85484 57302 85496
rect 160830 85484 160836 85496
rect 160888 85484 160894 85536
rect 220630 85484 220636 85536
rect 220688 85524 220694 85536
rect 263686 85524 263692 85536
rect 220688 85496 263692 85524
rect 220688 85484 220694 85496
rect 263686 85484 263692 85496
rect 263744 85484 263750 85536
rect 69198 85416 69204 85468
rect 69256 85456 69262 85468
rect 107470 85456 107476 85468
rect 69256 85428 107476 85456
rect 69256 85416 69262 85428
rect 107470 85416 107476 85428
rect 107528 85416 107534 85468
rect 108114 85416 108120 85468
rect 108172 85456 108178 85468
rect 204990 85456 204996 85468
rect 108172 85428 204996 85456
rect 108172 85416 108178 85428
rect 204990 85416 204996 85428
rect 205048 85416 205054 85468
rect 242802 85416 242808 85468
rect 242860 85456 242866 85468
rect 243538 85456 243544 85468
rect 242860 85428 243544 85456
rect 242860 85416 242866 85428
rect 243538 85416 243544 85428
rect 243596 85416 243602 85468
rect 206830 84804 206836 84856
rect 206888 84844 206894 84856
rect 220078 84844 220084 84856
rect 206888 84816 220084 84844
rect 206888 84804 206894 84816
rect 220078 84804 220084 84816
rect 220136 84804 220142 84856
rect 216030 84192 216036 84244
rect 216088 84232 216094 84244
rect 242802 84232 242808 84244
rect 216088 84204 242808 84232
rect 216088 84192 216094 84204
rect 242802 84192 242808 84204
rect 242860 84192 242866 84244
rect 67818 84124 67824 84176
rect 67876 84164 67882 84176
rect 94590 84164 94596 84176
rect 67876 84136 94596 84164
rect 67876 84124 67882 84136
rect 94590 84124 94596 84136
rect 94648 84124 94654 84176
rect 104158 84124 104164 84176
rect 104216 84164 104222 84176
rect 213914 84164 213920 84176
rect 104216 84136 213920 84164
rect 104216 84124 104222 84136
rect 213914 84124 213920 84136
rect 213972 84124 213978 84176
rect 70394 84056 70400 84108
rect 70452 84096 70458 84108
rect 169662 84096 169668 84108
rect 70452 84068 169668 84096
rect 70452 84056 70458 84068
rect 169662 84056 169668 84068
rect 169720 84096 169726 84108
rect 195974 84096 195980 84108
rect 169720 84068 195980 84096
rect 169720 84056 169726 84068
rect 195974 84056 195980 84068
rect 196032 84056 196038 84108
rect 209866 84056 209872 84108
rect 209924 84096 209930 84108
rect 210418 84096 210424 84108
rect 209924 84068 210424 84096
rect 209924 84056 209930 84068
rect 210418 84056 210424 84068
rect 210476 84096 210482 84108
rect 275002 84096 275008 84108
rect 210476 84068 275008 84096
rect 210476 84056 210482 84068
rect 275002 84056 275008 84068
rect 275060 84056 275066 84108
rect 275002 83444 275008 83496
rect 275060 83484 275066 83496
rect 322934 83484 322940 83496
rect 275060 83456 322940 83484
rect 275060 83444 275066 83456
rect 322934 83444 322940 83456
rect 322992 83444 322998 83496
rect 195974 82832 195980 82884
rect 196032 82872 196038 82884
rect 196618 82872 196624 82884
rect 196032 82844 196624 82872
rect 196032 82832 196038 82844
rect 196618 82832 196624 82844
rect 196676 82832 196682 82884
rect 75914 82764 75920 82816
rect 75972 82804 75978 82816
rect 102778 82804 102784 82816
rect 75972 82776 102784 82804
rect 75972 82764 75978 82776
rect 102778 82764 102784 82776
rect 102836 82764 102842 82816
rect 115290 82764 115296 82816
rect 115348 82804 115354 82816
rect 224954 82804 224960 82816
rect 115348 82776 224960 82804
rect 115348 82764 115354 82776
rect 224954 82764 224960 82776
rect 225012 82764 225018 82816
rect 84194 82696 84200 82748
rect 84252 82736 84258 82748
rect 105538 82736 105544 82748
rect 84252 82708 105544 82736
rect 84252 82696 84258 82708
rect 105538 82696 105544 82708
rect 105596 82696 105602 82748
rect 155402 82696 155408 82748
rect 155460 82736 155466 82748
rect 252738 82736 252744 82748
rect 155460 82708 252744 82736
rect 155460 82696 155466 82708
rect 252738 82696 252744 82708
rect 252796 82696 252802 82748
rect 252738 81404 252744 81456
rect 252796 81444 252802 81456
rect 253198 81444 253204 81456
rect 252796 81416 253204 81444
rect 252796 81404 252802 81416
rect 253198 81404 253204 81416
rect 253256 81404 253262 81456
rect 80146 81336 80152 81388
rect 80204 81376 80210 81388
rect 112438 81376 112444 81388
rect 80204 81348 112444 81376
rect 80204 81336 80210 81348
rect 112438 81336 112444 81348
rect 112496 81336 112502 81388
rect 183002 81336 183008 81388
rect 183060 81376 183066 81388
rect 233326 81376 233332 81388
rect 183060 81348 233332 81376
rect 183060 81336 183066 81348
rect 233326 81336 233332 81348
rect 233384 81336 233390 81388
rect 89714 81268 89720 81320
rect 89772 81308 89778 81320
rect 100110 81308 100116 81320
rect 89772 81280 100116 81308
rect 89772 81268 89778 81280
rect 100110 81268 100116 81280
rect 100168 81268 100174 81320
rect 173802 81268 173808 81320
rect 173860 81308 173866 81320
rect 204898 81308 204904 81320
rect 173860 81280 204904 81308
rect 173860 81268 173866 81280
rect 204898 81268 204904 81280
rect 204956 81268 204962 81320
rect 262122 80044 262128 80096
rect 262180 80084 262186 80096
rect 263594 80084 263600 80096
rect 262180 80056 263600 80084
rect 262180 80044 262186 80056
rect 263594 80044 263600 80056
rect 263652 80044 263658 80096
rect 81710 79976 81716 80028
rect 81768 80016 81774 80028
rect 112530 80016 112536 80028
rect 81768 79988 112536 80016
rect 81768 79976 81774 79988
rect 112530 79976 112536 79988
rect 112588 79976 112594 80028
rect 169110 79976 169116 80028
rect 169168 80016 169174 80028
rect 230474 80016 230480 80028
rect 169168 79988 230480 80016
rect 169168 79976 169174 79988
rect 230474 79976 230480 79988
rect 230532 79976 230538 80028
rect 204162 79908 204168 79960
rect 204220 79948 204226 79960
rect 237374 79948 237380 79960
rect 204220 79920 237380 79948
rect 204220 79908 204226 79920
rect 237374 79908 237380 79920
rect 237432 79908 237438 79960
rect 203518 79500 203524 79552
rect 203576 79540 203582 79552
rect 204162 79540 204168 79552
rect 203576 79512 204168 79540
rect 203576 79500 203582 79512
rect 204162 79500 204168 79512
rect 204220 79500 204226 79552
rect 90358 79296 90364 79348
rect 90416 79336 90422 79348
rect 134610 79336 134616 79348
rect 90416 79308 134616 79336
rect 90416 79296 90422 79308
rect 134610 79296 134616 79308
rect 134668 79296 134674 79348
rect 64690 78616 64696 78668
rect 64748 78656 64754 78668
rect 191558 78656 191564 78668
rect 64748 78628 191564 78656
rect 64748 78616 64754 78628
rect 191558 78616 191564 78628
rect 191616 78656 191622 78668
rect 248414 78656 248420 78668
rect 191616 78628 248420 78656
rect 191616 78616 191622 78628
rect 248414 78616 248420 78628
rect 248472 78656 248478 78668
rect 249150 78656 249156 78668
rect 248472 78628 249156 78656
rect 248472 78616 248478 78628
rect 249150 78616 249156 78628
rect 249208 78616 249214 78668
rect 82814 78548 82820 78600
rect 82872 78588 82878 78600
rect 181254 78588 181260 78600
rect 82872 78560 181260 78588
rect 82872 78548 82878 78560
rect 181254 78548 181260 78560
rect 181312 78548 181318 78600
rect 190178 77936 190184 77988
rect 190236 77976 190242 77988
rect 214650 77976 214656 77988
rect 190236 77948 214656 77976
rect 190236 77936 190242 77948
rect 214650 77936 214656 77948
rect 214708 77936 214714 77988
rect 88334 77188 88340 77240
rect 88392 77228 88398 77240
rect 121546 77228 121552 77240
rect 88392 77200 121552 77228
rect 88392 77188 88398 77200
rect 121546 77188 121552 77200
rect 121604 77188 121610 77240
rect 133782 77188 133788 77240
rect 133840 77228 133846 77240
rect 229186 77228 229192 77240
rect 133840 77200 229192 77228
rect 133840 77188 133846 77200
rect 229186 77188 229192 77200
rect 229244 77188 229250 77240
rect 3142 76508 3148 76560
rect 3200 76548 3206 76560
rect 95326 76548 95332 76560
rect 3200 76520 95332 76548
rect 3200 76508 3206 76520
rect 95326 76508 95332 76520
rect 95384 76508 95390 76560
rect 200206 76508 200212 76560
rect 200264 76548 200270 76560
rect 245654 76548 245660 76560
rect 200264 76520 245660 76548
rect 200264 76508 200270 76520
rect 245654 76508 245660 76520
rect 245712 76508 245718 76560
rect 121546 76440 121552 76492
rect 121604 76480 121610 76492
rect 122098 76480 122104 76492
rect 121604 76452 122104 76480
rect 121604 76440 121610 76452
rect 122098 76440 122104 76452
rect 122156 76440 122162 76492
rect 57790 75828 57796 75880
rect 57848 75868 57854 75880
rect 188890 75868 188896 75880
rect 57848 75840 188896 75868
rect 57848 75828 57854 75840
rect 188890 75828 188896 75840
rect 188948 75868 188954 75880
rect 263594 75868 263600 75880
rect 188948 75840 263600 75868
rect 188948 75828 188954 75840
rect 263594 75828 263600 75840
rect 263652 75828 263658 75880
rect 65610 75760 65616 75812
rect 65668 75800 65674 75812
rect 66070 75800 66076 75812
rect 65668 75772 66076 75800
rect 65668 75760 65674 75772
rect 66070 75760 66076 75772
rect 66128 75800 66134 75812
rect 182910 75800 182916 75812
rect 66128 75772 182916 75800
rect 66128 75760 66134 75772
rect 182910 75760 182916 75772
rect 182968 75760 182974 75812
rect 81618 74468 81624 74520
rect 81676 74508 81682 74520
rect 106458 74508 106464 74520
rect 81676 74480 106464 74508
rect 81676 74468 81682 74480
rect 106458 74468 106464 74480
rect 106516 74508 106522 74520
rect 210418 74508 210424 74520
rect 106516 74480 210424 74508
rect 106516 74468 106522 74480
rect 210418 74468 210424 74480
rect 210476 74468 210482 74520
rect 212626 74468 212632 74520
rect 212684 74508 212690 74520
rect 269758 74508 269764 74520
rect 212684 74480 269764 74508
rect 212684 74468 212690 74480
rect 269758 74468 269764 74480
rect 269816 74468 269822 74520
rect 57882 73788 57888 73840
rect 57940 73828 57946 73840
rect 185578 73828 185584 73840
rect 57940 73800 185584 73828
rect 57940 73788 57946 73800
rect 185578 73788 185584 73800
rect 185636 73788 185642 73840
rect 212626 73176 212632 73228
rect 212684 73216 212690 73228
rect 213178 73216 213184 73228
rect 212684 73188 213184 73216
rect 212684 73176 212690 73188
rect 213178 73176 213184 73188
rect 213236 73176 213242 73228
rect 86954 73108 86960 73160
rect 87012 73148 87018 73160
rect 215294 73148 215300 73160
rect 87012 73120 215300 73148
rect 87012 73108 87018 73120
rect 215294 73108 215300 73120
rect 215352 73108 215358 73160
rect 162210 73040 162216 73092
rect 162268 73080 162274 73092
rect 237558 73080 237564 73092
rect 162268 73052 237564 73080
rect 162268 73040 162274 73052
rect 237558 73040 237564 73052
rect 237616 73040 237622 73092
rect 215294 71748 215300 71800
rect 215352 71788 215358 71800
rect 215938 71788 215944 71800
rect 215352 71760 215944 71788
rect 215352 71748 215358 71760
rect 215938 71748 215944 71760
rect 215996 71748 216002 71800
rect 237558 71748 237564 71800
rect 237616 71788 237622 71800
rect 238018 71788 238024 71800
rect 237616 71760 238024 71788
rect 237616 71748 237622 71760
rect 238018 71748 238024 71760
rect 238076 71748 238082 71800
rect 61930 71680 61936 71732
rect 61988 71720 61994 71732
rect 178862 71720 178868 71732
rect 61988 71692 178868 71720
rect 61988 71680 61994 71692
rect 178862 71680 178868 71692
rect 178920 71680 178926 71732
rect 180058 71680 180064 71732
rect 180116 71720 180122 71732
rect 228358 71720 228364 71732
rect 180116 71692 228364 71720
rect 180116 71680 180122 71692
rect 228358 71680 228364 71692
rect 228416 71680 228422 71732
rect 124858 71612 124864 71664
rect 124916 71652 124922 71664
rect 218054 71652 218060 71664
rect 124916 71624 218060 71652
rect 124916 71612 124922 71624
rect 218054 71612 218060 71624
rect 218112 71652 218118 71664
rect 218330 71652 218336 71664
rect 218112 71624 218336 71652
rect 218112 71612 218118 71624
rect 218330 71612 218336 71624
rect 218388 71612 218394 71664
rect 88242 71000 88248 71052
rect 88300 71040 88306 71052
rect 111150 71040 111156 71052
rect 88300 71012 111156 71040
rect 88300 71000 88306 71012
rect 111150 71000 111156 71012
rect 111208 71000 111214 71052
rect 218330 71000 218336 71052
rect 218388 71040 218394 71052
rect 351914 71040 351920 71052
rect 218388 71012 351920 71040
rect 218388 71000 218394 71012
rect 351914 71000 351920 71012
rect 351972 71000 351978 71052
rect 94498 70320 94504 70372
rect 94556 70360 94562 70372
rect 222286 70360 222292 70372
rect 94556 70332 222292 70360
rect 94556 70320 94562 70332
rect 222286 70320 222292 70332
rect 222344 70360 222350 70372
rect 222838 70360 222844 70372
rect 222344 70332 222844 70360
rect 222344 70320 222350 70332
rect 222838 70320 222844 70332
rect 222896 70320 222902 70372
rect 71682 69640 71688 69692
rect 71740 69680 71746 69692
rect 171778 69680 171784 69692
rect 71740 69652 171784 69680
rect 71740 69640 71746 69652
rect 171778 69640 171784 69652
rect 171836 69640 171842 69692
rect 193122 69640 193128 69692
rect 193180 69680 193186 69692
rect 270494 69680 270500 69692
rect 193180 69652 270500 69680
rect 193180 69640 193186 69652
rect 270494 69640 270500 69652
rect 270552 69640 270558 69692
rect 69198 68960 69204 69012
rect 69256 69000 69262 69012
rect 194778 69000 194784 69012
rect 69256 68972 194784 69000
rect 69256 68960 69262 68972
rect 194778 68960 194784 68972
rect 194836 69000 194842 69012
rect 195330 69000 195336 69012
rect 194836 68972 195336 69000
rect 194836 68960 194842 68972
rect 195330 68960 195336 68972
rect 195388 68960 195394 69012
rect 89622 68280 89628 68332
rect 89680 68320 89686 68332
rect 163498 68320 163504 68332
rect 89680 68292 163504 68320
rect 89680 68280 89686 68292
rect 163498 68280 163504 68292
rect 163556 68280 163562 68332
rect 192846 68280 192852 68332
rect 192904 68320 192910 68332
rect 281534 68320 281540 68332
rect 192904 68292 281540 68320
rect 192904 68280 192910 68292
rect 281534 68280 281540 68292
rect 281592 68280 281598 68332
rect 71866 67532 71872 67584
rect 71924 67572 71930 67584
rect 197354 67572 197360 67584
rect 71924 67544 197360 67572
rect 71924 67532 71930 67544
rect 197354 67532 197360 67544
rect 197412 67572 197418 67584
rect 197998 67572 198004 67584
rect 197412 67544 198004 67572
rect 197412 67532 197418 67544
rect 197998 67532 198004 67544
rect 198056 67532 198062 67584
rect 201494 67532 201500 67584
rect 201552 67572 201558 67584
rect 202138 67572 202144 67584
rect 201552 67544 202144 67572
rect 201552 67532 201558 67544
rect 202138 67532 202144 67544
rect 202196 67572 202202 67584
rect 293954 67572 293960 67584
rect 202196 67544 293960 67572
rect 202196 67532 202202 67544
rect 293954 67532 293960 67544
rect 294012 67532 294018 67584
rect 166350 67464 166356 67516
rect 166408 67504 166414 67516
rect 231854 67504 231860 67516
rect 166408 67476 231860 67504
rect 166408 67464 166414 67476
rect 231854 67464 231860 67476
rect 231912 67464 231918 67516
rect 100018 66172 100024 66224
rect 100076 66212 100082 66224
rect 241514 66212 241520 66224
rect 100076 66184 241520 66212
rect 100076 66172 100082 66184
rect 241514 66172 241520 66184
rect 241572 66172 241578 66224
rect 75822 65492 75828 65544
rect 75880 65532 75886 65544
rect 177298 65532 177304 65544
rect 75880 65504 177304 65532
rect 75880 65492 75886 65504
rect 177298 65492 177304 65504
rect 177356 65492 177362 65544
rect 187602 65492 187608 65544
rect 187660 65532 187666 65544
rect 214558 65532 214564 65544
rect 187660 65504 214564 65532
rect 187660 65492 187666 65504
rect 214558 65492 214564 65504
rect 214616 65492 214622 65544
rect 85574 64812 85580 64864
rect 85632 64852 85638 64864
rect 118786 64852 118792 64864
rect 85632 64824 118792 64852
rect 85632 64812 85638 64824
rect 118786 64812 118792 64824
rect 118844 64852 118850 64864
rect 213178 64852 213184 64864
rect 118844 64824 213184 64852
rect 118844 64812 118850 64824
rect 213178 64812 213184 64824
rect 213236 64812 213242 64864
rect 152550 64744 152556 64796
rect 152608 64784 152614 64796
rect 227714 64784 227720 64796
rect 152608 64756 227720 64784
rect 152608 64744 152614 64756
rect 227714 64744 227720 64756
rect 227772 64744 227778 64796
rect 106182 64132 106188 64184
rect 106240 64172 106246 64184
rect 126330 64172 126336 64184
rect 106240 64144 126336 64172
rect 106240 64132 106246 64144
rect 126330 64132 126336 64144
rect 126388 64132 126394 64184
rect 227714 63520 227720 63572
rect 227772 63560 227778 63572
rect 228358 63560 228364 63572
rect 227772 63532 228364 63560
rect 227772 63520 227778 63532
rect 228358 63520 228364 63532
rect 228416 63520 228422 63572
rect 193306 63452 193312 63504
rect 193364 63492 193370 63504
rect 295426 63492 295432 63504
rect 193364 63464 295432 63492
rect 193364 63452 193370 63464
rect 295426 63452 295432 63464
rect 295484 63452 295490 63504
rect 122098 63384 122104 63436
rect 122156 63424 122162 63436
rect 217318 63424 217324 63436
rect 122156 63396 217324 63424
rect 122156 63384 122162 63396
rect 217318 63384 217324 63396
rect 217376 63384 217382 63436
rect 85482 62840 85488 62892
rect 85540 62880 85546 62892
rect 115198 62880 115204 62892
rect 85540 62852 115204 62880
rect 85540 62840 85546 62852
rect 115198 62840 115204 62852
rect 115256 62840 115262 62892
rect 81342 62772 81348 62824
rect 81400 62812 81406 62824
rect 130470 62812 130476 62824
rect 81400 62784 130476 62812
rect 81400 62772 81406 62784
rect 130470 62772 130476 62784
rect 130528 62772 130534 62824
rect 88150 62024 88156 62076
rect 88208 62064 88214 62076
rect 216030 62064 216036 62076
rect 88208 62036 216036 62064
rect 88208 62024 88214 62036
rect 216030 62024 216036 62036
rect 216088 62024 216094 62076
rect 71038 61956 71044 62008
rect 71096 61996 71102 62008
rect 194686 61996 194692 62008
rect 71096 61968 194692 61996
rect 71096 61956 71102 61968
rect 194686 61956 194692 61968
rect 194744 61956 194750 62008
rect 195330 61956 195336 62008
rect 195388 61996 195394 62008
rect 285674 61996 285680 62008
rect 195388 61968 285680 61996
rect 195388 61956 195394 61968
rect 285674 61956 285680 61968
rect 285732 61996 285738 62008
rect 286594 61996 286600 62008
rect 285732 61968 286600 61996
rect 285732 61956 285738 61968
rect 286594 61956 286600 61968
rect 286652 61956 286658 62008
rect 286594 61344 286600 61396
rect 286652 61384 286658 61396
rect 345014 61384 345020 61396
rect 286652 61356 345020 61384
rect 286652 61344 286658 61356
rect 345014 61344 345020 61356
rect 345072 61344 345078 61396
rect 194686 60732 194692 60784
rect 194744 60772 194750 60784
rect 195238 60772 195244 60784
rect 194744 60744 195244 60772
rect 194744 60732 194750 60744
rect 195238 60732 195244 60744
rect 195296 60732 195302 60784
rect 67266 60664 67272 60716
rect 67324 60704 67330 60716
rect 183554 60704 183560 60716
rect 67324 60676 183560 60704
rect 67324 60664 67330 60676
rect 183554 60664 183560 60676
rect 183612 60704 183618 60716
rect 184290 60704 184296 60716
rect 183612 60676 184296 60704
rect 183612 60664 183618 60676
rect 184290 60664 184296 60676
rect 184348 60664 184354 60716
rect 97258 60596 97264 60648
rect 97316 60636 97322 60648
rect 204346 60636 204352 60648
rect 97316 60608 204352 60636
rect 97316 60596 97322 60608
rect 204346 60596 204352 60608
rect 204404 60596 204410 60648
rect 204346 60188 204352 60240
rect 204404 60228 204410 60240
rect 204990 60228 204996 60240
rect 204404 60200 204996 60228
rect 204404 60188 204410 60200
rect 204990 60188 204996 60200
rect 205048 60188 205054 60240
rect 193214 59984 193220 60036
rect 193272 60024 193278 60036
rect 264974 60024 264980 60036
rect 193272 59996 264980 60024
rect 193272 59984 193278 59996
rect 264974 59984 264980 59996
rect 265032 59984 265038 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 51718 59344 51724 59356
rect 3108 59316 51724 59344
rect 3108 59304 3114 59316
rect 51718 59304 51724 59316
rect 51776 59304 51782 59356
rect 67634 59304 67640 59356
rect 67692 59344 67698 59356
rect 193306 59344 193312 59356
rect 67692 59316 193312 59344
rect 67692 59304 67698 59316
rect 193306 59304 193312 59316
rect 193364 59344 193370 59356
rect 193858 59344 193864 59356
rect 193364 59316 193864 59344
rect 193364 59304 193370 59316
rect 193858 59304 193864 59316
rect 193916 59304 193922 59356
rect 207106 59344 207112 59356
rect 200086 59316 207112 59344
rect 112438 59236 112444 59288
rect 112496 59276 112502 59288
rect 200086 59276 200114 59316
rect 207106 59304 207112 59316
rect 207164 59344 207170 59356
rect 207658 59344 207664 59356
rect 207164 59316 207664 59344
rect 207164 59304 207170 59316
rect 207658 59304 207664 59316
rect 207716 59304 207722 59356
rect 289814 59344 289820 59356
rect 209746 59316 289820 59344
rect 112496 59248 200114 59276
rect 112496 59236 112502 59248
rect 200114 59168 200120 59220
rect 200172 59208 200178 59220
rect 209746 59208 209774 59316
rect 289814 59304 289820 59316
rect 289872 59304 289878 59356
rect 200172 59180 209774 59208
rect 200172 59168 200178 59180
rect 93762 57876 93768 57928
rect 93820 57916 93826 57928
rect 222194 57916 222200 57928
rect 93820 57888 222200 57916
rect 93820 57876 93826 57888
rect 222194 57876 222200 57888
rect 222252 57916 222258 57928
rect 222930 57916 222936 57928
rect 222252 57888 222936 57916
rect 222252 57876 222258 57888
rect 222930 57876 222936 57888
rect 222988 57876 222994 57928
rect 73798 57808 73804 57860
rect 73856 57848 73862 57860
rect 200114 57848 200120 57860
rect 73856 57820 200120 57848
rect 73856 57808 73862 57820
rect 200114 57808 200120 57820
rect 200172 57848 200178 57860
rect 200758 57848 200764 57860
rect 200172 57820 200764 57848
rect 200172 57808 200178 57820
rect 200758 57808 200764 57820
rect 200816 57808 200822 57860
rect 74534 56516 74540 56568
rect 74592 56556 74598 56568
rect 202138 56556 202144 56568
rect 74592 56528 202144 56556
rect 74592 56516 74598 56528
rect 202138 56516 202144 56528
rect 202196 56516 202202 56568
rect 197998 56448 198004 56500
rect 198056 56488 198062 56500
rect 247034 56488 247040 56500
rect 198056 56460 247040 56488
rect 198056 56448 198062 56460
rect 247034 56448 247040 56460
rect 247092 56488 247098 56500
rect 247586 56488 247592 56500
rect 247092 56460 247592 56488
rect 247092 56448 247098 56460
rect 247586 56448 247592 56460
rect 247644 56448 247650 56500
rect 247586 55836 247592 55888
rect 247644 55876 247650 55888
rect 342254 55876 342260 55888
rect 247644 55848 342260 55876
rect 247644 55836 247650 55848
rect 342254 55836 342260 55848
rect 342312 55836 342318 55888
rect 103330 54544 103336 54596
rect 103388 54584 103394 54596
rect 133230 54584 133236 54596
rect 103388 54556 133236 54584
rect 103388 54544 103394 54556
rect 133230 54544 133236 54556
rect 133288 54544 133294 54596
rect 73062 54476 73068 54528
rect 73120 54516 73126 54528
rect 145558 54516 145564 54528
rect 73120 54488 145564 54516
rect 73120 54476 73126 54488
rect 145558 54476 145564 54488
rect 145616 54476 145622 54528
rect 184290 54476 184296 54528
rect 184348 54516 184354 54528
rect 320174 54516 320180 54528
rect 184348 54488 320180 54516
rect 184348 54476 184354 54488
rect 320174 54476 320180 54488
rect 320232 54476 320238 54528
rect 97258 53048 97264 53100
rect 97316 53088 97322 53100
rect 141510 53088 141516 53100
rect 97316 53060 141516 53088
rect 97316 53048 97322 53060
rect 141510 53048 141516 53060
rect 141568 53048 141574 53100
rect 214650 53048 214656 53100
rect 214708 53088 214714 53100
rect 286318 53088 286324 53100
rect 214708 53060 286324 53088
rect 214708 53048 214714 53060
rect 286318 53048 286324 53060
rect 286376 53048 286382 53100
rect 61930 51688 61936 51740
rect 61988 51728 61994 51740
rect 144178 51728 144184 51740
rect 61988 51700 144184 51728
rect 61988 51688 61994 51700
rect 144178 51688 144184 51700
rect 144236 51688 144242 51740
rect 186958 51688 186964 51740
rect 187016 51728 187022 51740
rect 580166 51728 580172 51740
rect 187016 51700 580172 51728
rect 187016 51688 187022 51700
rect 580166 51688 580172 51700
rect 580224 51688 580230 51740
rect 3970 50328 3976 50380
rect 4028 50368 4034 50380
rect 142890 50368 142896 50380
rect 4028 50340 142896 50368
rect 4028 50328 4034 50340
rect 142890 50328 142896 50340
rect 142948 50328 142954 50380
rect 182818 50328 182824 50380
rect 182876 50368 182882 50380
rect 335354 50368 335360 50380
rect 182876 50340 335360 50368
rect 182876 50328 182882 50340
rect 335354 50328 335360 50340
rect 335412 50328 335418 50380
rect 59262 48968 59268 49020
rect 59320 49008 59326 49020
rect 151170 49008 151176 49020
rect 59320 48980 151176 49008
rect 59320 48968 59326 48980
rect 151170 48968 151176 48980
rect 151228 48968 151234 49020
rect 193030 48968 193036 49020
rect 193088 49008 193094 49020
rect 310514 49008 310520 49020
rect 193088 48980 310520 49008
rect 193088 48968 193094 48980
rect 310514 48968 310520 48980
rect 310572 48968 310578 49020
rect 65518 47540 65524 47592
rect 65576 47580 65582 47592
rect 149698 47580 149704 47592
rect 65576 47552 149704 47580
rect 65576 47540 65582 47552
rect 149698 47540 149704 47552
rect 149756 47540 149762 47592
rect 181990 47540 181996 47592
rect 182048 47580 182054 47592
rect 226978 47580 226984 47592
rect 182048 47552 226984 47580
rect 182048 47540 182054 47552
rect 226978 47540 226984 47552
rect 227036 47540 227042 47592
rect 119890 46248 119896 46300
rect 119948 46288 119954 46300
rect 153838 46288 153844 46300
rect 119948 46260 153844 46288
rect 119948 46248 119954 46260
rect 153838 46248 153844 46260
rect 153896 46248 153902 46300
rect 3326 46180 3332 46232
rect 3384 46220 3390 46232
rect 65610 46220 65616 46232
rect 3384 46192 65616 46220
rect 3384 46180 3390 46192
rect 65610 46180 65616 46192
rect 65668 46180 65674 46232
rect 67542 46180 67548 46232
rect 67600 46220 67606 46232
rect 128998 46220 129004 46232
rect 67600 46192 129004 46220
rect 67600 46180 67606 46192
rect 128998 46180 129004 46192
rect 129056 46180 129062 46232
rect 217318 46180 217324 46232
rect 217376 46220 217382 46232
rect 291930 46220 291936 46232
rect 217376 46192 291936 46220
rect 217376 46180 217382 46192
rect 291930 46180 291936 46192
rect 291988 46180 291994 46232
rect 190270 44820 190276 44872
rect 190328 44860 190334 44872
rect 288434 44860 288440 44872
rect 190328 44832 288440 44860
rect 190328 44820 190334 44832
rect 288434 44820 288440 44832
rect 288492 44820 288498 44872
rect 77202 43392 77208 43444
rect 77260 43432 77266 43444
rect 146938 43432 146944 43444
rect 77260 43404 146944 43432
rect 77260 43392 77266 43404
rect 146938 43392 146944 43404
rect 146996 43392 147002 43444
rect 191650 43392 191656 43444
rect 191708 43432 191714 43444
rect 305730 43432 305736 43444
rect 191708 43404 305736 43432
rect 191708 43392 191714 43404
rect 305730 43392 305736 43404
rect 305788 43392 305794 43444
rect 79318 42032 79324 42084
rect 79376 42072 79382 42084
rect 137370 42072 137376 42084
rect 79376 42044 137376 42072
rect 79376 42032 79382 42044
rect 137370 42032 137376 42044
rect 137428 42032 137434 42084
rect 305638 42032 305644 42084
rect 305696 42072 305702 42084
rect 329834 42072 329840 42084
rect 305696 42044 329840 42072
rect 305696 42032 305702 42044
rect 329834 42032 329840 42044
rect 329892 42032 329898 42084
rect 99282 40672 99288 40724
rect 99340 40712 99346 40724
rect 162118 40712 162124 40724
rect 99340 40684 162124 40712
rect 99340 40672 99346 40684
rect 162118 40672 162124 40684
rect 162176 40672 162182 40724
rect 239398 40672 239404 40724
rect 239456 40712 239462 40724
rect 349798 40712 349804 40724
rect 239456 40684 349804 40712
rect 239456 40672 239462 40684
rect 349798 40672 349804 40684
rect 349856 40672 349862 40724
rect 82722 39312 82728 39364
rect 82780 39352 82786 39364
rect 167638 39352 167644 39364
rect 82780 39324 167644 39352
rect 82780 39312 82786 39324
rect 167638 39312 167644 39324
rect 167696 39312 167702 39364
rect 199378 39312 199384 39364
rect 199436 39352 199442 39364
rect 233878 39352 233884 39364
rect 199436 39324 233884 39352
rect 199436 39312 199442 39324
rect 233878 39312 233884 39324
rect 233936 39312 233942 39364
rect 244918 37952 244924 38004
rect 244976 37992 244982 38004
rect 258810 37992 258816 38004
rect 244976 37964 258816 37992
rect 244976 37952 244982 37964
rect 258810 37952 258816 37964
rect 258868 37952 258874 38004
rect 68922 37884 68928 37936
rect 68980 37924 68986 37936
rect 174538 37924 174544 37936
rect 68980 37896 174544 37924
rect 68980 37884 68986 37896
rect 174538 37884 174544 37896
rect 174596 37884 174602 37936
rect 184198 37884 184204 37936
rect 184256 37924 184262 37936
rect 249794 37924 249800 37936
rect 184256 37896 249800 37924
rect 184256 37884 184262 37896
rect 249794 37884 249800 37896
rect 249852 37884 249858 37936
rect 67726 36524 67732 36576
rect 67784 36564 67790 36576
rect 125594 36564 125600 36576
rect 67784 36536 125600 36564
rect 67784 36524 67790 36536
rect 125594 36524 125600 36536
rect 125652 36524 125658 36576
rect 214558 36524 214564 36576
rect 214616 36564 214622 36576
rect 327074 36564 327080 36576
rect 214616 36536 327080 36564
rect 214616 36524 214622 36536
rect 327074 36524 327080 36536
rect 327132 36524 327138 36576
rect 75178 35164 75184 35216
rect 75236 35204 75242 35216
rect 155310 35204 155316 35216
rect 75236 35176 155316 35204
rect 75236 35164 75242 35176
rect 155310 35164 155316 35176
rect 155368 35164 155374 35216
rect 222930 35164 222936 35216
rect 222988 35204 222994 35216
rect 301498 35204 301504 35216
rect 222988 35176 301504 35204
rect 222988 35164 222994 35176
rect 301498 35164 301504 35176
rect 301556 35164 301562 35216
rect 55122 33736 55128 33788
rect 55180 33776 55186 33788
rect 140038 33776 140044 33788
rect 55180 33748 140044 33776
rect 55180 33736 55186 33748
rect 140038 33736 140044 33748
rect 140096 33736 140102 33788
rect 200758 33736 200764 33788
rect 200816 33776 200822 33788
rect 340966 33776 340972 33788
rect 200816 33748 340972 33776
rect 200816 33736 200822 33748
rect 340966 33736 340972 33748
rect 341024 33736 341030 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 54478 33096 54484 33108
rect 3568 33068 54484 33096
rect 3568 33056 3574 33068
rect 54478 33056 54484 33068
rect 54536 33056 54542 33108
rect 64782 32376 64788 32428
rect 64840 32416 64846 32428
rect 175918 32416 175924 32428
rect 64840 32388 175924 32416
rect 64840 32376 64846 32388
rect 175918 32376 175924 32388
rect 175976 32376 175982 32428
rect 44082 31016 44088 31068
rect 44140 31056 44146 31068
rect 169018 31056 169024 31068
rect 44140 31028 169024 31056
rect 44140 31016 44146 31028
rect 169018 31016 169024 31028
rect 169076 31016 169082 31068
rect 195238 31016 195244 31068
rect 195296 31056 195302 31068
rect 311894 31056 311900 31068
rect 195296 31028 311900 31056
rect 195296 31016 195302 31028
rect 311894 31016 311900 31028
rect 311952 31016 311958 31068
rect 46842 29588 46848 29640
rect 46900 29628 46906 29640
rect 166258 29628 166264 29640
rect 46900 29600 166264 29628
rect 46900 29588 46906 29600
rect 166258 29588 166264 29600
rect 166316 29588 166322 29640
rect 193858 29588 193864 29640
rect 193916 29628 193922 29640
rect 291194 29628 291200 29640
rect 193916 29600 291200 29628
rect 193916 29588 193922 29600
rect 291194 29588 291200 29600
rect 291252 29588 291258 29640
rect 291838 29588 291844 29640
rect 291896 29628 291902 29640
rect 325694 29628 325700 29640
rect 291896 29600 325700 29628
rect 291896 29588 291902 29600
rect 325694 29588 325700 29600
rect 325752 29588 325758 29640
rect 86770 28228 86776 28280
rect 86828 28268 86834 28280
rect 164878 28268 164884 28280
rect 86828 28240 164884 28268
rect 86828 28228 86834 28240
rect 164878 28228 164884 28240
rect 164936 28228 164942 28280
rect 213178 28228 213184 28280
rect 213236 28268 213242 28280
rect 287054 28268 287060 28280
rect 213236 28240 287060 28268
rect 213236 28228 213242 28240
rect 287054 28228 287060 28240
rect 287112 28228 287118 28280
rect 93762 26868 93768 26920
rect 93820 26908 93826 26920
rect 157978 26908 157984 26920
rect 93820 26880 157984 26908
rect 93820 26868 93826 26880
rect 157978 26868 157984 26880
rect 158036 26868 158042 26920
rect 56502 25508 56508 25560
rect 56560 25548 56566 25560
rect 135898 25548 135904 25560
rect 56560 25520 135904 25548
rect 56560 25508 56566 25520
rect 135898 25508 135904 25520
rect 135956 25508 135962 25560
rect 209682 25508 209688 25560
rect 209740 25548 209746 25560
rect 278774 25548 278780 25560
rect 209740 25520 278780 25548
rect 209740 25508 209746 25520
rect 278774 25508 278780 25520
rect 278832 25508 278838 25560
rect 66162 24080 66168 24132
rect 66220 24120 66226 24132
rect 138658 24120 138664 24132
rect 66220 24092 138664 24120
rect 66220 24080 66226 24092
rect 138658 24080 138664 24092
rect 138716 24080 138722 24132
rect 207658 24080 207664 24132
rect 207716 24120 207722 24132
rect 246298 24120 246304 24132
rect 207716 24092 246304 24120
rect 207716 24080 207722 24092
rect 246298 24080 246304 24092
rect 246356 24080 246362 24132
rect 78582 22720 78588 22772
rect 78640 22760 78646 22772
rect 178678 22760 178684 22772
rect 78640 22732 178684 22760
rect 78640 22720 78646 22732
rect 178678 22720 178684 22732
rect 178736 22720 178742 22772
rect 213822 22720 213828 22772
rect 213880 22760 213886 22772
rect 334066 22760 334072 22772
rect 213880 22732 334072 22760
rect 213880 22720 213886 22732
rect 334066 22720 334072 22732
rect 334124 22720 334130 22772
rect 74442 21360 74448 21412
rect 74500 21400 74506 21412
rect 108390 21400 108396 21412
rect 74500 21372 108396 21400
rect 74500 21360 74506 21372
rect 108390 21360 108396 21372
rect 108448 21360 108454 21412
rect 111610 21360 111616 21412
rect 111668 21400 111674 21412
rect 127710 21400 127716 21412
rect 111668 21372 127716 21400
rect 111668 21360 111674 21372
rect 127710 21360 127716 21372
rect 127768 21360 127774 21412
rect 204162 21360 204168 21412
rect 204220 21400 204226 21412
rect 324406 21400 324412 21412
rect 204220 21372 324412 21400
rect 204220 21360 204226 21372
rect 324406 21360 324412 21372
rect 324464 21360 324470 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 93118 20652 93124 20664
rect 3476 20624 93124 20652
rect 3476 20612 3482 20624
rect 93118 20612 93124 20624
rect 93176 20612 93182 20664
rect 242802 20000 242808 20052
rect 242860 20040 242866 20052
rect 284386 20040 284392 20052
rect 242860 20012 284392 20040
rect 242860 20000 242866 20012
rect 284386 20000 284392 20012
rect 284444 20000 284450 20052
rect 91002 19932 91008 19984
rect 91060 19972 91066 19984
rect 141418 19972 141424 19984
rect 91060 19944 141424 19972
rect 91060 19932 91066 19944
rect 141418 19932 141424 19944
rect 141476 19932 141482 19984
rect 185670 19932 185676 19984
rect 185728 19972 185734 19984
rect 242986 19972 242992 19984
rect 185728 19944 242992 19972
rect 185728 19932 185734 19944
rect 242986 19932 242992 19944
rect 243044 19932 243050 19984
rect 50982 18572 50988 18624
rect 51040 18612 51046 18624
rect 170398 18612 170404 18624
rect 51040 18584 170404 18612
rect 51040 18572 51046 18584
rect 170398 18572 170404 18584
rect 170456 18572 170462 18624
rect 222838 18572 222844 18624
rect 222896 18612 222902 18624
rect 339494 18612 339500 18624
rect 222896 18584 339500 18612
rect 222896 18572 222902 18584
rect 339494 18572 339500 18584
rect 339552 18572 339558 18624
rect 228358 17212 228364 17264
rect 228416 17252 228422 17264
rect 331214 17252 331220 17264
rect 228416 17224 331220 17252
rect 228416 17212 228422 17224
rect 331214 17212 331220 17224
rect 331272 17212 331278 17264
rect 240778 15852 240784 15904
rect 240836 15892 240842 15904
rect 253474 15892 253480 15904
rect 240836 15864 253480 15892
rect 240836 15852 240842 15864
rect 253474 15852 253480 15864
rect 253532 15852 253538 15904
rect 253198 15172 253204 15224
rect 253256 15212 253262 15224
rect 256694 15212 256700 15224
rect 253256 15184 256700 15212
rect 253256 15172 253262 15184
rect 256694 15172 256700 15184
rect 256752 15172 256758 15224
rect 95050 14424 95056 14476
rect 95108 14464 95114 14476
rect 152458 14464 152464 14476
rect 95108 14436 152464 14464
rect 95108 14424 95114 14436
rect 152458 14424 152464 14436
rect 152516 14424 152522 14476
rect 204990 14424 204996 14476
rect 205048 14464 205054 14476
rect 344554 14464 344560 14476
rect 205048 14436 344560 14464
rect 205048 14424 205054 14436
rect 344554 14424 344560 14436
rect 344612 14424 344618 14476
rect 70210 13064 70216 13116
rect 70268 13104 70274 13116
rect 142798 13104 142804 13116
rect 70268 13076 142804 13104
rect 70268 13064 70274 13076
rect 142798 13064 142804 13076
rect 142856 13064 142862 13116
rect 249058 13064 249064 13116
rect 249116 13104 249122 13116
rect 302878 13104 302884 13116
rect 249116 13076 302884 13104
rect 249116 13064 249122 13076
rect 302878 13064 302884 13076
rect 302936 13064 302942 13116
rect 84102 11704 84108 11756
rect 84160 11744 84166 11756
rect 131758 11744 131764 11756
rect 84160 11716 131764 11744
rect 84160 11704 84166 11716
rect 131758 11704 131764 11716
rect 131816 11704 131822 11756
rect 215938 11704 215944 11756
rect 215996 11744 216002 11756
rect 266538 11744 266544 11756
rect 215996 11716 266544 11744
rect 215996 11704 216002 11716
rect 266538 11704 266544 11716
rect 266596 11704 266602 11756
rect 79686 10276 79692 10328
rect 79744 10316 79750 10328
rect 148410 10316 148416 10328
rect 79744 10288 148416 10316
rect 79744 10276 79750 10288
rect 148410 10276 148416 10288
rect 148468 10276 148474 10328
rect 202138 10276 202144 10328
rect 202196 10316 202202 10328
rect 321554 10316 321560 10328
rect 202196 10288 321560 10316
rect 202196 10276 202202 10288
rect 321554 10276 321560 10288
rect 321612 10276 321618 10328
rect 99834 8984 99840 9036
rect 99892 9024 99898 9036
rect 173158 9024 173164 9036
rect 99892 8996 173164 9024
rect 99892 8984 99898 8996
rect 173158 8984 173164 8996
rect 173216 8984 173222 9036
rect 566 8916 572 8968
rect 624 8956 630 8968
rect 101398 8956 101404 8968
rect 624 8928 101404 8956
rect 624 8916 630 8928
rect 101398 8916 101404 8928
rect 101456 8916 101462 8968
rect 196618 8916 196624 8968
rect 196676 8956 196682 8968
rect 258258 8956 258264 8968
rect 196676 8928 258264 8956
rect 196676 8916 196682 8928
rect 258258 8916 258264 8928
rect 258316 8916 258322 8968
rect 320818 8916 320824 8968
rect 320876 8956 320882 8968
rect 332686 8956 332692 8968
rect 320876 8928 332692 8956
rect 320876 8916 320882 8928
rect 332686 8916 332692 8928
rect 332744 8916 332750 8968
rect 250530 7624 250536 7676
rect 250588 7664 250594 7676
rect 261754 7664 261760 7676
rect 250588 7636 261760 7664
rect 250588 7624 250594 7636
rect 261754 7624 261760 7636
rect 261812 7624 261818 7676
rect 266998 7624 267004 7676
rect 267056 7664 267062 7676
rect 276014 7664 276020 7676
rect 267056 7636 276020 7664
rect 267056 7624 267062 7636
rect 276014 7624 276020 7636
rect 276072 7624 276078 7676
rect 59630 7556 59636 7608
rect 59688 7596 59694 7608
rect 155218 7596 155224 7608
rect 59688 7568 155224 7596
rect 59688 7556 59694 7568
rect 155218 7556 155224 7568
rect 155276 7556 155282 7608
rect 191742 7556 191748 7608
rect 191800 7596 191806 7608
rect 249794 7596 249800 7608
rect 191800 7568 249800 7596
rect 191800 7556 191806 7568
rect 249794 7556 249800 7568
rect 249852 7556 249858 7608
rect 258718 7556 258724 7608
rect 258776 7596 258782 7608
rect 269114 7596 269120 7608
rect 258776 7568 269120 7596
rect 258776 7556 258782 7568
rect 269114 7556 269120 7568
rect 269172 7556 269178 7608
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 52546 6128 52552 6180
rect 52604 6168 52610 6180
rect 159358 6168 159364 6180
rect 52604 6140 159364 6168
rect 52604 6128 52610 6140
rect 159358 6128 159364 6140
rect 159416 6128 159422 6180
rect 224862 6128 224868 6180
rect 224920 6168 224926 6180
rect 254670 6168 254676 6180
rect 224920 6140 254676 6168
rect 224920 6128 224926 6140
rect 254670 6128 254676 6140
rect 254728 6128 254734 6180
rect 271138 6128 271144 6180
rect 271196 6168 271202 6180
rect 297266 6168 297272 6180
rect 271196 6140 297272 6168
rect 271196 6128 271202 6140
rect 297266 6128 297272 6140
rect 297324 6128 297330 6180
rect 305730 5516 305736 5568
rect 305788 5556 305794 5568
rect 309042 5556 309048 5568
rect 305788 5528 309048 5556
rect 305788 5516 305794 5528
rect 309042 5516 309048 5528
rect 309100 5516 309106 5568
rect 349798 5516 349804 5568
rect 349856 5556 349862 5568
rect 351638 5556 351644 5568
rect 349856 5528 351644 5556
rect 349856 5516 349862 5528
rect 351638 5516 351644 5528
rect 351696 5516 351702 5568
rect 96246 4836 96252 4888
rect 96304 4876 96310 4888
rect 151078 4876 151084 4888
rect 96304 4848 151084 4876
rect 96304 4836 96310 4848
rect 151078 4836 151084 4848
rect 151136 4836 151142 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 97258 4808 97264 4820
rect 1728 4780 97264 4808
rect 1728 4768 1734 4780
rect 97258 4768 97264 4780
rect 97316 4768 97322 4820
rect 204898 4768 204904 4820
rect 204956 4808 204962 4820
rect 274818 4808 274824 4820
rect 204956 4780 274824 4808
rect 204956 4768 204962 4780
rect 274818 4768 274824 4780
rect 274876 4768 274882 4820
rect 331858 4496 331864 4548
rect 331916 4536 331922 4548
rect 337470 4536 337476 4548
rect 331916 4508 337476 4536
rect 331916 4496 331922 4508
rect 337470 4496 337476 4508
rect 337528 4496 337534 4548
rect 238018 4360 238024 4412
rect 238076 4400 238082 4412
rect 239306 4400 239312 4412
rect 238076 4372 239312 4400
rect 238076 4360 238082 4372
rect 239306 4360 239312 4372
rect 239364 4360 239370 4412
rect 134518 4156 134524 4208
rect 134576 4196 134582 4208
rect 136450 4196 136456 4208
rect 134576 4168 136456 4196
rect 134576 4156 134582 4168
rect 136450 4156 136456 4168
rect 136508 4156 136514 4208
rect 342990 4088 342996 4140
rect 343048 4128 343054 4140
rect 346946 4128 346952 4140
rect 343048 4100 346952 4128
rect 343048 4088 343054 4100
rect 346946 4088 346952 4100
rect 347004 4088 347010 4140
rect 233878 4020 233884 4072
rect 233936 4060 233942 4072
rect 240502 4060 240508 4072
rect 233936 4032 240508 4060
rect 233936 4020 233942 4032
rect 240502 4020 240508 4032
rect 240560 4020 240566 4072
rect 44266 3884 44272 3936
rect 44324 3924 44330 3936
rect 47578 3924 47584 3936
rect 44324 3896 47584 3924
rect 44324 3884 44330 3896
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 304350 3748 304356 3800
rect 304408 3788 304414 3800
rect 307938 3788 307944 3800
rect 304408 3760 307944 3788
rect 304408 3748 304414 3760
rect 307938 3748 307944 3760
rect 307996 3748 308002 3800
rect 27706 3612 27712 3664
rect 27764 3652 27770 3664
rect 32398 3652 32404 3664
rect 27764 3624 32404 3652
rect 27764 3612 27770 3624
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 60826 3544 60832 3596
rect 60884 3584 60890 3596
rect 61930 3584 61936 3596
rect 60884 3556 61936 3584
rect 60884 3544 60890 3556
rect 61930 3544 61936 3556
rect 61988 3544 61994 3596
rect 101030 3544 101036 3596
rect 101088 3584 101094 3596
rect 101088 3556 103514 3584
rect 101088 3544 101094 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20622 3516 20628 3528
rect 19484 3488 20628 3516
rect 19484 3476 19490 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 44082 3516 44088 3528
rect 43128 3488 44088 3516
rect 43128 3476 43134 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 64322 3476 64328 3528
rect 64380 3516 64386 3528
rect 64782 3516 64788 3528
rect 64380 3488 64788 3516
rect 64380 3476 64386 3488
rect 64782 3476 64788 3488
rect 64840 3476 64846 3528
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 70210 3516 70216 3528
rect 69164 3488 70216 3516
rect 69164 3476 69170 3488
rect 70210 3476 70216 3488
rect 70268 3476 70274 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 73798 3476 73804 3528
rect 73856 3516 73862 3528
rect 74442 3516 74448 3528
rect 73856 3488 74448 3516
rect 73856 3476 73862 3488
rect 74442 3476 74448 3488
rect 74500 3476 74506 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 80882 3476 80888 3528
rect 80940 3516 80946 3528
rect 81342 3516 81348 3528
rect 80940 3488 81348 3516
rect 80940 3476 80946 3488
rect 81342 3476 81348 3488
rect 81400 3476 81406 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 82722 3516 82728 3528
rect 82136 3488 82728 3516
rect 82136 3476 82142 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 84102 3516 84108 3528
rect 83332 3488 84108 3516
rect 83332 3476 83338 3488
rect 84102 3476 84108 3488
rect 84160 3476 84166 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 85666 3476 85672 3528
rect 85724 3516 85730 3528
rect 86770 3516 86776 3528
rect 85724 3488 86776 3516
rect 85724 3476 85730 3488
rect 86770 3476 86776 3488
rect 86828 3476 86834 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 89622 3516 89628 3528
rect 89220 3488 89628 3516
rect 89220 3476 89226 3488
rect 89622 3476 89628 3488
rect 89680 3476 89686 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 92750 3476 92756 3528
rect 92808 3516 92814 3528
rect 93762 3516 93768 3528
rect 92808 3488 93768 3516
rect 92808 3476 92814 3488
rect 93762 3476 93768 3488
rect 93820 3476 93826 3528
rect 93946 3476 93952 3528
rect 94004 3516 94010 3528
rect 95050 3516 95056 3528
rect 94004 3488 95056 3516
rect 94004 3476 94010 3488
rect 95050 3476 95056 3488
rect 95108 3476 95114 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 102226 3476 102232 3528
rect 102284 3516 102290 3528
rect 103238 3516 103244 3528
rect 102284 3488 103244 3516
rect 102284 3476 102290 3488
rect 103238 3476 103244 3488
rect 103296 3476 103302 3528
rect 103486 3516 103514 3556
rect 114002 3544 114008 3596
rect 114060 3584 114066 3596
rect 114462 3584 114468 3596
rect 114060 3556 114468 3584
rect 114060 3544 114066 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 115198 3544 115204 3596
rect 115256 3584 115262 3596
rect 115842 3584 115848 3596
rect 115256 3556 115848 3584
rect 115256 3544 115262 3556
rect 115842 3544 115848 3556
rect 115900 3544 115906 3596
rect 116394 3544 116400 3596
rect 116452 3584 116458 3596
rect 117222 3584 117228 3596
rect 116452 3556 117228 3584
rect 116452 3544 116458 3556
rect 117222 3544 117228 3556
rect 117280 3544 117286 3596
rect 117590 3544 117596 3596
rect 117648 3584 117654 3596
rect 118602 3584 118608 3596
rect 117648 3556 118608 3584
rect 117648 3544 117654 3556
rect 118602 3544 118608 3556
rect 118660 3544 118666 3596
rect 122282 3544 122288 3596
rect 122340 3584 122346 3596
rect 122742 3584 122748 3596
rect 122340 3556 122748 3584
rect 122340 3544 122346 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 126238 3584 126244 3596
rect 123404 3556 126244 3584
rect 123404 3516 123432 3556
rect 126238 3544 126244 3556
rect 126296 3544 126302 3596
rect 103486 3488 123432 3516
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 128262 3476 128268 3528
rect 128320 3516 128326 3528
rect 129366 3516 129372 3528
rect 128320 3488 129372 3516
rect 128320 3476 128326 3488
rect 129366 3476 129372 3488
rect 129424 3476 129430 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 147582 3516 147588 3528
rect 147180 3488 147588 3516
rect 147180 3476 147186 3488
rect 147582 3476 147588 3488
rect 147640 3476 147646 3528
rect 258810 3476 258816 3528
rect 258868 3516 258874 3528
rect 260650 3516 260656 3528
rect 258868 3488 260656 3516
rect 258868 3476 258874 3488
rect 260650 3476 260656 3488
rect 260708 3476 260714 3528
rect 269114 3476 269120 3528
rect 269172 3516 269178 3528
rect 272426 3516 272432 3528
rect 269172 3488 272432 3516
rect 269172 3476 269178 3488
rect 272426 3476 272432 3488
rect 272484 3476 272490 3528
rect 281442 3476 281448 3528
rect 281500 3516 281506 3528
rect 286594 3516 286600 3528
rect 281500 3488 286600 3516
rect 281500 3476 281506 3488
rect 286594 3476 286600 3488
rect 286652 3476 286658 3528
rect 291930 3476 291936 3528
rect 291988 3516 291994 3528
rect 294874 3516 294880 3528
rect 291988 3488 294880 3516
rect 291988 3476 291994 3488
rect 294874 3476 294880 3488
rect 294932 3476 294938 3528
rect 301498 3476 301504 3528
rect 301556 3516 301562 3528
rect 303154 3516 303160 3528
rect 301556 3488 303160 3516
rect 301556 3476 301562 3488
rect 303154 3476 303160 3488
rect 303212 3476 303218 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 327074 3476 327080 3528
rect 327132 3516 327138 3528
rect 327994 3516 328000 3528
rect 327132 3488 328000 3516
rect 327132 3476 327138 3488
rect 327994 3476 328000 3488
rect 328052 3476 328058 3528
rect 340138 3476 340144 3528
rect 340196 3516 340202 3528
rect 342162 3516 342168 3528
rect 340196 3488 342168 3516
rect 340196 3476 340202 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 583110 3516 583116 3528
rect 582248 3488 583116 3516
rect 582248 3476 582254 3488
rect 583110 3476 583116 3488
rect 583168 3476 583174 3528
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 43438 3448 43444 3460
rect 15988 3420 43444 3448
rect 15988 3408 15994 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 63218 3408 63224 3460
rect 63276 3448 63282 3460
rect 75178 3448 75184 3460
rect 63276 3420 75184 3448
rect 63276 3408 63282 3420
rect 75178 3408 75184 3420
rect 75236 3408 75242 3460
rect 77386 3408 77392 3460
rect 77444 3448 77450 3460
rect 90266 3448 90272 3460
rect 77444 3420 90272 3448
rect 77444 3408 77450 3420
rect 90266 3408 90272 3420
rect 90324 3408 90330 3460
rect 91554 3408 91560 3460
rect 91612 3448 91618 3460
rect 104342 3448 104348 3460
rect 91612 3420 104348 3448
rect 91612 3408 91618 3420
rect 104342 3408 104348 3420
rect 104400 3408 104406 3460
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 106182 3448 106188 3460
rect 105780 3420 106188 3448
rect 105780 3408 105786 3420
rect 106182 3408 106188 3420
rect 106240 3408 106246 3460
rect 106918 3408 106924 3460
rect 106976 3448 106982 3460
rect 107562 3448 107568 3460
rect 106976 3420 107568 3448
rect 106976 3408 106982 3420
rect 107562 3408 107568 3420
rect 107620 3408 107626 3460
rect 109310 3408 109316 3460
rect 109368 3448 109374 3460
rect 110322 3448 110328 3460
rect 109368 3420 110328 3448
rect 109368 3408 109374 3420
rect 110322 3408 110328 3420
rect 110380 3408 110386 3460
rect 110506 3408 110512 3460
rect 110564 3448 110570 3460
rect 111702 3448 111708 3460
rect 110564 3420 111708 3448
rect 110564 3408 110570 3420
rect 111702 3408 111708 3420
rect 111760 3408 111766 3460
rect 137278 3448 137284 3460
rect 113146 3420 137284 3448
rect 108114 3340 108120 3392
rect 108172 3380 108178 3392
rect 113146 3380 113174 3420
rect 137278 3408 137284 3420
rect 137336 3408 137342 3460
rect 220078 3408 220084 3460
rect 220136 3448 220142 3460
rect 242894 3448 242900 3460
rect 220136 3420 242900 3448
rect 220136 3408 220142 3420
rect 242894 3408 242900 3420
rect 242952 3408 242958 3460
rect 260098 3408 260104 3460
rect 260156 3448 260162 3460
rect 267734 3448 267740 3460
rect 260156 3420 267740 3448
rect 260156 3408 260162 3420
rect 267734 3408 267740 3420
rect 267792 3408 267798 3460
rect 304258 3408 304264 3460
rect 304316 3448 304322 3460
rect 310238 3448 310244 3460
rect 304316 3420 310244 3448
rect 304316 3408 304322 3420
rect 310238 3408 310244 3420
rect 310296 3408 310302 3460
rect 327718 3408 327724 3460
rect 327776 3448 327782 3460
rect 329190 3448 329196 3460
rect 327776 3420 329196 3448
rect 327776 3408 327782 3420
rect 329190 3408 329196 3420
rect 329248 3408 329254 3460
rect 341518 3408 341524 3460
rect 341576 3448 341582 3460
rect 350442 3448 350448 3460
rect 341576 3420 350448 3448
rect 341576 3408 341582 3420
rect 350442 3408 350448 3420
rect 350500 3408 350506 3460
rect 108172 3352 113174 3380
rect 108172 3340 108178 3352
rect 287698 3340 287704 3392
rect 287756 3380 287762 3392
rect 290182 3380 290188 3392
rect 287756 3352 290188 3380
rect 287756 3340 287762 3352
rect 290182 3340 290188 3352
rect 290240 3340 290246 3392
rect 20622 3272 20628 3324
rect 20680 3312 20686 3324
rect 25498 3312 25504 3324
rect 20680 3284 25504 3312
rect 20680 3272 20686 3284
rect 25498 3272 25504 3284
rect 25556 3272 25562 3324
rect 249794 3272 249800 3324
rect 249852 3312 249858 3324
rect 251174 3312 251180 3324
rect 249852 3284 251180 3312
rect 249852 3272 249858 3284
rect 251174 3272 251180 3284
rect 251232 3272 251238 3324
rect 298738 3272 298744 3324
rect 298796 3312 298802 3324
rect 301958 3312 301964 3324
rect 298796 3284 301964 3312
rect 298796 3272 298802 3284
rect 301958 3272 301964 3284
rect 302016 3272 302022 3324
rect 317322 3272 317328 3324
rect 317380 3312 317386 3324
rect 321646 3312 321652 3324
rect 317380 3284 321652 3312
rect 317380 3272 317386 3284
rect 321646 3272 321652 3284
rect 321704 3272 321710 3324
rect 76190 3204 76196 3256
rect 76248 3244 76254 3256
rect 77202 3244 77208 3256
rect 76248 3216 77208 3244
rect 76248 3204 76254 3216
rect 77202 3204 77208 3216
rect 77260 3204 77266 3256
rect 289078 3204 289084 3256
rect 289136 3244 289142 3256
rect 292574 3244 292580 3256
rect 289136 3216 292580 3244
rect 289136 3204 289142 3216
rect 292574 3204 292580 3216
rect 292632 3204 292638 3256
rect 349246 3136 349252 3188
rect 349304 3176 349310 3188
rect 351914 3176 351920 3188
rect 349304 3148 351920 3176
rect 349304 3136 349310 3148
rect 351914 3136 351920 3148
rect 351972 3136 351978 3188
rect 299658 3068 299664 3120
rect 299716 3108 299722 3120
rect 302234 3108 302240 3120
rect 299716 3080 302240 3108
rect 299716 3068 299722 3080
rect 302234 3068 302240 3080
rect 302292 3068 302298 3120
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 15838 3040 15844 3052
rect 11204 3012 15844 3040
rect 11204 3000 11210 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 118786 3000 118792 3052
rect 118844 3040 118850 3052
rect 119798 3040 119804 3052
rect 118844 3012 119804 3040
rect 118844 3000 118850 3012
rect 119798 3000 119804 3012
rect 119856 3000 119862 3052
rect 309778 3000 309784 3052
rect 309836 3040 309842 3052
rect 315022 3040 315028 3052
rect 309836 3012 315028 3040
rect 309836 3000 309842 3012
rect 315022 3000 315028 3012
rect 315080 3000 315086 3052
rect 348050 3000 348056 3052
rect 348108 3040 348114 3052
rect 353294 3040 353300 3052
rect 348108 3012 353300 3040
rect 348108 3000 348114 3012
rect 353294 3000 353300 3012
rect 353352 3000 353358 3052
rect 580994 3000 581000 3052
rect 581052 3040 581058 3052
rect 582558 3040 582564 3052
rect 581052 3012 582564 3040
rect 581052 3000 581058 3012
rect 582558 3000 582564 3012
rect 582616 3000 582622 3052
rect 246298 2932 246304 2984
rect 246356 2972 246362 2984
rect 247586 2972 247592 2984
rect 246356 2944 247592 2972
rect 246356 2932 246362 2944
rect 247586 2932 247592 2944
rect 247644 2932 247650 2984
rect 282178 2932 282184 2984
rect 282236 2972 282242 2984
rect 283098 2972 283104 2984
rect 282236 2944 283104 2972
rect 282236 2932 282242 2944
rect 283098 2932 283104 2944
rect 283156 2932 283162 2984
rect 299474 2184 299480 2236
rect 299532 2224 299538 2236
rect 300762 2224 300768 2236
rect 299532 2196 300768 2224
rect 299532 2184 299538 2196
rect 300762 2184 300768 2196
rect 300820 2184 300826 2236
rect 51350 2116 51356 2168
rect 51408 2156 51414 2168
rect 79318 2156 79324 2168
rect 51408 2128 79324 2156
rect 51408 2116 51414 2128
rect 79318 2116 79324 2128
rect 79376 2116 79382 2168
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 65426 2088 65432 2100
rect 7708 2060 65432 2088
rect 7708 2048 7714 2060
rect 65426 2048 65432 2060
rect 65484 2048 65490 2100
rect 140038 2048 140044 2100
rect 140096 2088 140102 2100
rect 160738 2088 160744 2100
rect 140096 2060 160744 2088
rect 140096 2048 140102 2060
rect 160738 2048 160744 2060
rect 160796 2048 160802 2100
rect 226978 2048 226984 2100
rect 227036 2088 227042 2100
rect 280706 2088 280712 2100
rect 227036 2060 280712 2088
rect 227036 2048 227042 2060
rect 280706 2048 280712 2060
rect 280764 2048 280770 2100
<< via1 >>
rect 191748 703400 191800 703452
rect 283840 703400 283892 703452
rect 282828 703332 282880 703384
rect 348792 703332 348844 703384
rect 214564 703264 214616 703316
rect 364984 703264 365036 703316
rect 240784 703196 240836 703248
rect 332508 703196 332560 703248
rect 249064 703128 249116 703180
rect 413652 703128 413704 703180
rect 273904 703060 273956 703112
rect 462320 703060 462372 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 102048 702992 102100 703044
rect 300124 702992 300176 703044
rect 271144 702924 271196 702976
rect 478512 702924 478564 702976
rect 8116 702856 8168 702908
rect 96620 702856 96672 702908
rect 213184 702856 213236 702908
rect 429844 702856 429896 702908
rect 24308 702788 24360 702840
rect 86224 702788 86276 702840
rect 177304 702788 177356 702840
rect 397460 702788 397512 702840
rect 69664 702720 69716 702772
rect 154120 702720 154172 702772
rect 280804 702720 280856 702772
rect 543464 702720 543516 702772
rect 90364 702652 90416 702704
rect 235172 702652 235224 702704
rect 258724 702652 258776 702704
rect 559656 702652 559708 702704
rect 84108 702584 84160 702636
rect 202788 702584 202840 702636
rect 215944 702584 215996 702636
rect 527088 702584 527140 702636
rect 67640 702516 67692 702568
rect 170312 702516 170364 702568
rect 184848 702516 184900 702568
rect 580908 702516 580960 702568
rect 79968 702448 80020 702500
rect 494796 702448 494848 702500
rect 71688 700272 71740 700324
rect 105452 700272 105504 700324
rect 220084 700272 220136 700324
rect 267648 700272 267700 700324
rect 218980 698912 219032 698964
rect 241520 698912 241572 698964
rect 3424 683136 3476 683188
rect 11704 683136 11756 683188
rect 3516 670692 3568 670744
rect 14464 670692 14516 670744
rect 3424 656888 3476 656940
rect 74540 656888 74592 656940
rect 3516 618604 3568 618656
rect 7564 618604 7616 618656
rect 3516 605820 3568 605872
rect 93124 605820 93176 605872
rect 81440 592628 81492 592680
rect 84108 592628 84160 592680
rect 143540 592628 143592 592680
rect 79324 589840 79376 589892
rect 79968 589840 80020 589892
rect 79968 589296 80020 589348
rect 124220 589296 124272 589348
rect 67548 588548 67600 588600
rect 71688 588548 71740 588600
rect 128360 588548 128412 588600
rect 40040 587120 40092 587172
rect 96712 587120 96764 587172
rect 82728 586508 82780 586560
rect 123484 586508 123536 586560
rect 78128 585760 78180 585812
rect 88340 585760 88392 585812
rect 112444 585760 112496 585812
rect 121736 585760 121788 585812
rect 582748 585760 582800 585812
rect 52368 585148 52420 585200
rect 84292 585148 84344 585200
rect 87512 585148 87564 585200
rect 121460 585148 121512 585200
rect 121736 585148 121788 585200
rect 93124 584400 93176 584452
rect 97264 584400 97316 584452
rect 76288 583720 76340 583772
rect 108304 583720 108356 583772
rect 77208 582768 77260 582820
rect 79324 582768 79376 582820
rect 86224 582496 86276 582548
rect 106924 582496 106976 582548
rect 79048 582428 79100 582480
rect 86868 582428 86920 582480
rect 50988 582360 51040 582412
rect 69940 582360 69992 582412
rect 73528 582360 73580 582412
rect 95884 582360 95936 582412
rect 62028 581068 62080 581120
rect 90548 581068 90600 581120
rect 60648 581000 60700 581052
rect 69020 581000 69072 581052
rect 3148 580932 3200 580984
rect 80244 581000 80296 581052
rect 90272 581000 90324 581052
rect 104256 581000 104308 581052
rect 86868 580660 86920 580712
rect 93768 580660 93820 580712
rect 102784 580252 102836 580304
rect 141424 579640 141476 579692
rect 97172 578212 97224 578264
rect 134524 578212 134576 578264
rect 98000 576852 98052 576904
rect 132592 576852 132644 576904
rect 3424 576784 3476 576836
rect 67732 576784 67784 576836
rect 97908 576716 97960 576768
rect 102048 576716 102100 576768
rect 102048 576104 102100 576156
rect 125600 576104 125652 576156
rect 94688 573316 94740 573368
rect 126980 573316 127032 573368
rect 96988 572704 97040 572756
rect 100852 572704 100904 572756
rect 53656 571344 53708 571396
rect 66812 571344 66864 571396
rect 97540 571344 97592 571396
rect 99380 571344 99432 571396
rect 97264 570664 97316 570716
rect 98736 570664 98788 570716
rect 55036 570596 55088 570648
rect 66720 570596 66772 570648
rect 59268 569984 59320 570036
rect 66904 569984 66956 570036
rect 97908 569916 97960 569968
rect 109684 569916 109736 569968
rect 64696 568556 64748 568608
rect 66536 568556 66588 568608
rect 95884 567808 95936 567860
rect 111064 567808 111116 567860
rect 57704 565836 57756 565888
rect 67640 565836 67692 565888
rect 56508 564408 56560 564460
rect 66904 564408 66956 564460
rect 52276 563048 52328 563100
rect 66904 563048 66956 563100
rect 96804 561688 96856 561740
rect 113180 561688 113232 561740
rect 48136 560260 48188 560312
rect 66812 560260 66864 560312
rect 96804 560260 96856 560312
rect 117320 560260 117372 560312
rect 97080 558968 97132 559020
rect 100024 558968 100076 559020
rect 57888 558900 57940 558952
rect 66812 558900 66864 558952
rect 97908 558152 97960 558204
rect 122840 558152 122892 558204
rect 61936 557540 61988 557592
rect 66812 557540 66864 557592
rect 96620 556928 96672 556980
rect 97080 556928 97132 556980
rect 96712 554752 96764 554804
rect 129004 554752 129056 554804
rect 2780 553800 2832 553852
rect 4804 553800 4856 553852
rect 63316 553392 63368 553444
rect 66904 553392 66956 553444
rect 96988 552032 97040 552084
rect 112536 552032 112588 552084
rect 96620 551828 96672 551880
rect 96896 551828 96948 551880
rect 97448 549312 97500 549364
rect 100760 549312 100812 549364
rect 53748 549244 53800 549296
rect 66720 549244 66772 549296
rect 55128 546456 55180 546508
rect 66812 546456 66864 546508
rect 59176 545096 59228 545148
rect 66812 545096 66864 545148
rect 97080 543736 97132 543788
rect 108396 543736 108448 543788
rect 11704 543668 11756 543720
rect 67640 543668 67692 543720
rect 68376 543668 68428 543720
rect 97080 542376 97132 542428
rect 125692 542376 125744 542428
rect 14464 541628 14516 541680
rect 42800 541628 42852 541680
rect 42800 540948 42852 541000
rect 43996 540948 44048 541000
rect 66628 540948 66680 541000
rect 96620 540948 96672 541000
rect 130384 540948 130436 541000
rect 3424 540200 3476 540252
rect 69388 539792 69440 539844
rect 91008 539792 91060 539844
rect 96804 539792 96856 539844
rect 70308 539656 70360 539708
rect 76564 539656 76616 539708
rect 86592 539588 86644 539640
rect 94320 539588 94372 539640
rect 67272 539044 67324 539096
rect 71872 539044 71924 539096
rect 11704 538228 11756 538280
rect 93952 538228 94004 538280
rect 4804 538160 4856 538212
rect 70676 538160 70728 538212
rect 70676 536800 70728 536852
rect 71044 536800 71096 536852
rect 7564 536732 7616 536784
rect 73528 536732 73580 536784
rect 68928 536120 68980 536172
rect 80704 536120 80756 536172
rect 82820 536120 82872 536172
rect 87604 536120 87656 536172
rect 93400 536120 93452 536172
rect 98644 536120 98696 536172
rect 73528 536052 73580 536104
rect 77944 536052 77996 536104
rect 80060 536052 80112 536104
rect 93124 536052 93176 536104
rect 88984 535440 89036 535492
rect 91100 535440 91152 535492
rect 67824 534692 67876 534744
rect 83464 534692 83516 534744
rect 48228 533332 48280 533384
rect 76748 533332 76800 533384
rect 78312 533332 78364 533384
rect 111156 533332 111208 533384
rect 64788 531972 64840 532024
rect 96896 531972 96948 532024
rect 67364 530612 67416 530664
rect 147680 530612 147732 530664
rect 3516 530544 3568 530596
rect 98000 530544 98052 530596
rect 50896 529184 50948 529236
rect 84200 529184 84252 529236
rect 64696 527824 64748 527876
rect 115940 527824 115992 527876
rect 3424 526396 3476 526448
rect 94504 526396 94556 526448
rect 95148 525784 95200 525836
rect 95424 525784 95476 525836
rect 71780 525036 71832 525088
rect 136732 525036 136784 525088
rect 85672 522384 85724 522436
rect 105544 522384 105596 522436
rect 61936 522248 61988 522300
rect 85672 522248 85724 522300
rect 59084 518168 59136 518220
rect 100852 518168 100904 518220
rect 3516 514768 3568 514820
rect 21364 514768 21416 514820
rect 71044 497428 71096 497480
rect 120724 497428 120776 497480
rect 85580 494708 85632 494760
rect 118792 494708 118844 494760
rect 73160 493280 73212 493332
rect 133880 493280 133932 493332
rect 65984 490560 66036 490612
rect 92572 490560 92624 490612
rect 77944 487772 77996 487824
rect 102876 487772 102928 487824
rect 80704 486412 80756 486464
rect 99472 486412 99524 486464
rect 188988 484372 189040 484424
rect 580172 484372 580224 484424
rect 67824 484304 67876 484356
rect 69020 484304 69072 484356
rect 106924 483624 106976 483676
rect 131120 483624 131172 483676
rect 77300 482264 77352 482316
rect 88984 482264 89036 482316
rect 258172 481584 258224 481636
rect 258724 481584 258776 481636
rect 93124 480904 93176 480956
rect 121552 480904 121604 480956
rect 122748 480224 122800 480276
rect 258172 480224 258224 480276
rect 110420 478864 110472 478916
rect 111064 478864 111116 478916
rect 251824 478864 251876 478916
rect 98736 478116 98788 478168
rect 124312 478116 124364 478168
rect 48136 477504 48188 477556
rect 202144 477504 202196 477556
rect 85580 476756 85632 476808
rect 95240 476756 95292 476808
rect 8208 476076 8260 476128
rect 11704 476076 11756 476128
rect 109776 476076 109828 476128
rect 249064 476076 249116 476128
rect 59176 476008 59228 476060
rect 122748 476008 122800 476060
rect 123024 476008 123076 476060
rect 3424 475192 3476 475244
rect 7564 475192 7616 475244
rect 8208 475192 8260 475244
rect 104256 474716 104308 474768
rect 238024 474716 238076 474768
rect 90916 473356 90968 473408
rect 226984 473356 227036 473408
rect 94504 473288 94556 473340
rect 95056 473288 95108 473340
rect 202880 472064 202932 472116
rect 295340 472064 295392 472116
rect 95056 471996 95108 472048
rect 231860 471996 231912 472048
rect 240140 471928 240192 471980
rect 240784 471928 240836 471980
rect 102140 471248 102192 471300
rect 102784 471248 102836 471300
rect 240140 471248 240192 471300
rect 155776 470568 155828 470620
rect 251180 470568 251232 470620
rect 70308 469820 70360 469872
rect 91192 469820 91244 469872
rect 105544 469820 105596 469872
rect 241520 469820 241572 469872
rect 241520 469276 241572 469328
rect 242164 469276 242216 469328
rect 85488 469208 85540 469260
rect 86224 469208 86276 469260
rect 104900 469208 104952 469260
rect 105544 469208 105596 469260
rect 123484 469208 123536 469260
rect 255412 469208 255464 469260
rect 111156 468460 111208 468512
rect 117780 468460 117832 468512
rect 93860 467848 93912 467900
rect 95148 467848 95200 467900
rect 227812 467916 227864 467968
rect 117412 467848 117464 467900
rect 117780 467848 117832 467900
rect 258264 467848 258316 467900
rect 164148 466488 164200 466540
rect 242900 466488 242952 466540
rect 112536 466420 112588 466472
rect 142068 466420 142120 466472
rect 252560 466420 252612 466472
rect 170496 465128 170548 465180
rect 259552 465128 259604 465180
rect 142804 465060 142856 465112
rect 245660 465060 245712 465112
rect 119344 463768 119396 463820
rect 255320 463768 255372 463820
rect 115204 463700 115256 463752
rect 262220 463700 262272 463752
rect 212632 463632 212684 463684
rect 213184 463632 213236 463684
rect 67640 463020 67692 463072
rect 81348 463020 81400 463072
rect 80060 462952 80112 463004
rect 113272 462952 113324 463004
rect 184204 462408 184256 462460
rect 212632 462408 212684 462460
rect 3240 462340 3292 462392
rect 11704 462340 11756 462392
rect 64788 462340 64840 462392
rect 186964 462340 187016 462392
rect 187056 462340 187108 462392
rect 260840 462340 260892 462392
rect 215392 462272 215444 462324
rect 215944 462272 215996 462324
rect 78680 461592 78732 461644
rect 91744 461592 91796 461644
rect 286324 461592 286376 461644
rect 583300 461592 583352 461644
rect 201500 461320 201552 461372
rect 202144 461320 202196 461372
rect 182824 460980 182876 461032
rect 215392 460980 215444 461032
rect 62028 460912 62080 460964
rect 185584 460912 185636 460964
rect 202144 460912 202196 460964
rect 286324 460912 286376 460964
rect 87604 460844 87656 460896
rect 109040 460844 109092 460896
rect 109040 460164 109092 460216
rect 109776 460164 109828 460216
rect 141424 459620 141476 459672
rect 256792 459620 256844 459672
rect 81348 459552 81400 459604
rect 208400 459552 208452 459604
rect 226984 459552 227036 459604
rect 227628 459552 227680 459604
rect 258356 459552 258408 459604
rect 77208 458804 77260 458856
rect 90364 458804 90416 458856
rect 95240 458260 95292 458312
rect 195796 458260 195848 458312
rect 227720 458260 227772 458312
rect 237380 458260 237432 458312
rect 291200 458260 291252 458312
rect 111708 458192 111760 458244
rect 259460 458192 259512 458244
rect 193404 456832 193456 456884
rect 218980 456832 219032 456884
rect 78680 456764 78732 456816
rect 173624 456764 173676 456816
rect 173808 456764 173860 456816
rect 179328 456764 179380 456816
rect 204536 456764 204588 456816
rect 230480 456764 230532 456816
rect 287152 456764 287204 456816
rect 580172 456764 580224 456816
rect 251180 456084 251232 456136
rect 252100 456084 252152 456136
rect 238024 456016 238076 456068
rect 241520 456016 241572 456068
rect 72424 455472 72476 455524
rect 160100 455472 160152 455524
rect 197360 455472 197412 455524
rect 225512 455472 225564 455524
rect 261484 455472 261536 455524
rect 98000 455404 98052 455456
rect 233240 455404 233292 455456
rect 82820 455336 82872 455388
rect 111708 455336 111760 455388
rect 112720 455336 112772 455388
rect 191196 454112 191248 454164
rect 218152 454112 218204 454164
rect 76564 454044 76616 454096
rect 159456 454044 159508 454096
rect 200120 454044 200172 454096
rect 222568 454044 222620 454096
rect 267004 454044 267056 454096
rect 227628 453976 227680 454028
rect 228732 453976 228784 454028
rect 212724 453364 212776 453416
rect 215484 453364 215536 453416
rect 195980 453296 196032 453348
rect 212448 453296 212500 453348
rect 193312 452752 193364 452804
rect 213644 452752 213696 452804
rect 251824 452752 251876 452804
rect 268384 452752 268436 452804
rect 222108 452684 222160 452736
rect 251456 452684 251508 452736
rect 60464 452616 60516 452668
rect 170404 452616 170456 452668
rect 192484 452616 192536 452668
rect 196532 452616 196584 452668
rect 211252 452616 211304 452668
rect 226892 452616 226944 452668
rect 227720 452616 227772 452668
rect 229652 452616 229704 452668
rect 237380 452616 237432 452668
rect 274640 452616 274692 452668
rect 82728 451936 82780 451988
rect 122840 451936 122892 451988
rect 124128 451936 124180 451988
rect 87604 451868 87656 451920
rect 187608 451868 187660 451920
rect 188344 451868 188396 451920
rect 240232 451392 240284 451444
rect 189816 451324 189868 451376
rect 241060 451324 241112 451376
rect 256700 451324 256752 451376
rect 191840 451256 191892 451308
rect 199292 451256 199344 451308
rect 210424 451256 210476 451308
rect 583300 451256 583352 451308
rect 101404 450508 101456 450560
rect 117964 450508 118016 450560
rect 192576 450508 192628 450560
rect 211252 450508 211304 450560
rect 231860 449964 231912 450016
rect 232872 449964 232924 450016
rect 267740 449964 267792 450016
rect 59268 449896 59320 449948
rect 151084 449896 151136 449948
rect 178684 449896 178736 449948
rect 240232 449896 240284 449948
rect 242440 449896 242492 449948
rect 254584 449896 254636 449948
rect 73804 449828 73856 449880
rect 200948 449828 201000 449880
rect 3240 449760 3292 449812
rect 100760 449760 100812 449812
rect 251456 449692 251508 449744
rect 173808 449148 173860 449200
rect 193404 449148 193456 449200
rect 255504 449216 255556 449268
rect 271236 449216 271288 449268
rect 269120 449148 269172 449200
rect 64696 448536 64748 448588
rect 74540 448536 74592 448588
rect 75828 448536 75880 448588
rect 53656 447856 53708 447908
rect 106924 447856 106976 447908
rect 112444 447856 112496 447908
rect 122932 447856 122984 447908
rect 169024 447856 169076 447908
rect 191656 447856 191708 447908
rect 75828 447788 75880 447840
rect 181444 447788 181496 447840
rect 255412 447788 255464 447840
rect 287060 447788 287112 447840
rect 188436 447108 188488 447160
rect 191012 447108 191064 447160
rect 176568 446360 176620 446412
rect 191840 446360 191892 446412
rect 59176 445816 59228 445868
rect 152464 445816 152516 445868
rect 71136 445748 71188 445800
rect 191656 445748 191708 445800
rect 186320 445680 186372 445732
rect 187608 445680 187660 445732
rect 191196 445680 191248 445732
rect 52276 445000 52328 445052
rect 60556 445000 60608 445052
rect 88248 445000 88300 445052
rect 91008 445000 91060 445052
rect 186320 445000 186372 445052
rect 60556 444388 60608 444440
rect 88524 444388 88576 444440
rect 255412 444388 255464 444440
rect 263784 444388 263836 444440
rect 111892 444320 111944 444372
rect 112536 444320 112588 444372
rect 107660 443776 107712 443828
rect 108396 443776 108448 443828
rect 142804 443640 142856 443692
rect 65984 443504 66036 443556
rect 70492 443504 70544 443556
rect 255412 443368 255464 443420
rect 259460 443368 259512 443420
rect 3424 442960 3476 443012
rect 111892 442960 111944 443012
rect 117320 442892 117372 442944
rect 117780 442892 117832 442944
rect 192484 442892 192536 442944
rect 70400 442212 70452 442264
rect 117780 442212 117832 442264
rect 125692 442076 125744 442128
rect 126244 442076 126296 442128
rect 255412 442008 255464 442060
rect 258172 442008 258224 442060
rect 258724 442008 258776 442060
rect 63224 441600 63276 441652
rect 125692 441600 125744 441652
rect 67088 440852 67140 440904
rect 122840 440852 122892 440904
rect 67364 440240 67416 440292
rect 166356 440240 166408 440292
rect 176660 440240 176712 440292
rect 191380 440240 191432 440292
rect 185768 439492 185820 439544
rect 193312 439492 193364 439544
rect 255320 439492 255372 439544
rect 288532 439492 288584 439544
rect 583024 439492 583076 439544
rect 44088 438948 44140 439000
rect 69664 438948 69716 439000
rect 83464 438948 83516 439000
rect 83740 438948 83792 439000
rect 185768 438948 185820 439000
rect 186136 438948 186188 439000
rect 68284 438880 68336 438932
rect 191380 438880 191432 438932
rect 65984 438132 66036 438184
rect 191564 438132 191616 438184
rect 255412 438132 255464 438184
rect 258264 438132 258316 438184
rect 266360 438132 266412 438184
rect 95056 437588 95108 437640
rect 96988 437588 97040 437640
rect 48136 437452 48188 437504
rect 50988 437452 51040 437504
rect 74816 437452 74868 437504
rect 71688 437384 71740 437436
rect 72424 437384 72476 437436
rect 82820 437384 82872 437436
rect 83924 437384 83976 437436
rect 87604 437384 87656 437436
rect 90916 437384 90968 437436
rect 94228 437384 94280 437436
rect 102876 437384 102928 437436
rect 178684 437384 178736 437436
rect 263416 437384 263468 437436
rect 582472 437384 582524 437436
rect 80980 437316 81032 437368
rect 86224 437316 86276 437368
rect 68928 437112 68980 437164
rect 69756 437112 69808 437164
rect 91744 436704 91796 436756
rect 104440 436704 104492 436756
rect 136640 436704 136692 436756
rect 189816 436704 189868 436756
rect 255412 436704 255464 436756
rect 262312 436704 262364 436756
rect 120724 436500 120776 436552
rect 122104 436500 122156 436552
rect 74080 436432 74132 436484
rect 76564 436432 76616 436484
rect 87328 436296 87380 436348
rect 88248 436296 88300 436348
rect 52184 436092 52236 436144
rect 68928 436092 68980 436144
rect 69664 436092 69716 436144
rect 71044 436092 71096 436144
rect 75828 436092 75880 436144
rect 80428 436092 80480 436144
rect 108304 436092 108356 436144
rect 120724 436092 120776 436144
rect 186964 436024 187016 436076
rect 191564 436024 191616 436076
rect 103888 435412 103940 435464
rect 104440 435412 104492 435464
rect 136640 435412 136692 435464
rect 67272 435344 67324 435396
rect 176660 435344 176712 435396
rect 255412 435344 255464 435396
rect 259644 435344 259696 435396
rect 271880 435344 271932 435396
rect 15844 434732 15896 434784
rect 70584 434732 70636 434784
rect 115756 434664 115808 434716
rect 180156 434664 180208 434716
rect 255412 434664 255464 434716
rect 262220 434664 262272 434716
rect 263692 434664 263744 434716
rect 57612 434052 57664 434104
rect 60648 434052 60700 434104
rect 66812 434052 66864 434104
rect 104164 433984 104216 434036
rect 115296 433984 115348 434036
rect 180708 433984 180760 434036
rect 191104 433984 191156 434036
rect 68376 433644 68428 433696
rect 71136 433644 71188 433696
rect 112352 433644 112404 433696
rect 114008 433644 114060 433696
rect 68652 433236 68704 433288
rect 188436 433236 188488 433288
rect 115848 433168 115900 433220
rect 123484 433168 123536 433220
rect 185584 433168 185636 433220
rect 190644 433168 190696 433220
rect 64604 431944 64656 431996
rect 67548 431944 67600 431996
rect 255412 431944 255464 431996
rect 262220 431944 262272 431996
rect 115848 431196 115900 431248
rect 118700 431196 118752 431248
rect 152464 431196 152516 431248
rect 191196 431196 191248 431248
rect 170404 430516 170456 430568
rect 191104 430516 191156 430568
rect 114008 429836 114060 429888
rect 143632 429836 143684 429888
rect 255504 429496 255556 429548
rect 259552 429496 259604 429548
rect 181444 429088 181496 429140
rect 191748 429088 191800 429140
rect 115848 428408 115900 428460
rect 122840 428408 122892 428460
rect 123024 428408 123076 428460
rect 255412 428408 255464 428460
rect 270592 428408 270644 428460
rect 67548 428340 67600 428392
rect 68284 428340 68336 428392
rect 255412 427796 255464 427848
rect 288440 427796 288492 427848
rect 255504 427728 255556 427780
rect 260840 427728 260892 427780
rect 262128 427728 262180 427780
rect 116584 427048 116636 427100
rect 162124 427048 162176 427100
rect 262128 427048 262180 427100
rect 285680 427048 285732 427100
rect 63408 426436 63460 426488
rect 66996 426436 67048 426488
rect 151084 426368 151136 426420
rect 170404 426368 170456 426420
rect 190644 426436 190696 426488
rect 285680 426436 285732 426488
rect 582656 426436 582708 426488
rect 115388 426232 115440 426284
rect 119344 426232 119396 426284
rect 57796 425688 57848 425740
rect 67272 425688 67324 425740
rect 126336 425688 126388 425740
rect 141424 425688 141476 425740
rect 174544 425688 174596 425740
rect 191748 425688 191800 425740
rect 255872 425688 255924 425740
rect 256792 425688 256844 425740
rect 269212 425688 269264 425740
rect 115020 425008 115072 425060
rect 117504 425008 117556 425060
rect 115388 424940 115440 424992
rect 117412 424940 117464 424992
rect 54944 423648 54996 423700
rect 66628 423648 66680 423700
rect 115020 423512 115072 423564
rect 120816 423512 120868 423564
rect 49608 422900 49660 422952
rect 64788 422900 64840 422952
rect 66812 422900 66864 422952
rect 126244 422900 126296 422952
rect 166264 422900 166316 422952
rect 166264 422288 166316 422340
rect 190644 422288 190696 422340
rect 255504 422288 255556 422340
rect 276112 422288 276164 422340
rect 62028 422220 62080 422272
rect 66628 422220 66680 422272
rect 52276 421540 52328 421592
rect 62028 421540 62080 421592
rect 255964 421540 256016 421592
rect 262864 421540 262916 421592
rect 115296 420928 115348 420980
rect 188436 420928 188488 420980
rect 255504 420928 255556 420980
rect 283012 420928 283064 420980
rect 60464 420860 60516 420912
rect 66812 420860 66864 420912
rect 64788 420248 64840 420300
rect 67088 420248 67140 420300
rect 115756 419500 115808 419552
rect 129832 419500 129884 419552
rect 171876 419500 171928 419552
rect 191748 419500 191800 419552
rect 255504 419500 255556 419552
rect 260840 419500 260892 419552
rect 59268 418752 59320 418804
rect 67640 418752 67692 418804
rect 123484 418752 123536 418804
rect 136732 418752 136784 418804
rect 187056 418752 187108 418804
rect 289728 418752 289780 418804
rect 583116 418752 583168 418804
rect 59176 418276 59228 418328
rect 66812 418276 66864 418328
rect 178684 418140 178736 418192
rect 191748 418140 191800 418192
rect 255412 418140 255464 418192
rect 288624 418140 288676 418192
rect 289728 418140 289780 418192
rect 64696 418072 64748 418124
rect 67088 418072 67140 418124
rect 112720 418072 112772 418124
rect 170496 418072 170548 418124
rect 265256 417460 265308 417512
rect 271144 417460 271196 417512
rect 162124 417392 162176 417444
rect 162768 417392 162820 417444
rect 191748 417392 191800 417444
rect 270408 417392 270460 417444
rect 583208 417392 583260 417444
rect 113916 417052 113968 417104
rect 117964 417052 118016 417104
rect 255412 416848 255464 416900
rect 265072 416848 265124 416900
rect 265256 416848 265308 416900
rect 255504 416780 255556 416832
rect 269304 416780 269356 416832
rect 270408 416780 270460 416832
rect 63316 416712 63368 416764
rect 66260 416712 66312 416764
rect 116124 416100 116176 416152
rect 126336 416100 126388 416152
rect 116584 416032 116636 416084
rect 142160 416032 142212 416084
rect 173164 416032 173216 416084
rect 187700 415896 187752 415948
rect 188988 415896 189040 415948
rect 190644 415896 190696 415948
rect 63224 415012 63276 415064
rect 66904 415012 66956 415064
rect 115848 414672 115900 414724
rect 125692 414672 125744 414724
rect 53656 413992 53708 414044
rect 66812 413992 66864 414044
rect 142160 413992 142212 414044
rect 191748 413992 191800 414044
rect 255412 413516 255464 413568
rect 258172 413516 258224 413568
rect 113180 412972 113232 413024
rect 117320 412972 117372 413024
rect 46848 412632 46900 412684
rect 66260 412632 66312 412684
rect 121644 412632 121696 412684
rect 148324 412632 148376 412684
rect 115848 412564 115900 412616
rect 123484 412564 123536 412616
rect 166356 411884 166408 411936
rect 166908 411884 166960 411936
rect 191748 411884 191800 411936
rect 39948 411272 40000 411324
rect 66260 411272 66312 411324
rect 50804 411204 50856 411256
rect 57704 411204 57756 411256
rect 66628 411204 66680 411256
rect 114744 410592 114796 410644
rect 116584 410592 116636 410644
rect 118700 410524 118752 410576
rect 131120 410524 131172 410576
rect 180156 410524 180208 410576
rect 3148 409844 3200 409896
rect 7656 409844 7708 409896
rect 188896 409844 188948 409896
rect 191012 409844 191064 409896
rect 255412 409844 255464 409896
rect 266452 409844 266504 409896
rect 125508 409096 125560 409148
rect 143540 409096 143592 409148
rect 187148 409096 187200 409148
rect 59084 408416 59136 408468
rect 62764 408484 62816 408536
rect 66812 408484 66864 408536
rect 115848 408484 115900 408536
rect 152464 408484 152516 408536
rect 186228 408484 186280 408536
rect 191012 408484 191064 408536
rect 255412 408484 255464 408536
rect 273352 408484 273404 408536
rect 130384 408416 130436 408468
rect 142160 408416 142212 408468
rect 115388 408348 115440 408400
rect 121644 408348 121696 408400
rect 48136 407124 48188 407176
rect 66904 407124 66956 407176
rect 53840 407056 53892 407108
rect 55036 407056 55088 407108
rect 66812 407056 66864 407108
rect 254584 407056 254636 407108
rect 259552 407056 259604 407108
rect 41236 406376 41288 406428
rect 53840 406376 53892 406428
rect 255412 406240 255464 406292
rect 259644 406240 259696 406292
rect 159364 405696 159416 405748
rect 191748 405696 191800 405748
rect 115848 405628 115900 405680
rect 125508 405628 125560 405680
rect 115756 405560 115808 405612
rect 118700 405560 118752 405612
rect 64696 404336 64748 404388
rect 66812 404336 66864 404388
rect 162124 404336 162176 404388
rect 191748 404336 191800 404388
rect 147680 403724 147732 403776
rect 148416 403724 148468 403776
rect 117228 403044 117280 403096
rect 147680 403044 147732 403096
rect 55036 402976 55088 403028
rect 66812 402976 66864 403028
rect 115848 402976 115900 403028
rect 155224 402976 155276 403028
rect 156604 402976 156656 403028
rect 191748 402976 191800 403028
rect 113456 402364 113508 402416
rect 118792 402364 118844 402416
rect 64604 401616 64656 401668
rect 66260 401616 66312 401668
rect 114744 401072 114796 401124
rect 117228 401072 117280 401124
rect 121644 400868 121696 400920
rect 128360 400868 128412 400920
rect 60648 400188 60700 400240
rect 66720 400188 66772 400240
rect 115572 400188 115624 400240
rect 119344 400188 119396 400240
rect 255412 400188 255464 400240
rect 277492 400188 277544 400240
rect 255412 399440 255464 399492
rect 258264 399440 258316 399492
rect 582840 399440 582892 399492
rect 115848 398828 115900 398880
rect 192668 398896 192720 398948
rect 184296 398828 184348 398880
rect 191748 398828 191800 398880
rect 4804 397468 4856 397520
rect 63316 397468 63368 397520
rect 67180 397468 67232 397520
rect 115388 397468 115440 397520
rect 118608 397468 118660 397520
rect 121644 397468 121696 397520
rect 159548 397468 159600 397520
rect 190828 397468 190880 397520
rect 115296 397128 115348 397180
rect 119436 397128 119488 397180
rect 53380 396720 53432 396772
rect 66812 396720 66864 396772
rect 160744 396720 160796 396772
rect 184848 396720 184900 396772
rect 191748 396720 191800 396772
rect 50896 395972 50948 396024
rect 67180 395972 67232 396024
rect 271236 395292 271288 395344
rect 287244 395292 287296 395344
rect 157984 394748 158036 394800
rect 190828 394748 190880 394800
rect 115848 394680 115900 394732
rect 189816 394680 189868 394732
rect 61844 393388 61896 393440
rect 67640 393388 67692 393440
rect 131764 393388 131816 393440
rect 132592 393388 132644 393440
rect 115756 393320 115808 393372
rect 151176 393320 151228 393372
rect 188528 393320 188580 393372
rect 190828 393320 190880 393372
rect 256884 393320 256936 393372
rect 271972 393320 272024 393372
rect 67364 393252 67416 393304
rect 67640 393252 67692 393304
rect 115572 392028 115624 392080
rect 116032 392028 116084 392080
rect 131764 392028 131816 392080
rect 184388 392028 184440 392080
rect 191564 392028 191616 392080
rect 56416 391960 56468 392012
rect 66812 391960 66864 392012
rect 115756 391960 115808 392012
rect 193404 391960 193456 392012
rect 267004 391212 267056 391264
rect 273444 391212 273496 391264
rect 114836 390736 114888 390788
rect 116584 390736 116636 390788
rect 111984 390600 112036 390652
rect 117228 390600 117280 390652
rect 67732 390532 67784 390584
rect 68652 390532 68704 390584
rect 73712 390532 73764 390584
rect 178040 390532 178092 390584
rect 196900 390600 196952 390652
rect 196072 390260 196124 390312
rect 247684 389784 247736 389836
rect 254032 389784 254084 389836
rect 109408 389240 109460 389292
rect 165620 389240 165672 389292
rect 248328 389240 248380 389292
rect 53748 389172 53800 389224
rect 83004 389172 83056 389224
rect 103152 389172 103204 389224
rect 238760 389172 238812 389224
rect 239956 389172 240008 389224
rect 249156 389172 249208 389224
rect 254216 389172 254268 389224
rect 11704 389104 11756 389156
rect 51448 389104 51500 389156
rect 52368 389104 52420 389156
rect 69664 389104 69716 389156
rect 73712 389104 73764 389156
rect 107844 389104 107896 389156
rect 246396 389104 246448 389156
rect 246580 389104 246632 389156
rect 48228 389036 48280 389088
rect 72516 389036 72568 389088
rect 111984 389036 112036 389088
rect 133880 389036 133932 389088
rect 251824 389036 251876 389088
rect 87604 387880 87656 387932
rect 92020 387880 92072 387932
rect 71136 387812 71188 387864
rect 71688 387812 71740 387864
rect 78128 387812 78180 387864
rect 78588 387812 78640 387864
rect 79968 387812 80020 387864
rect 81532 387812 81584 387864
rect 86224 387812 86276 387864
rect 87788 387812 87840 387864
rect 249248 387812 249300 387864
rect 251364 387812 251416 387864
rect 7564 387744 7616 387796
rect 93952 387744 94004 387796
rect 94504 387744 94556 387796
rect 100392 387744 100444 387796
rect 121552 387744 121604 387796
rect 122196 387744 122248 387796
rect 186044 387132 186096 387184
rect 221004 387132 221056 387184
rect 110420 387064 110472 387116
rect 186964 387064 187016 387116
rect 192668 387064 192720 387116
rect 214012 387064 214064 387116
rect 253480 387064 253532 387116
rect 226340 386996 226392 387048
rect 227260 386996 227312 387048
rect 231216 386384 231268 386436
rect 270500 386384 270552 386436
rect 43996 386316 44048 386368
rect 89260 386316 89312 386368
rect 99656 386316 99708 386368
rect 100852 386316 100904 386368
rect 105176 386316 105228 386368
rect 124312 386316 124364 386368
rect 124864 386316 124916 386368
rect 131764 386316 131816 386368
rect 256884 386316 256936 386368
rect 240784 386248 240836 386300
rect 247040 386248 247092 386300
rect 82084 385636 82136 385688
rect 91100 385636 91152 385688
rect 101956 385636 102008 385688
rect 112720 385636 112772 385688
rect 198004 385636 198056 385688
rect 203892 385636 203944 385688
rect 232504 385024 232556 385076
rect 239036 385024 239088 385076
rect 289912 385024 289964 385076
rect 582564 385024 582616 385076
rect 56508 384956 56560 385008
rect 86224 384956 86276 385008
rect 100944 384956 100996 385008
rect 236644 384956 236696 385008
rect 66168 384888 66220 384940
rect 87604 384888 87656 384940
rect 89168 384888 89220 384940
rect 126888 384888 126940 384940
rect 148324 384888 148376 384940
rect 148968 384888 149020 384940
rect 258172 384888 258224 384940
rect 236644 384276 236696 384328
rect 266544 384276 266596 384328
rect 279424 384276 279476 384328
rect 582932 384276 582984 384328
rect 189816 383596 189868 383648
rect 252744 383596 252796 383648
rect 255320 383596 255372 383648
rect 97908 382916 97960 382968
rect 128360 382916 128412 382968
rect 251824 382916 251876 382968
rect 267832 382916 267884 382968
rect 3516 382236 3568 382288
rect 113180 382236 113232 382288
rect 113456 382236 113508 382288
rect 128360 382236 128412 382288
rect 231860 382236 231912 382288
rect 252744 382236 252796 382288
rect 101036 382168 101088 382220
rect 122104 382168 122156 382220
rect 126888 382168 126940 382220
rect 186044 382168 186096 382220
rect 251824 382168 251876 382220
rect 187516 381556 187568 381608
rect 194600 381556 194652 381608
rect 101404 381488 101456 381540
rect 113548 381488 113600 381540
rect 191748 381488 191800 381540
rect 264980 381488 265032 381540
rect 186044 380876 186096 380928
rect 186320 380876 186372 380928
rect 198740 380876 198792 380928
rect 276020 380876 276072 380928
rect 105544 380808 105596 380860
rect 231216 380808 231268 380860
rect 274732 380808 274784 380860
rect 582380 380808 582432 380860
rect 193404 380740 193456 380792
rect 255596 380740 255648 380792
rect 188988 380264 189040 380316
rect 192576 380264 192628 380316
rect 60556 380196 60608 380248
rect 77484 380196 77536 380248
rect 73160 380128 73212 380180
rect 168380 380128 168432 380180
rect 106004 379448 106056 379500
rect 243084 379448 243136 379500
rect 67548 379380 67600 379432
rect 155960 379380 156012 379432
rect 156604 379380 156656 379432
rect 173072 379380 173124 379432
rect 173716 379380 173768 379432
rect 207020 379380 207072 379432
rect 243084 378972 243136 379024
rect 243544 378972 243596 379024
rect 231860 378768 231912 378820
rect 281724 378768 281776 378820
rect 106924 377476 106976 377528
rect 116032 377476 116084 377528
rect 78588 377408 78640 377460
rect 176476 377408 176528 377460
rect 205640 377408 205692 377460
rect 3424 376660 3476 376712
rect 116124 376660 116176 376712
rect 152464 376660 152516 376712
rect 247040 376660 247092 376712
rect 247684 376660 247736 376712
rect 92480 376592 92532 376644
rect 122932 376592 122984 376644
rect 123484 376592 123536 376644
rect 118608 375980 118660 376032
rect 277492 375980 277544 376032
rect 87604 375300 87656 375352
rect 88248 375300 88300 375352
rect 107476 375300 107528 375352
rect 245752 375300 245804 375352
rect 224960 375232 225012 375284
rect 255688 374620 255740 374672
rect 256792 374620 256844 374672
rect 291292 374620 291344 374672
rect 245752 374552 245804 374604
rect 246304 374552 246356 374604
rect 122196 373940 122248 373992
rect 236000 373940 236052 373992
rect 100576 373260 100628 373312
rect 118608 373260 118660 373312
rect 208492 373260 208544 373312
rect 284392 373260 284444 373312
rect 236000 372580 236052 372632
rect 236644 372580 236696 372632
rect 111800 372512 111852 372564
rect 112536 372512 112588 372564
rect 252652 372512 252704 372564
rect 75920 372444 75972 372496
rect 198004 372444 198056 372496
rect 209780 371832 209832 371884
rect 278872 371832 278924 371884
rect 114468 371152 114520 371204
rect 259644 371152 259696 371204
rect 260748 371152 260800 371204
rect 104164 370540 104216 370592
rect 113180 370540 113232 370592
rect 114468 370540 114520 370592
rect 94044 370472 94096 370524
rect 107660 370472 107712 370524
rect 155224 370472 155276 370524
rect 252468 370472 252520 370524
rect 255412 370472 255464 370524
rect 260748 370472 260800 370524
rect 281816 370472 281868 370524
rect 196072 369180 196124 369232
rect 240232 369180 240284 369232
rect 102140 369112 102192 369164
rect 137468 369112 137520 369164
rect 232504 369112 232556 369164
rect 130476 368432 130528 368484
rect 231124 368432 231176 368484
rect 89076 367820 89128 367872
rect 129004 367820 129056 367872
rect 232504 367820 232556 367872
rect 262220 367820 262272 367872
rect 74632 367752 74684 367804
rect 152556 367752 152608 367804
rect 201500 367752 201552 367804
rect 254584 367752 254636 367804
rect 582748 367752 582800 367804
rect 204260 367004 204312 367056
rect 582472 367004 582524 367056
rect 107752 366392 107804 366444
rect 180800 366392 180852 366444
rect 181352 366392 181404 366444
rect 45376 366324 45428 366376
rect 75920 366324 75972 366376
rect 82820 366324 82872 366376
rect 156604 366324 156656 366376
rect 213920 366324 213972 366376
rect 63316 365644 63368 365696
rect 184296 365644 184348 365696
rect 220728 365644 220780 365696
rect 240784 365644 240836 365696
rect 182916 364964 182968 365016
rect 229100 364964 229152 365016
rect 193404 363740 193456 363792
rect 195980 363740 196032 363792
rect 151176 363672 151228 363724
rect 253848 363740 253900 363792
rect 255504 363740 255556 363792
rect 71688 363604 71740 363656
rect 193404 363604 193456 363656
rect 116584 362856 116636 362908
rect 252560 362856 252612 362908
rect 86224 362788 86276 362840
rect 219532 362788 219584 362840
rect 220084 362788 220136 362840
rect 85580 361496 85632 361548
rect 216680 361496 216732 361548
rect 123484 361428 123536 361480
rect 226432 361428 226484 361480
rect 232596 360816 232648 360868
rect 263784 360816 263836 360868
rect 226432 360204 226484 360256
rect 226984 360204 227036 360256
rect 94504 359524 94556 359576
rect 124220 359524 124272 359576
rect 125048 359524 125100 359576
rect 56416 359456 56468 359508
rect 184388 359456 184440 359508
rect 215392 359456 215444 359508
rect 242900 359456 242952 359508
rect 125048 358776 125100 358828
rect 226340 358776 226392 358828
rect 84200 358708 84252 358760
rect 215300 358708 215352 358760
rect 215944 358708 215996 358760
rect 2780 358436 2832 358488
rect 4804 358436 4856 358488
rect 103520 357348 103572 357400
rect 240140 357348 240192 357400
rect 240784 357348 240836 357400
rect 226340 356668 226392 356720
rect 262220 356668 262272 356720
rect 129004 355988 129056 356040
rect 220912 355988 220964 356040
rect 221556 355988 221608 356040
rect 75736 355308 75788 355360
rect 193312 355308 193364 355360
rect 202880 355308 202932 355360
rect 79968 354628 80020 354680
rect 211160 354628 211212 354680
rect 81532 353948 81584 354000
rect 102140 353948 102192 354000
rect 212540 353948 212592 354000
rect 222200 353268 222252 353320
rect 231124 353268 231176 353320
rect 249708 353268 249760 353320
rect 252560 353268 252612 353320
rect 111064 353200 111116 353252
rect 249248 353200 249300 353252
rect 110512 352860 110564 352912
rect 111064 352860 111116 352912
rect 155868 352520 155920 352572
rect 194600 352520 194652 352572
rect 222844 352520 222896 352572
rect 95148 351840 95200 351892
rect 182180 351840 182232 351892
rect 182916 351840 182968 351892
rect 186964 351840 187016 351892
rect 187516 351840 187568 351892
rect 249800 351840 249852 351892
rect 195244 349868 195296 349920
rect 249156 349868 249208 349920
rect 154488 349800 154540 349852
rect 270592 349800 270644 349852
rect 196624 348372 196676 348424
rect 238024 348372 238076 348424
rect 67456 347760 67508 347812
rect 294052 347760 294104 347812
rect 123576 346468 123628 346520
rect 211160 346468 211212 346520
rect 211804 346468 211856 346520
rect 142988 346400 143040 346452
rect 234804 346400 234856 346452
rect 141608 345108 141660 345160
rect 234712 345108 234764 345160
rect 3332 345040 3384 345092
rect 11704 345040 11756 345092
rect 88984 345040 89036 345092
rect 292580 345040 292632 345092
rect 141424 343680 141476 343732
rect 142068 343680 142120 343732
rect 291384 343680 291436 343732
rect 37188 343612 37240 343664
rect 204260 343612 204312 343664
rect 172428 342864 172480 342916
rect 183468 342864 183520 342916
rect 224224 342864 224276 342916
rect 227720 342864 227772 342916
rect 253204 342864 253256 342916
rect 88248 342252 88300 342304
rect 233976 342252 234028 342304
rect 184756 341504 184808 341556
rect 208400 341504 208452 341556
rect 244372 341504 244424 341556
rect 263600 341504 263652 341556
rect 130476 340892 130528 340944
rect 244372 340892 244424 340944
rect 170956 340144 171008 340196
rect 244280 340144 244332 340196
rect 159548 339464 159600 339516
rect 295524 339464 295576 339516
rect 124864 338172 124916 338224
rect 229100 338172 229152 338224
rect 112444 338104 112496 338156
rect 238760 338104 238812 338156
rect 239404 338104 239456 338156
rect 184848 337424 184900 337476
rect 232596 337424 232648 337476
rect 223488 337356 223540 337408
rect 272064 337356 272116 337408
rect 42708 336744 42760 336796
rect 221464 336744 221516 336796
rect 190368 335996 190420 336048
rect 280252 335996 280304 336048
rect 108948 335724 109000 335776
rect 112536 335724 112588 335776
rect 155316 335316 155368 335368
rect 251824 335316 251876 335368
rect 184296 334568 184348 334620
rect 274732 334568 274784 334620
rect 145656 333956 145708 334008
rect 247040 333956 247092 334008
rect 247684 333956 247736 334008
rect 183468 333208 183520 333260
rect 232504 333208 232556 333260
rect 152648 332596 152700 332648
rect 233148 332596 233200 332648
rect 233884 332596 233936 332648
rect 174636 331304 174688 331356
rect 242900 331304 242952 331356
rect 173624 331236 173676 331288
rect 245660 331236 245712 331288
rect 246396 330488 246448 330540
rect 270592 330488 270644 330540
rect 177488 329876 177540 329928
rect 177948 329876 178000 329928
rect 232504 329876 232556 329928
rect 177304 329808 177356 329860
rect 240232 329808 240284 329860
rect 166356 329332 166408 329384
rect 166908 329332 166960 329384
rect 115204 329128 115256 329180
rect 115848 329128 115900 329180
rect 115848 328516 115900 328568
rect 192576 328516 192628 328568
rect 166356 328448 166408 328500
rect 256792 328448 256844 328500
rect 242808 328040 242860 328092
rect 244372 328040 244424 328092
rect 253848 327768 253900 327820
rect 265256 327768 265308 327820
rect 181996 327700 182048 327752
rect 192484 327700 192536 327752
rect 141700 327088 141752 327140
rect 189080 327088 189132 327140
rect 170404 326340 170456 326392
rect 184204 326340 184256 326392
rect 188344 326340 188396 326392
rect 227076 326340 227128 326392
rect 236644 326340 236696 326392
rect 259828 326340 259880 326392
rect 261484 326340 261536 326392
rect 283104 326340 283156 326392
rect 163596 325660 163648 325712
rect 242992 325660 243044 325712
rect 239404 324912 239456 324964
rect 249800 324912 249852 324964
rect 159364 324300 159416 324352
rect 259736 324300 259788 324352
rect 144276 323620 144328 323672
rect 159364 323620 159416 323672
rect 162400 323620 162452 323672
rect 259460 323620 259512 323672
rect 108396 323552 108448 323604
rect 120724 323552 120776 323604
rect 273536 323552 273588 323604
rect 125692 322872 125744 322924
rect 276112 322872 276164 322924
rect 104256 322260 104308 322312
rect 125692 322260 125744 322312
rect 86224 322192 86276 322244
rect 166264 322192 166316 322244
rect 258080 322192 258132 322244
rect 193128 320900 193180 320952
rect 216680 320900 216732 320952
rect 226984 320900 227036 320952
rect 262404 320900 262456 320952
rect 126888 320832 126940 320884
rect 136640 320832 136692 320884
rect 263600 320832 263652 320884
rect 268384 320832 268436 320884
rect 286416 320832 286468 320884
rect 104348 320220 104400 320272
rect 126888 320220 126940 320272
rect 75828 320152 75880 320204
rect 108304 320152 108356 320204
rect 175924 319472 175976 319524
rect 176568 319472 176620 319524
rect 4068 319404 4120 319456
rect 15844 319404 15896 319456
rect 98000 319404 98052 319456
rect 141424 319404 141476 319456
rect 182088 319404 182140 319456
rect 215300 319404 215352 319456
rect 233976 319404 234028 319456
rect 276204 319404 276256 319456
rect 259368 319336 259420 319388
rect 263784 319336 263836 319388
rect 175924 318792 175976 318844
rect 246488 318792 246540 318844
rect 71964 318044 72016 318096
rect 88984 318044 89036 318096
rect 103428 318044 103480 318096
rect 114560 318044 114612 318096
rect 144828 317500 144880 317552
rect 197452 317500 197504 317552
rect 142804 317432 142856 317484
rect 261024 317432 261076 317484
rect 184204 317364 184256 317416
rect 184664 317364 184716 317416
rect 214012 316752 214064 316804
rect 214564 316752 214616 316804
rect 119344 316684 119396 316736
rect 190460 316684 190512 316736
rect 215300 316684 215352 316736
rect 254676 316684 254728 316736
rect 579620 316684 579672 316736
rect 87604 316616 87656 316668
rect 88248 316616 88300 316668
rect 192484 316072 192536 316124
rect 214564 316072 214616 316124
rect 88248 316004 88300 316056
rect 110512 316004 110564 316056
rect 184664 316004 184716 316056
rect 257344 316004 257396 316056
rect 228364 315256 228416 315308
rect 265072 315256 265124 315308
rect 190460 315188 190512 315240
rect 191564 315188 191616 315240
rect 195244 315188 195296 315240
rect 178684 314644 178736 314696
rect 179328 314644 179380 314696
rect 226340 314644 226392 314696
rect 216036 313896 216088 313948
rect 236552 313896 236604 313948
rect 239404 313896 239456 313948
rect 269396 313896 269448 313948
rect 167644 313352 167696 313404
rect 208400 313352 208452 313404
rect 164884 313284 164936 313336
rect 211344 313284 211396 313336
rect 238668 313284 238720 313336
rect 279056 313284 279108 313336
rect 246488 312536 246540 312588
rect 273260 312536 273312 312588
rect 185584 311924 185636 311976
rect 186136 311924 186188 311976
rect 262496 311924 262548 311976
rect 151268 311856 151320 311908
rect 231860 311856 231912 311908
rect 218060 311108 218112 311160
rect 249616 311108 249668 311160
rect 181444 310564 181496 310616
rect 267740 310564 267792 310616
rect 115848 310496 115900 310548
rect 217416 310496 217468 310548
rect 57612 310428 57664 310480
rect 57888 310428 57940 310480
rect 112536 310428 112588 310480
rect 114652 310428 114704 310480
rect 168380 310428 168432 310480
rect 169024 310428 169076 310480
rect 57520 309884 57572 309936
rect 80060 309884 80112 309936
rect 57888 309748 57940 309800
rect 168380 309748 168432 309800
rect 187056 309204 187108 309256
rect 259552 309204 259604 309256
rect 170404 309136 170456 309188
rect 271880 309136 271932 309188
rect 184572 309068 184624 309120
rect 187700 309068 187752 309120
rect 84200 308388 84252 308440
rect 151176 308388 151228 308440
rect 223580 308388 223632 308440
rect 255964 308388 256016 308440
rect 4068 307776 4120 307828
rect 7564 307776 7616 307828
rect 148324 307776 148376 307828
rect 216036 307776 216088 307828
rect 251824 307776 251876 307828
rect 282920 307776 282972 307828
rect 233240 307096 233292 307148
rect 252560 307096 252612 307148
rect 199384 307028 199436 307080
rect 203984 307028 204036 307080
rect 226340 307028 226392 307080
rect 262312 307028 262364 307080
rect 253204 306552 253256 306604
rect 258264 306552 258316 306604
rect 152464 306416 152516 306468
rect 214196 306416 214248 306468
rect 9588 306348 9640 306400
rect 197360 306348 197412 306400
rect 213276 305736 213328 305788
rect 231584 305736 231636 305788
rect 222844 305600 222896 305652
rect 246028 305600 246080 305652
rect 191380 305056 191432 305108
rect 193312 305056 193364 305108
rect 193496 305056 193548 305108
rect 202788 305056 202840 305108
rect 249248 305056 249300 305108
rect 249708 305056 249760 305108
rect 278780 305056 278832 305108
rect 137284 304988 137336 305040
rect 216588 304988 216640 305040
rect 240048 304988 240100 305040
rect 270684 304988 270736 305040
rect 218704 304920 218756 304972
rect 220820 304920 220872 304972
rect 97908 304308 97960 304360
rect 108396 304308 108448 304360
rect 123484 304308 123536 304360
rect 151084 304308 151136 304360
rect 151360 304308 151412 304360
rect 164884 304308 164936 304360
rect 226984 304308 227036 304360
rect 236368 304308 236420 304360
rect 60464 304240 60516 304292
rect 170496 304240 170548 304292
rect 213184 304240 213236 304292
rect 223212 304240 223264 304292
rect 231124 304240 231176 304292
rect 253204 304240 253256 304292
rect 226524 303764 226576 303816
rect 231032 303764 231084 303816
rect 186044 303696 186096 303748
rect 196256 303696 196308 303748
rect 221464 303696 221516 303748
rect 224408 303696 224460 303748
rect 193220 303628 193272 303680
rect 193588 303628 193640 303680
rect 211344 303628 211396 303680
rect 212172 303628 212224 303680
rect 215944 303628 215996 303680
rect 217232 303628 217284 303680
rect 220912 303628 220964 303680
rect 221740 303628 221792 303680
rect 222936 303628 222988 303680
rect 226248 303628 226300 303680
rect 243084 303628 243136 303680
rect 243820 303628 243872 303680
rect 248420 303628 248472 303680
rect 248972 303628 249024 303680
rect 265164 303628 265216 303680
rect 176660 302880 176712 302932
rect 177396 302880 177448 302932
rect 192668 302880 192720 302932
rect 197360 302880 197412 302932
rect 211252 302880 211304 302932
rect 233148 302880 233200 302932
rect 254124 302880 254176 302932
rect 257436 302880 257488 302932
rect 261116 302880 261168 302932
rect 87696 302268 87748 302320
rect 176660 302268 176712 302320
rect 192576 302268 192628 302320
rect 218428 302268 218480 302320
rect 15844 302200 15896 302252
rect 198004 302200 198056 302252
rect 247684 302200 247736 302252
rect 281540 302200 281592 302252
rect 252468 302132 252520 302184
rect 258448 302132 258500 302184
rect 240876 301656 240928 301708
rect 73068 301452 73120 301504
rect 173624 301452 173676 301504
rect 176108 301452 176160 301504
rect 252928 301452 252980 301504
rect 193312 301044 193364 301096
rect 195244 301044 195296 301096
rect 188528 300976 188580 301028
rect 206928 300976 206980 301028
rect 178868 300908 178920 300960
rect 192484 300908 192536 300960
rect 199476 300908 199528 300960
rect 214564 300908 214616 300960
rect 191472 300772 191524 300824
rect 245108 301044 245160 301096
rect 242072 300976 242124 301028
rect 258724 300908 258776 300960
rect 259460 300908 259512 300960
rect 255412 300840 255464 300892
rect 278044 300840 278096 300892
rect 252468 300772 252520 300824
rect 124956 300092 125008 300144
rect 159456 300092 159508 300144
rect 164240 300092 164292 300144
rect 255780 299548 255832 299600
rect 259368 299548 259420 299600
rect 164240 299480 164292 299532
rect 191748 299480 191800 299532
rect 255412 299480 255464 299532
rect 288716 299480 288768 299532
rect 281356 299412 281408 299464
rect 580172 299412 580224 299464
rect 92848 298732 92900 298784
rect 130476 298732 130528 298784
rect 170496 298732 170548 298784
rect 187516 298732 187568 298784
rect 191012 298800 191064 298852
rect 275284 298800 275336 298852
rect 280252 298800 280304 298852
rect 281356 298800 281408 298852
rect 259368 298732 259420 298784
rect 293960 298732 294012 298784
rect 257344 298188 257396 298240
rect 258172 298188 258224 298240
rect 255412 298120 255464 298172
rect 266636 298120 266688 298172
rect 164148 298052 164200 298104
rect 191748 298052 191800 298104
rect 255412 297712 255464 297764
rect 259460 297712 259512 297764
rect 91192 297372 91244 297424
rect 104348 297372 104400 297424
rect 117228 297372 117280 297424
rect 164148 297372 164200 297424
rect 253296 296692 253348 296744
rect 296720 296692 296772 296744
rect 255504 296080 255556 296132
rect 255688 296080 255740 296132
rect 130568 296012 130620 296064
rect 191564 296012 191616 296064
rect 78588 295944 78640 295996
rect 255504 295944 255556 295996
rect 265256 295944 265308 295996
rect 284484 295944 284536 295996
rect 189080 295876 189132 295928
rect 189724 295876 189776 295928
rect 77392 295332 77444 295384
rect 78588 295332 78640 295384
rect 191288 295332 191340 295384
rect 193404 295332 193456 295384
rect 86960 294652 87012 294704
rect 152648 294652 152700 294704
rect 19248 294584 19300 294636
rect 149704 294584 149756 294636
rect 152740 294584 152792 294636
rect 189908 294584 189960 294636
rect 255412 294584 255464 294636
rect 258264 294584 258316 294636
rect 280344 294584 280396 294636
rect 255412 293972 255464 294024
rect 277584 293972 277636 294024
rect 93768 293904 93820 293956
rect 117228 293904 117280 293956
rect 138020 293904 138072 293956
rect 143632 293904 143684 293956
rect 155776 293904 155828 293956
rect 191196 293904 191248 293956
rect 253848 293904 253900 293956
rect 269120 293904 269172 293956
rect 58992 293224 59044 293276
rect 78680 293224 78732 293276
rect 96712 293224 96764 293276
rect 141700 293224 141752 293276
rect 166908 293224 166960 293276
rect 187700 293224 187752 293276
rect 255504 293224 255556 293276
rect 258448 293224 258500 293276
rect 290004 293224 290056 293276
rect 3516 292544 3568 292596
rect 14464 292544 14516 292596
rect 65800 291796 65852 291848
rect 86224 291796 86276 291848
rect 163688 291796 163740 291848
rect 178960 291796 179012 291848
rect 256424 291796 256476 291848
rect 264980 291796 265032 291848
rect 253848 291728 253900 291780
rect 256608 291728 256660 291780
rect 85856 291184 85908 291236
rect 86776 291184 86828 291236
rect 104900 291252 104952 291304
rect 95148 291184 95200 291236
rect 127716 291184 127768 291236
rect 256516 291048 256568 291100
rect 263876 291048 263928 291100
rect 98460 290504 98512 290556
rect 138020 290504 138072 290556
rect 173164 290504 173216 290556
rect 184204 290504 184256 290556
rect 33784 290436 33836 290488
rect 87604 290436 87656 290488
rect 106188 290436 106240 290488
rect 177488 290436 177540 290488
rect 71872 289824 71924 289876
rect 104992 289824 105044 289876
rect 106188 289824 106240 289876
rect 177580 289824 177632 289876
rect 191748 289824 191800 289876
rect 79968 289756 80020 289808
rect 173808 289756 173860 289808
rect 191656 289756 191708 289808
rect 61844 289076 61896 289128
rect 77484 289076 77536 289128
rect 80152 289076 80204 289128
rect 180708 289076 180760 289128
rect 184204 289076 184256 289128
rect 255964 288872 256016 288924
rect 259736 288872 259788 288924
rect 97540 288396 97592 288448
rect 97908 288396 97960 288448
rect 109040 288396 109092 288448
rect 259368 288396 259420 288448
rect 261116 288396 261168 288448
rect 255872 288328 255924 288380
rect 276112 288328 276164 288380
rect 255780 288260 255832 288312
rect 258080 288260 258132 288312
rect 116492 287716 116544 287768
rect 184848 287716 184900 287768
rect 191748 287716 191800 287768
rect 78588 287648 78640 287700
rect 186964 287648 187016 287700
rect 87880 287036 87932 287088
rect 88156 287036 88208 287088
rect 104348 287036 104400 287088
rect 276756 287036 276808 287088
rect 279056 287036 279108 287088
rect 61936 286968 61988 287020
rect 65984 286968 66036 287020
rect 95792 286968 95844 287020
rect 97540 286968 97592 287020
rect 127716 286968 127768 287020
rect 142896 286968 142948 287020
rect 256608 286628 256660 286680
rect 261024 286628 261076 286680
rect 75736 286288 75788 286340
rect 185584 286288 185636 286340
rect 90916 286220 90968 286272
rect 94504 286220 94556 286272
rect 85304 285880 85356 285932
rect 87696 285880 87748 285932
rect 68652 285744 68704 285796
rect 81256 285812 81308 285864
rect 83464 285812 83516 285864
rect 71320 285676 71372 285728
rect 72424 285676 72476 285728
rect 74816 285676 74868 285728
rect 75828 285676 75880 285728
rect 79232 285676 79284 285728
rect 79968 285676 80020 285728
rect 256424 285676 256476 285728
rect 262496 285676 262548 285728
rect 263968 285676 264020 285728
rect 256608 285608 256660 285660
rect 263600 285608 263652 285660
rect 140044 284996 140096 285048
rect 149796 284996 149848 285048
rect 75920 284928 75972 284980
rect 76380 284928 76432 284980
rect 149704 284928 149756 284980
rect 180156 284928 180208 284980
rect 266636 284792 266688 284844
rect 267832 284792 267884 284844
rect 53564 284452 53616 284504
rect 71320 284452 71372 284504
rect 70860 284384 70912 284436
rect 99380 284384 99432 284436
rect 67364 284316 67416 284368
rect 160100 284316 160152 284368
rect 167828 284316 167880 284368
rect 191748 284316 191800 284368
rect 149060 284248 149112 284300
rect 256608 284248 256660 284300
rect 294052 284248 294104 284300
rect 191748 284180 191800 284232
rect 256332 284180 256384 284232
rect 273260 284180 273312 284232
rect 88294 283704 88346 283756
rect 89536 283704 89588 283756
rect 92710 283704 92762 283756
rect 93768 283704 93820 283756
rect 96896 283364 96948 283416
rect 97264 283364 97316 283416
rect 184664 283228 184716 283280
rect 187700 283228 187752 283280
rect 86868 283024 86920 283076
rect 98920 283024 98972 283076
rect 63224 282956 63276 283008
rect 76012 282956 76064 283008
rect 94136 282956 94188 283008
rect 98828 282956 98880 283008
rect 56416 282888 56468 282940
rect 66260 282888 66312 282940
rect 68836 282888 68888 282940
rect 173808 282888 173860 282940
rect 175924 282888 175976 282940
rect 119344 282820 119396 282872
rect 124956 282820 125008 282872
rect 44088 282140 44140 282192
rect 63500 282140 63552 282192
rect 135904 282140 135956 282192
rect 191840 282140 191892 282192
rect 255504 282140 255556 282192
rect 259828 282140 259880 282192
rect 263692 282140 263744 282192
rect 63500 281596 63552 281648
rect 64604 281596 64656 281648
rect 102784 281596 102836 281648
rect 100760 281528 100812 281580
rect 180340 281528 180392 281580
rect 181536 281528 181588 281580
rect 190460 281528 190512 281580
rect 255320 281460 255372 281512
rect 281816 281460 281868 281512
rect 255504 281392 255556 281444
rect 262312 281392 262364 281444
rect 119344 280848 119396 280900
rect 155316 280848 155368 280900
rect 176476 280848 176528 280900
rect 190552 280848 190604 280900
rect 99380 280780 99432 280832
rect 162676 280780 162728 280832
rect 178684 280780 178736 280832
rect 4804 280168 4856 280220
rect 67548 280168 67600 280220
rect 68836 280168 68888 280220
rect 100852 280100 100904 280152
rect 162124 280100 162176 280152
rect 165528 280100 165580 280152
rect 175280 280100 175332 280152
rect 255504 280100 255556 280152
rect 291384 280100 291436 280152
rect 159456 280032 159508 280084
rect 160100 280032 160152 280084
rect 190460 280032 190512 280084
rect 3424 279624 3476 279676
rect 7656 279624 7708 279676
rect 7564 279420 7616 279472
rect 37096 279420 37148 279472
rect 60464 279420 60516 279472
rect 66812 279420 66864 279472
rect 179328 279420 179380 279472
rect 191288 279420 191340 279472
rect 262312 279420 262364 279472
rect 270592 279420 270644 279472
rect 255320 278740 255372 278792
rect 262312 278740 262364 278792
rect 64604 278672 64656 278724
rect 66812 278672 66864 278724
rect 100760 278604 100812 278656
rect 104440 278604 104492 278656
rect 112812 278060 112864 278112
rect 116584 278060 116636 278112
rect 144184 278060 144236 278112
rect 167644 278060 167696 278112
rect 255504 278060 255556 278112
rect 266544 278060 266596 278112
rect 112628 277992 112680 278044
rect 152556 277992 152608 278044
rect 190276 277992 190328 278044
rect 190460 277992 190512 278044
rect 258080 277992 258132 278044
rect 295524 277992 295576 278044
rect 52368 277312 52420 277364
rect 66812 277312 66864 277364
rect 100760 277312 100812 277364
rect 123484 277312 123536 277364
rect 255320 277312 255372 277364
rect 271972 277312 272024 277364
rect 255504 277244 255556 277296
rect 267740 277244 267792 277296
rect 98920 276632 98972 276684
rect 176660 276632 176712 276684
rect 63316 276020 63368 276072
rect 67640 276020 67692 276072
rect 148508 276020 148560 276072
rect 190460 276020 190512 276072
rect 57888 275952 57940 276004
rect 66812 275952 66864 276004
rect 176660 275952 176712 276004
rect 177856 275952 177908 276004
rect 181444 275952 181496 276004
rect 255320 275952 255372 276004
rect 270500 275952 270552 276004
rect 255504 275476 255556 275528
rect 258080 275476 258132 275528
rect 101680 275340 101732 275392
rect 136088 275340 136140 275392
rect 57704 275272 57756 275324
rect 66444 275272 66496 275324
rect 66720 275272 66772 275324
rect 100944 275272 100996 275324
rect 169208 275272 169260 275324
rect 259368 275272 259420 275324
rect 292580 275272 292632 275324
rect 184848 274728 184900 274780
rect 186412 274728 186464 274780
rect 187056 274728 187108 274780
rect 190552 274728 190604 274780
rect 171968 274660 172020 274712
rect 190460 274660 190512 274712
rect 100760 274592 100812 274644
rect 170404 274592 170456 274644
rect 255320 274592 255372 274644
rect 281724 274592 281776 274644
rect 100852 274524 100904 274576
rect 135996 274524 136048 274576
rect 255504 274252 255556 274304
rect 259276 274252 259328 274304
rect 259552 274252 259604 274304
rect 145748 273912 145800 273964
rect 159548 273912 159600 273964
rect 58900 273300 58952 273352
rect 60648 273300 60700 273352
rect 66812 273300 66864 273352
rect 182916 273232 182968 273284
rect 190460 273232 190512 273284
rect 100760 273164 100812 273216
rect 129740 273164 129792 273216
rect 278688 272960 278740 273012
rect 281724 272960 281776 273012
rect 255504 272892 255556 272944
rect 259368 272892 259420 272944
rect 146944 272552 146996 272604
rect 173164 272552 173216 272604
rect 100024 272484 100076 272536
rect 115940 272484 115992 272536
rect 129740 272484 129792 272536
rect 159548 272484 159600 272536
rect 61660 271940 61712 271992
rect 61936 271940 61988 271992
rect 66812 271940 66864 271992
rect 181444 271872 181496 271924
rect 190828 271872 190880 271924
rect 101128 271804 101180 271856
rect 101864 271804 101916 271856
rect 128728 271804 128780 271856
rect 271972 271804 272024 271856
rect 276020 271804 276072 271856
rect 128728 271192 128780 271244
rect 129648 271192 129700 271244
rect 135996 271192 136048 271244
rect 137376 271192 137428 271244
rect 188528 271192 188580 271244
rect 98828 271124 98880 271176
rect 155316 271124 155368 271176
rect 255504 270920 255556 270972
rect 258724 270920 258776 270972
rect 63408 270580 63460 270632
rect 64604 270580 64656 270632
rect 66812 270580 66864 270632
rect 188436 270580 188488 270632
rect 191656 270580 191708 270632
rect 255504 270512 255556 270564
rect 271972 270512 272024 270564
rect 57244 270444 57296 270496
rect 57796 270444 57848 270496
rect 66628 270444 66680 270496
rect 100760 270444 100812 270496
rect 112536 270444 112588 270496
rect 255320 270444 255372 270496
rect 277492 270444 277544 270496
rect 255504 270376 255556 270428
rect 262404 270376 262456 270428
rect 262680 270376 262732 270428
rect 152648 269832 152700 269884
rect 171784 269832 171836 269884
rect 98736 269764 98788 269816
rect 160928 269764 160980 269816
rect 187148 269152 187200 269204
rect 191564 269152 191616 269204
rect 53288 269084 53340 269136
rect 57244 269084 57296 269136
rect 170588 269084 170640 269136
rect 190828 269084 190880 269136
rect 262680 269084 262732 269136
rect 269304 269084 269356 269136
rect 267832 269016 267884 269068
rect 270776 269016 270828 269068
rect 166816 268608 166868 268660
rect 168380 268608 168432 268660
rect 100116 268404 100168 268456
rect 134708 268404 134760 268456
rect 145564 268404 145616 268456
rect 173256 268404 173308 268456
rect 113824 268336 113876 268388
rect 166356 268336 166408 268388
rect 100760 267996 100812 268048
rect 104256 267996 104308 268048
rect 255504 267792 255556 267844
rect 267832 267792 267884 267844
rect 54944 267724 54996 267776
rect 57796 267724 57848 267776
rect 66812 267724 66864 267776
rect 173164 267724 173216 267776
rect 191656 267724 191708 267776
rect 3516 267656 3568 267708
rect 33784 267656 33836 267708
rect 291292 267656 291344 267708
rect 580264 267656 580316 267708
rect 174544 267112 174596 267164
rect 180800 267112 180852 267164
rect 102232 266976 102284 267028
rect 115204 266976 115256 267028
rect 175188 266976 175240 267028
rect 189080 266976 189132 267028
rect 257344 266976 257396 267028
rect 291292 266976 291344 267028
rect 62028 266364 62080 266416
rect 64788 266364 64840 266416
rect 66812 266364 66864 266416
rect 100760 266364 100812 266416
rect 147128 266364 147180 266416
rect 255320 266364 255372 266416
rect 262404 266364 262456 266416
rect 255504 266296 255556 266348
rect 265072 266296 265124 266348
rect 117320 266024 117372 266076
rect 123484 266024 123536 266076
rect 130476 265616 130528 265668
rect 147036 265616 147088 265668
rect 266728 265616 266780 265668
rect 280160 265616 280212 265668
rect 52276 265004 52328 265056
rect 54852 265004 54904 265056
rect 163504 265004 163556 265056
rect 190828 265004 190880 265056
rect 64788 264936 64840 264988
rect 66536 264936 66588 264988
rect 100760 264936 100812 264988
rect 138848 264936 138900 264988
rect 157984 264936 158036 264988
rect 191656 264936 191708 264988
rect 255504 264936 255556 264988
rect 266452 264936 266504 264988
rect 266728 264936 266780 264988
rect 147680 264868 147732 264920
rect 148968 264868 149020 264920
rect 181536 264868 181588 264920
rect 131764 264256 131816 264308
rect 151360 264256 151412 264308
rect 53656 264188 53708 264240
rect 66260 264188 66312 264240
rect 100944 264188 100996 264240
rect 147680 264188 147732 264240
rect 276940 264188 276992 264240
rect 284576 264188 284628 264240
rect 59176 263644 59228 263696
rect 66812 263644 66864 263696
rect 255320 263644 255372 263696
rect 260840 263644 260892 263696
rect 100852 263576 100904 263628
rect 104440 263576 104492 263628
rect 164884 263576 164936 263628
rect 191656 263576 191708 263628
rect 255504 263576 255556 263628
rect 276020 263576 276072 263628
rect 276940 263576 276992 263628
rect 100760 263508 100812 263560
rect 145656 263508 145708 263560
rect 273352 262828 273404 262880
rect 281264 262828 281316 262880
rect 256424 262284 256476 262336
rect 265348 262284 265400 262336
rect 265808 262284 265860 262336
rect 7748 262216 7800 262268
rect 65892 262216 65944 262268
rect 66536 262216 66588 262268
rect 167644 262216 167696 262268
rect 191656 262216 191708 262268
rect 280804 262148 280856 262200
rect 281264 262148 281316 262200
rect 287336 262148 287388 262200
rect 52368 261536 52420 261588
rect 61016 261536 61068 261588
rect 61752 261536 61804 261588
rect 104348 261536 104400 261588
rect 117964 261536 118016 261588
rect 124956 261536 125008 261588
rect 169576 261536 169628 261588
rect 7564 261468 7616 261520
rect 67088 261468 67140 261520
rect 103428 261468 103480 261520
rect 106280 261468 106332 261520
rect 113088 261468 113140 261520
rect 166264 261468 166316 261520
rect 258724 261536 258776 261588
rect 279056 261536 279108 261588
rect 182824 261468 182876 261520
rect 256608 261468 256660 261520
rect 280252 261468 280304 261520
rect 281448 261468 281500 261520
rect 178684 260856 178736 260908
rect 191656 260856 191708 260908
rect 281448 260856 281500 260908
rect 295340 260856 295392 260908
rect 50896 260176 50948 260228
rect 65800 260176 65852 260228
rect 66536 260176 66588 260228
rect 39948 260108 40000 260160
rect 60464 260108 60516 260160
rect 256608 260108 256660 260160
rect 263232 260108 263284 260160
rect 285680 260108 285732 260160
rect 288532 260108 288584 260160
rect 100760 259496 100812 259548
rect 155408 259496 155460 259548
rect 177304 259496 177356 259548
rect 191656 259496 191708 259548
rect 100852 259428 100904 259480
rect 185676 259428 185728 259480
rect 258724 259428 258776 259480
rect 285680 259428 285732 259480
rect 101404 259360 101456 259412
rect 154488 259360 154540 259412
rect 104808 258816 104860 258868
rect 111064 258816 111116 258868
rect 46848 258748 46900 258800
rect 64512 258748 64564 258800
rect 66352 258748 66404 258800
rect 255964 258748 256016 258800
rect 265072 258748 265124 258800
rect 41144 258680 41196 258732
rect 66260 258680 66312 258732
rect 156696 258680 156748 258732
rect 171876 258680 171928 258732
rect 256608 258680 256660 258732
rect 271880 258680 271932 258732
rect 274732 258680 274784 258732
rect 287152 258680 287204 258732
rect 265072 258612 265124 258664
rect 265348 258612 265400 258664
rect 174544 258068 174596 258120
rect 190460 258068 190512 258120
rect 50804 258000 50856 258052
rect 66444 258000 66496 258052
rect 100760 258000 100812 258052
rect 104164 258000 104216 258052
rect 256332 258000 256384 258052
rect 258724 258000 258776 258052
rect 267740 258000 267792 258052
rect 288624 258000 288676 258052
rect 66352 257932 66404 257984
rect 68192 257932 68244 257984
rect 102048 257388 102100 257440
rect 130568 257388 130620 257440
rect 256608 257388 256660 257440
rect 267740 257388 267792 257440
rect 44088 257320 44140 257372
rect 50804 257320 50856 257372
rect 113916 257320 113968 257372
rect 184296 257320 184348 257372
rect 258172 257320 258224 257372
rect 286232 257320 286284 257372
rect 175924 256708 175976 256760
rect 191656 256708 191708 256760
rect 286232 256708 286284 256760
rect 287152 256708 287204 256760
rect 286324 256640 286376 256692
rect 580908 256640 580960 256692
rect 184204 256164 184256 256216
rect 192668 256164 192720 256216
rect 41236 255960 41288 256012
rect 53472 255960 53524 256012
rect 60004 255960 60056 256012
rect 100852 255960 100904 256012
rect 178868 255960 178920 256012
rect 256608 255960 256660 256012
rect 276388 255960 276440 256012
rect 278964 255960 279016 256012
rect 278044 255824 278096 255876
rect 285680 255824 285732 255876
rect 63132 255416 63184 255468
rect 66260 255416 66312 255468
rect 100760 255280 100812 255332
rect 164976 255280 165028 255332
rect 180156 255280 180208 255332
rect 190644 255280 190696 255332
rect 256608 255280 256660 255332
rect 262496 255280 262548 255332
rect 48136 255212 48188 255264
rect 66812 255212 66864 255264
rect 137468 255212 137520 255264
rect 177580 255212 177632 255264
rect 2780 255144 2832 255196
rect 4804 255144 4856 255196
rect 100760 254872 100812 254924
rect 104256 254872 104308 254924
rect 256608 254600 256660 254652
rect 274732 254600 274784 254652
rect 60004 254532 60056 254584
rect 66812 254532 66864 254584
rect 115296 254532 115348 254584
rect 137468 254532 137520 254584
rect 171048 254532 171100 254584
rect 176016 254532 176068 254584
rect 259368 254532 259420 254584
rect 289912 254532 289964 254584
rect 185584 253988 185636 254040
rect 191656 253988 191708 254040
rect 46848 253920 46900 253972
rect 48136 253920 48188 253972
rect 100760 253920 100812 253972
rect 115204 253920 115256 253972
rect 182824 253920 182876 253972
rect 191564 253920 191616 253972
rect 111064 253240 111116 253292
rect 122196 253240 122248 253292
rect 7656 253172 7708 253224
rect 66996 253172 67048 253224
rect 67364 253172 67416 253224
rect 108396 253172 108448 253224
rect 123576 253172 123628 253224
rect 138664 253172 138716 253224
rect 162308 253172 162360 253224
rect 254124 253036 254176 253088
rect 259368 253036 259420 253088
rect 158168 252764 158220 252816
rect 161020 252764 161072 252816
rect 100760 252560 100812 252612
rect 111156 252560 111208 252612
rect 170404 252560 170456 252612
rect 191656 252560 191708 252612
rect 255780 252560 255832 252612
rect 258356 252560 258408 252612
rect 273352 252560 273404 252612
rect 275284 252560 275336 252612
rect 100852 252492 100904 252544
rect 119344 252492 119396 252544
rect 116768 251880 116820 251932
rect 158168 251880 158220 251932
rect 55036 251812 55088 251864
rect 66076 251812 66128 251864
rect 66628 251812 66680 251864
rect 129188 251812 129240 251864
rect 180248 251812 180300 251864
rect 189816 251812 189868 251864
rect 190368 251812 190420 251864
rect 193220 251812 193272 251864
rect 270408 251812 270460 251864
rect 582472 251812 582524 251864
rect 100760 251336 100812 251388
rect 103520 251336 103572 251388
rect 256424 251268 256476 251320
rect 269396 251268 269448 251320
rect 270408 251268 270460 251320
rect 166264 251200 166316 251252
rect 191656 251200 191708 251252
rect 256608 251200 256660 251252
rect 271880 251200 271932 251252
rect 60556 250724 60608 250776
rect 66812 250724 66864 250776
rect 100760 250520 100812 250572
rect 106924 250520 106976 250572
rect 102784 250452 102836 250504
rect 153844 250452 153896 250504
rect 256608 250452 256660 250504
rect 273352 250452 273404 250504
rect 256700 250316 256752 250368
rect 257344 250316 257396 250368
rect 169024 249772 169076 249824
rect 190644 249772 190696 249824
rect 100944 249704 100996 249756
rect 108488 249704 108540 249756
rect 108948 249704 109000 249756
rect 162124 249704 162176 249756
rect 163688 249704 163740 249756
rect 108488 249092 108540 249144
rect 129096 249092 129148 249144
rect 148508 249092 148560 249144
rect 120816 249024 120868 249076
rect 160836 249024 160888 249076
rect 256608 248480 256660 248532
rect 278044 248480 278096 248532
rect 53380 248412 53432 248464
rect 57888 248412 57940 248464
rect 66812 248412 66864 248464
rect 188344 248412 188396 248464
rect 190828 248412 190880 248464
rect 256240 248412 256292 248464
rect 291292 248412 291344 248464
rect 582380 248412 582432 248464
rect 254676 248344 254728 248396
rect 286324 248344 286376 248396
rect 135168 247664 135220 247716
rect 167828 247664 167880 247716
rect 60556 247052 60608 247104
rect 66536 247052 66588 247104
rect 100944 246984 100996 247036
rect 104808 247052 104860 247104
rect 133880 247052 133932 247104
rect 135168 247052 135220 247104
rect 256608 246984 256660 247036
rect 283012 246984 283064 247036
rect 288532 246984 288584 247036
rect 102324 246304 102376 246356
rect 155960 246304 156012 246356
rect 162768 246304 162820 246356
rect 168288 246304 168340 246356
rect 175280 246304 175332 246356
rect 186228 246304 186280 246356
rect 193588 246304 193640 246356
rect 253940 246032 253992 246084
rect 258172 246032 258224 246084
rect 183468 245624 183520 245676
rect 191288 245624 191340 245676
rect 159548 245556 159600 245608
rect 190276 245556 190328 245608
rect 191840 245556 191892 245608
rect 100944 244944 100996 244996
rect 106280 244944 106332 244996
rect 107016 244944 107068 244996
rect 101036 244876 101088 244928
rect 165620 244876 165672 244928
rect 58900 244264 58952 244316
rect 66812 244264 66864 244316
rect 165620 244264 165672 244316
rect 166448 244264 166500 244316
rect 56508 244196 56560 244248
rect 66720 244196 66772 244248
rect 276388 244196 276440 244248
rect 278872 244196 278924 244248
rect 113916 243584 113968 243636
rect 140136 243584 140188 243636
rect 98000 243516 98052 243568
rect 98276 243516 98328 243568
rect 98276 243380 98328 243432
rect 192576 243516 192628 243568
rect 255320 243516 255372 243568
rect 287060 243516 287112 243568
rect 61752 242904 61804 242956
rect 66904 242904 66956 242956
rect 162768 242904 162820 242956
rect 192116 242904 192168 242956
rect 192484 242904 192536 242956
rect 67732 242496 67784 242548
rect 68790 242496 68842 242548
rect 112536 242224 112588 242276
rect 145748 242224 145800 242276
rect 134708 242156 134760 242208
rect 252836 242904 252888 242956
rect 255688 242904 255740 242956
rect 276388 242904 276440 242956
rect 276664 242904 276716 242956
rect 252376 242292 252428 242344
rect 252836 242292 252888 242344
rect 259644 242156 259696 242208
rect 195336 242020 195388 242072
rect 195796 242020 195848 242072
rect 248512 242020 248564 242072
rect 250444 242020 250496 242072
rect 155316 241884 155368 241936
rect 160744 241884 160796 241936
rect 68560 241748 68612 241800
rect 69388 241748 69440 241800
rect 94964 241612 95016 241664
rect 115296 241612 115348 241664
rect 59268 241544 59320 241596
rect 66812 241544 66864 241596
rect 58992 241476 59044 241528
rect 77438 241476 77490 241528
rect 93952 241476 94004 241528
rect 95976 241476 96028 241528
rect 99104 241476 99156 241528
rect 181996 241476 182048 241528
rect 201500 241476 201552 241528
rect 201960 241476 202012 241528
rect 255504 241476 255556 241528
rect 261116 241476 261168 241528
rect 73528 241408 73580 241460
rect 112628 241408 112680 241460
rect 192116 241408 192168 241460
rect 204352 241408 204404 241460
rect 268292 241408 268344 241460
rect 298100 241408 298152 241460
rect 67824 241340 67876 241392
rect 102324 241340 102376 241392
rect 3424 241068 3476 241120
rect 7748 241068 7800 241120
rect 136088 240796 136140 240848
rect 171140 240796 171192 240848
rect 164976 240728 165028 240780
rect 234620 240796 234672 240848
rect 256700 240796 256752 240848
rect 251824 240728 251876 240780
rect 276756 240728 276808 240780
rect 181536 240320 181588 240372
rect 186320 240320 186372 240372
rect 74540 240116 74592 240168
rect 75460 240116 75512 240168
rect 78680 240116 78732 240168
rect 79324 240116 79376 240168
rect 80060 240116 80112 240168
rect 80980 240116 81032 240168
rect 82820 240116 82872 240168
rect 83740 240116 83792 240168
rect 84200 240116 84252 240168
rect 84844 240116 84896 240168
rect 86960 240116 87012 240168
rect 87604 240116 87656 240168
rect 95240 240116 95292 240168
rect 95884 240116 95936 240168
rect 96620 240116 96672 240168
rect 97632 240116 97684 240168
rect 65984 240048 66036 240100
rect 70400 240048 70452 240100
rect 76104 240048 76156 240100
rect 77484 240048 77536 240100
rect 82176 240048 82228 240100
rect 86868 240048 86920 240100
rect 89628 240048 89680 240100
rect 182180 240048 182232 240100
rect 211804 240048 211856 240100
rect 233884 240048 233936 240100
rect 234620 240048 234672 240100
rect 242164 240048 242216 240100
rect 242716 240048 242768 240100
rect 272064 240048 272116 240100
rect 192668 239980 192720 240032
rect 196164 239980 196216 240032
rect 177948 239640 178000 239692
rect 178776 239640 178828 239692
rect 219440 239640 219492 239692
rect 221096 239640 221148 239692
rect 69480 239368 69532 239420
rect 89076 239368 89128 239420
rect 196164 239368 196216 239420
rect 206744 239368 206796 239420
rect 249064 239368 249116 239420
rect 267004 239368 267056 239420
rect 89352 238756 89404 238808
rect 219440 238756 219492 238808
rect 227076 238756 227128 238808
rect 230756 238756 230808 238808
rect 233148 238756 233200 238808
rect 237380 238756 237432 238808
rect 93768 238688 93820 238740
rect 107660 238688 107712 238740
rect 188988 238688 189040 238740
rect 80152 238620 80204 238672
rect 95976 238620 96028 238672
rect 177948 238620 178000 238672
rect 209136 238620 209188 238672
rect 74356 238484 74408 238536
rect 76656 238484 76708 238536
rect 170496 238076 170548 238128
rect 177948 238076 178000 238128
rect 45376 238008 45428 238060
rect 46756 238008 46808 238060
rect 74632 238008 74684 238060
rect 107568 238008 107620 238060
rect 170588 238008 170640 238060
rect 215300 238008 215352 238060
rect 261024 238008 261076 238060
rect 79416 237396 79468 237448
rect 80152 237396 80204 237448
rect 95056 237396 95108 237448
rect 98092 237396 98144 237448
rect 59084 237328 59136 237380
rect 76104 237328 76156 237380
rect 78772 237328 78824 237380
rect 108396 237328 108448 237380
rect 184756 237328 184808 237380
rect 233148 237328 233200 237380
rect 252284 237328 252336 237380
rect 287244 237328 287296 237380
rect 193772 237260 193824 237312
rect 215484 237260 215536 237312
rect 85580 237124 85632 237176
rect 88984 237124 89036 237176
rect 106924 237056 106976 237108
rect 113272 237056 113324 237108
rect 228364 236988 228416 237040
rect 230480 236988 230532 237040
rect 72976 236648 73028 236700
rect 79324 236648 79376 236700
rect 122196 236648 122248 236700
rect 124220 236648 124272 236700
rect 125508 236648 125560 236700
rect 171968 236648 172020 236700
rect 215484 236580 215536 236632
rect 216312 236580 216364 236632
rect 217968 236580 218020 236632
rect 220912 236580 220964 236632
rect 222108 236580 222160 236632
rect 107660 236444 107712 236496
rect 108396 236444 108448 236496
rect 76104 235968 76156 236020
rect 76748 235968 76800 236020
rect 97908 235968 97960 236020
rect 98184 235968 98236 236020
rect 249156 235968 249208 236020
rect 252376 235968 252428 236020
rect 191288 235900 191340 235952
rect 213920 235900 213972 235952
rect 249892 235832 249944 235884
rect 250536 235832 250588 235884
rect 288440 235900 288492 235952
rect 82912 235288 82964 235340
rect 112996 235288 113048 235340
rect 116676 235288 116728 235340
rect 64512 235220 64564 235272
rect 156788 235220 156840 235272
rect 164976 235220 165028 235272
rect 197176 235220 197228 235272
rect 243636 235220 243688 235272
rect 269212 235220 269264 235272
rect 213920 234608 213972 234660
rect 214656 234608 214708 234660
rect 283564 234608 283616 234660
rect 580264 234608 580316 234660
rect 166816 234540 166868 234592
rect 256792 234540 256844 234592
rect 166356 234132 166408 234184
rect 166816 234132 166868 234184
rect 94688 233928 94740 233980
rect 95332 233928 95384 233980
rect 61844 233860 61896 233912
rect 76564 233860 76616 233912
rect 77392 233860 77444 233912
rect 87696 233860 87748 233912
rect 91008 233860 91060 233912
rect 125416 233860 125468 233912
rect 128360 233860 128412 233912
rect 184296 233860 184348 233912
rect 215944 233860 215996 233912
rect 257988 233860 258040 233912
rect 265164 233860 265216 233912
rect 269764 233656 269816 233708
rect 274824 233656 274876 233708
rect 108304 233180 108356 233232
rect 108948 233180 109000 233232
rect 278044 233180 278096 233232
rect 278872 233180 278924 233232
rect 279056 233112 279108 233164
rect 73160 232500 73212 232552
rect 77300 232500 77352 232552
rect 78680 232500 78732 232552
rect 91008 232500 91060 232552
rect 102140 232500 102192 232552
rect 166448 232500 166500 232552
rect 196624 232500 196676 232552
rect 204904 232500 204956 232552
rect 252744 232500 252796 232552
rect 258724 232500 258776 232552
rect 270684 232500 270736 232552
rect 7656 231820 7708 231872
rect 96620 231820 96672 231872
rect 97264 231820 97316 231872
rect 278872 231820 278924 231872
rect 580172 231820 580224 231872
rect 89076 231752 89128 231804
rect 170496 231752 170548 231804
rect 215944 231752 215996 231804
rect 266452 231752 266504 231804
rect 67456 231684 67508 231736
rect 112536 231684 112588 231736
rect 63224 231072 63276 231124
rect 73436 231072 73488 231124
rect 138848 231072 138900 231124
rect 213828 231072 213880 231124
rect 224316 231072 224368 231124
rect 280804 231072 280856 231124
rect 80336 230392 80388 230444
rect 156604 230392 156656 230444
rect 164976 230392 165028 230444
rect 185676 230392 185728 230444
rect 262220 230392 262272 230444
rect 77576 229712 77628 229764
rect 105636 229712 105688 229764
rect 120724 229712 120776 229764
rect 160928 229712 160980 229764
rect 161020 229712 161072 229764
rect 204444 229712 204496 229764
rect 235908 229712 235960 229764
rect 255596 229712 255648 229764
rect 89720 229032 89772 229084
rect 105544 229032 105596 229084
rect 156788 229032 156840 229084
rect 273352 229032 273404 229084
rect 65892 228352 65944 228404
rect 76104 228352 76156 228404
rect 77208 228352 77260 228404
rect 156788 227808 156840 227860
rect 157248 227808 157300 227860
rect 77208 227740 77260 227792
rect 187700 227740 187752 227792
rect 188344 227740 188396 227792
rect 155408 227672 155460 227724
rect 277400 227672 277452 227724
rect 105544 227060 105596 227112
rect 118700 227060 118752 227112
rect 84016 226992 84068 227044
rect 84200 226992 84252 227044
rect 87052 226992 87104 227044
rect 104164 226992 104216 227044
rect 110512 226992 110564 227044
rect 195336 226992 195388 227044
rect 224224 226992 224276 227044
rect 254584 226992 254636 227044
rect 95148 226312 95200 226364
rect 100852 226312 100904 226364
rect 80060 226244 80112 226296
rect 113180 226244 113232 226296
rect 113916 226244 113968 226296
rect 245568 225632 245620 225684
rect 257344 225632 257396 225684
rect 242808 225564 242860 225616
rect 290004 225564 290056 225616
rect 100024 224952 100076 225004
rect 242256 224952 242308 225004
rect 242808 224952 242860 225004
rect 176016 224884 176068 224936
rect 259736 224884 259788 224936
rect 76748 224204 76800 224256
rect 108304 224204 108356 224256
rect 121368 224204 121420 224256
rect 187056 224204 187108 224256
rect 196624 223524 196676 223576
rect 234620 223524 234672 223576
rect 235540 223524 235592 223576
rect 237472 223524 237524 223576
rect 237932 223524 237984 223576
rect 204444 223456 204496 223508
rect 80704 222844 80756 222896
rect 104992 222844 105044 222896
rect 111708 222844 111760 222896
rect 188436 222844 188488 222896
rect 255320 222844 255372 222896
rect 287336 222844 287388 222896
rect 580356 222844 580408 222896
rect 153844 222096 153896 222148
rect 252836 222096 252888 222148
rect 133236 221484 133288 221536
rect 148416 221484 148468 221536
rect 82820 221416 82872 221468
rect 204996 221416 205048 221468
rect 227812 221416 227864 221468
rect 255320 221416 255372 221468
rect 88340 220736 88392 220788
rect 121460 220736 121512 220788
rect 122196 220736 122248 220788
rect 163688 220736 163740 220788
rect 164148 220736 164200 220788
rect 227076 220736 227128 220788
rect 118608 220056 118660 220108
rect 182916 220056 182968 220108
rect 226984 220056 227036 220108
rect 251916 220056 251968 220108
rect 232596 218764 232648 218816
rect 283564 218764 283616 218816
rect 147128 218696 147180 218748
rect 236000 218696 236052 218748
rect 101496 217948 101548 218000
rect 103520 217948 103572 218000
rect 284484 217948 284536 218000
rect 104348 217880 104400 217932
rect 245568 217880 245620 217932
rect 256608 217268 256660 217320
rect 273444 217268 273496 217320
rect 245568 216656 245620 216708
rect 246304 216656 246356 216708
rect 160928 216588 160980 216640
rect 161388 216588 161440 216640
rect 278872 216588 278924 216640
rect 49608 215908 49660 215960
rect 162124 215908 162176 215960
rect 3424 214956 3476 215008
rect 7564 214956 7616 215008
rect 8208 214956 8260 215008
rect 86960 214548 87012 214600
rect 111800 214548 111852 214600
rect 218704 214548 218756 214600
rect 237656 214548 237708 214600
rect 111800 213936 111852 213988
rect 196624 213936 196676 213988
rect 100116 213188 100168 213240
rect 266360 213188 266412 213240
rect 181536 212440 181588 212492
rect 182088 212440 182140 212492
rect 249156 212440 249208 212492
rect 236644 212236 236696 212288
rect 237472 212236 237524 212288
rect 58900 211760 58952 211812
rect 159548 211760 159600 211812
rect 259368 211760 259420 211812
rect 582656 211760 582708 211812
rect 253848 211148 253900 211200
rect 258172 211148 258224 211200
rect 259368 211148 259420 211200
rect 56508 211080 56560 211132
rect 167736 211080 167788 211132
rect 287060 211080 287112 211132
rect 161296 209720 161348 209772
rect 232596 209720 232648 209772
rect 160836 209516 160888 209568
rect 161296 209516 161348 209568
rect 97264 209040 97316 209092
rect 129740 209040 129792 209092
rect 129740 208360 129792 208412
rect 273352 208360 273404 208412
rect 102232 208292 102284 208344
rect 262312 208292 262364 208344
rect 93124 207068 93176 207120
rect 96068 207068 96120 207120
rect 98644 207000 98696 207052
rect 102232 207000 102284 207052
rect 263692 207000 263744 207052
rect 196624 206932 196676 206984
rect 197268 206932 197320 206984
rect 269304 206932 269356 206984
rect 95240 206252 95292 206304
rect 122840 206252 122892 206304
rect 123760 206252 123812 206304
rect 123760 205640 123812 205692
rect 280160 205640 280212 205692
rect 280436 205640 280488 205692
rect 93860 204960 93912 205012
rect 103520 204960 103572 205012
rect 104716 204960 104768 205012
rect 84016 204892 84068 204944
rect 115204 204892 115256 204944
rect 225788 204892 225840 204944
rect 266544 204892 266596 204944
rect 104716 204348 104768 204400
rect 225144 204348 225196 204400
rect 225788 204348 225840 204400
rect 114652 204280 114704 204332
rect 115204 204280 115256 204332
rect 258080 204280 258132 204332
rect 267004 203600 267056 203652
rect 284484 203600 284536 203652
rect 200028 203532 200080 203584
rect 582472 203532 582524 203584
rect 99472 202784 99524 202836
rect 100116 202784 100168 202836
rect 111248 202784 111300 202836
rect 201592 202784 201644 202836
rect 202236 202784 202288 202836
rect 201408 202716 201460 202768
rect 224316 202716 224368 202768
rect 3240 202104 3292 202156
rect 99472 202104 99524 202156
rect 214656 202104 214708 202156
rect 222292 202104 222344 202156
rect 243544 202104 243596 202156
rect 280344 202104 280396 202156
rect 148416 201492 148468 201544
rect 152648 201492 152700 201544
rect 54852 201424 54904 201476
rect 55036 201424 55088 201476
rect 247684 201424 247736 201476
rect 96528 200744 96580 200796
rect 109684 200744 109736 200796
rect 244924 200744 244976 200796
rect 277584 200744 277636 200796
rect 74540 199452 74592 199504
rect 95884 199452 95936 199504
rect 52276 199384 52328 199436
rect 79416 199384 79468 199436
rect 117228 199384 117280 199436
rect 126336 199384 126388 199436
rect 153844 199384 153896 199436
rect 173348 199384 173400 199436
rect 193128 199384 193180 199436
rect 226432 199384 226484 199436
rect 256056 199384 256108 199436
rect 267924 199384 267976 199436
rect 162584 198636 162636 198688
rect 291292 198636 291344 198688
rect 53472 198568 53524 198620
rect 169760 198568 169812 198620
rect 162124 198228 162176 198280
rect 162584 198228 162636 198280
rect 92388 197956 92440 198008
rect 125600 197956 125652 198008
rect 176108 197956 176160 198008
rect 196624 197956 196676 198008
rect 169760 197888 169812 197940
rect 171048 197888 171100 197940
rect 171876 197888 171928 197940
rect 195244 196596 195296 196648
rect 226340 196596 226392 196648
rect 49608 195236 49660 195288
rect 130476 195236 130528 195288
rect 204996 195236 205048 195288
rect 260840 195236 260892 195288
rect 87696 193808 87748 193860
rect 102784 193808 102836 193860
rect 111156 193808 111208 193860
rect 151268 193808 151320 193860
rect 195244 193808 195296 193860
rect 287152 193808 287204 193860
rect 27528 192448 27580 192500
rect 138756 192448 138808 192500
rect 195336 192448 195388 192500
rect 243636 192448 243688 192500
rect 246304 192448 246356 192500
rect 580172 192448 580224 192500
rect 184756 191088 184808 191140
rect 226984 191088 227036 191140
rect 213184 189728 213236 189780
rect 265072 189728 265124 189780
rect 3424 188844 3476 188896
rect 7656 188844 7708 188896
rect 194508 188300 194560 188352
rect 223580 188300 223632 188352
rect 231124 188300 231176 188352
rect 263784 188300 263836 188352
rect 60556 187688 60608 187740
rect 186228 187620 186280 187672
rect 232504 187620 232556 187672
rect 44088 186260 44140 186312
rect 292580 186260 292632 186312
rect 90916 184152 90968 184204
rect 121552 184152 121604 184204
rect 193496 184152 193548 184204
rect 225972 184152 226024 184204
rect 183468 182792 183520 182844
rect 295340 182792 295392 182844
rect 181536 181500 181588 181552
rect 201500 181500 201552 181552
rect 84108 181432 84160 181484
rect 106464 181432 106516 181484
rect 198096 181432 198148 181484
rect 244924 181432 244976 181484
rect 12348 180072 12400 180124
rect 153936 180072 153988 180124
rect 206284 180072 206336 180124
rect 226524 180072 226576 180124
rect 87604 178644 87656 178696
rect 120080 178644 120132 178696
rect 236736 178644 236788 178696
rect 237288 178644 237340 178696
rect 580172 178644 580224 178696
rect 95976 178032 96028 178084
rect 101496 178032 101548 178084
rect 88248 177284 88300 177336
rect 204904 177284 204956 177336
rect 209964 177284 210016 177336
rect 274732 177284 274784 177336
rect 87604 176672 87656 176724
rect 88248 176672 88300 176724
rect 91192 176672 91244 176724
rect 220820 176672 220872 176724
rect 221464 176672 221516 176724
rect 222844 176332 222896 176384
rect 224960 176332 225012 176384
rect 88984 175924 89036 175976
rect 105544 175924 105596 175976
rect 117964 175244 118016 175296
rect 213276 175244 213328 175296
rect 203524 174496 203576 174548
rect 281632 174496 281684 174548
rect 306380 174496 306432 174548
rect 89720 173884 89772 173936
rect 90824 173884 90876 173936
rect 220084 173884 220136 173936
rect 223580 173000 223632 173052
rect 224316 173000 224368 173052
rect 145656 172592 145708 172644
rect 223580 172592 223632 172644
rect 89168 172524 89220 172576
rect 201500 172524 201552 172576
rect 253204 172524 253256 172576
rect 583024 172524 583076 172576
rect 194784 172456 194836 172508
rect 195336 172456 195388 172508
rect 189724 171844 189776 171896
rect 288716 171844 288768 171896
rect 56416 171776 56468 171828
rect 194784 171776 194836 171828
rect 201500 171028 201552 171080
rect 269120 171028 269172 171080
rect 76656 170348 76708 170400
rect 202972 170348 203024 170400
rect 203524 170348 203576 170400
rect 75920 169736 75972 169788
rect 76656 169736 76708 169788
rect 195980 168376 196032 168428
rect 196624 168376 196676 168428
rect 300124 168376 300176 168428
rect 177948 167628 178000 167680
rect 191196 167628 191248 167680
rect 215392 167628 215444 167680
rect 259552 167628 259604 167680
rect 135996 167016 136048 167068
rect 215300 167016 215352 167068
rect 186320 166336 186372 166388
rect 187608 166336 187660 166388
rect 198096 166336 198148 166388
rect 82912 166268 82964 166320
rect 177856 166268 177908 166320
rect 207664 166268 207716 166320
rect 63316 165588 63368 165640
rect 186320 165588 186372 165640
rect 215300 164840 215352 164892
rect 231860 164840 231912 164892
rect 123484 164296 123536 164348
rect 233240 164296 233292 164348
rect 86960 164228 87012 164280
rect 215944 164228 215996 164280
rect 60464 164160 60516 164212
rect 60648 164160 60700 164212
rect 189080 164160 189132 164212
rect 189724 164160 189776 164212
rect 200120 163888 200172 163940
rect 204996 163888 205048 163940
rect 60464 163480 60516 163532
rect 189080 163480 189132 163532
rect 222200 163480 222252 163532
rect 276020 163480 276072 163532
rect 87144 162868 87196 162920
rect 215392 162868 215444 162920
rect 236000 162800 236052 162852
rect 236736 162800 236788 162852
rect 247132 162120 247184 162172
rect 280528 162120 280580 162172
rect 340144 162120 340196 162172
rect 183008 161508 183060 161560
rect 236000 161508 236052 161560
rect 147036 161440 147088 161492
rect 224960 161440 225012 161492
rect 191932 161372 191984 161424
rect 247132 161372 247184 161424
rect 91008 160692 91060 160744
rect 109040 160692 109092 160744
rect 220176 160692 220228 160744
rect 183468 160080 183520 160132
rect 184204 160080 184256 160132
rect 191656 160080 191708 160132
rect 191932 160080 191984 160132
rect 220360 160080 220412 160132
rect 302240 160080 302292 160132
rect 208584 159332 208636 159384
rect 270592 159332 270644 159384
rect 255412 158924 255464 158976
rect 255964 158924 256016 158976
rect 88984 158788 89036 158840
rect 127716 158788 127768 158840
rect 153936 158788 153988 158840
rect 255412 158788 255464 158840
rect 64696 158720 64748 158772
rect 193128 158720 193180 158772
rect 75276 157972 75328 158024
rect 89168 157972 89220 158024
rect 127716 157972 127768 158024
rect 220820 157972 220872 158024
rect 61936 157360 61988 157412
rect 191748 157360 191800 157412
rect 214564 157360 214616 157412
rect 215116 157360 215168 157412
rect 582748 157360 582800 157412
rect 65984 156612 66036 156664
rect 163596 156612 163648 156664
rect 209872 156408 209924 156460
rect 210424 156408 210476 156460
rect 152648 156000 152700 156052
rect 256976 156000 257028 156052
rect 210424 155932 210476 155984
rect 582380 155932 582432 155984
rect 191564 155864 191616 155916
rect 191748 155864 191800 155916
rect 230480 155864 230532 155916
rect 231768 155864 231820 155916
rect 231768 155252 231820 155304
rect 243636 155252 243688 155304
rect 37096 155184 37148 155236
rect 48136 155184 48188 155236
rect 97264 155116 97316 155168
rect 97816 155116 97868 155168
rect 249800 155184 249852 155236
rect 250536 155184 250588 155236
rect 48136 154572 48188 154624
rect 186964 154572 187016 154624
rect 164240 154504 164292 154556
rect 165068 154504 165120 154556
rect 193128 154504 193180 154556
rect 218060 154504 218112 154556
rect 61660 153824 61712 153876
rect 75184 153824 75236 153876
rect 65892 153280 65944 153332
rect 165068 153280 165120 153332
rect 93860 153212 93912 153264
rect 95056 153212 95108 153264
rect 223580 153212 223632 153264
rect 239956 153212 240008 153264
rect 333980 153212 334032 153264
rect 60648 152532 60700 152584
rect 82084 152532 82136 152584
rect 207020 152532 207072 152584
rect 220360 152532 220412 152584
rect 64604 152464 64656 152516
rect 64788 152464 64840 152516
rect 190460 152464 190512 152516
rect 191104 152464 191156 152516
rect 191196 152464 191248 152516
rect 239956 152464 240008 152516
rect 161480 151784 161532 151836
rect 162584 151784 162636 151836
rect 185768 151784 185820 151836
rect 281448 151716 281500 151768
rect 291476 151716 291528 151768
rect 81992 151036 82044 151088
rect 104900 151036 104952 151088
rect 199292 151036 199344 151088
rect 263968 151036 264020 151088
rect 61752 150424 61804 150476
rect 62028 150424 62080 150476
rect 131856 150492 131908 150544
rect 126888 150424 126940 150476
rect 216680 150424 216732 150476
rect 201408 149676 201460 149728
rect 271880 149676 271932 149728
rect 218060 149268 218112 149320
rect 218612 149268 218664 149320
rect 73068 149132 73120 149184
rect 199292 149132 199344 149184
rect 55036 149064 55088 149116
rect 181444 149064 181496 149116
rect 204536 149064 204588 149116
rect 244924 149064 244976 149116
rect 53748 148316 53800 148368
rect 182824 148316 182876 148368
rect 184664 148316 184716 148368
rect 191840 148316 191892 148368
rect 206928 147704 206980 147756
rect 232504 147704 232556 147756
rect 98736 147636 98788 147688
rect 99288 147636 99340 147688
rect 224960 147636 225012 147688
rect 207664 147568 207716 147620
rect 211160 147568 211212 147620
rect 227812 147160 227864 147212
rect 192484 147024 192536 147076
rect 215484 147024 215536 147076
rect 3424 146956 3476 147008
rect 88248 146956 88300 147008
rect 108488 146956 108540 147008
rect 108948 146956 109000 147008
rect 197912 146956 197964 147008
rect 208400 146956 208452 147008
rect 208860 146956 208912 147008
rect 209872 146956 209924 147008
rect 210700 146956 210752 147008
rect 215392 146956 215444 147008
rect 216220 146956 216272 147008
rect 223580 146956 223632 147008
rect 224500 146956 224552 147008
rect 227720 146956 227772 147008
rect 57796 146888 57848 146940
rect 181536 146888 181588 146940
rect 213460 146888 213512 146940
rect 257988 146888 258040 146940
rect 258816 146888 258868 146940
rect 252468 146276 252520 146328
rect 341524 146276 341576 146328
rect 87512 146208 87564 146260
rect 88248 146208 88300 146260
rect 126888 146208 126940 146260
rect 184296 146208 184348 146260
rect 184848 146208 184900 146260
rect 220176 146208 220228 146260
rect 220912 146208 220964 146260
rect 192576 145528 192628 145580
rect 245108 145528 245160 145580
rect 338120 145528 338172 145580
rect 67364 144916 67416 144968
rect 109776 144916 109828 144968
rect 184296 144916 184348 144968
rect 217232 144916 217284 144968
rect 80152 144780 80204 144832
rect 83464 144780 83516 144832
rect 85580 144440 85632 144492
rect 89076 144440 89128 144492
rect 240784 144168 240836 144220
rect 258724 144168 258776 144220
rect 286784 144168 286836 144220
rect 295340 144168 295392 144220
rect 97356 144032 97408 144084
rect 99380 144032 99432 144084
rect 82820 143692 82872 143744
rect 86316 143692 86368 143744
rect 161480 143624 161532 143676
rect 162676 143624 162728 143676
rect 194140 143624 194192 143676
rect 204996 143624 205048 143676
rect 209780 143624 209832 143676
rect 63132 143556 63184 143608
rect 182916 143556 182968 143608
rect 187148 143556 187200 143608
rect 225236 143556 225288 143608
rect 219532 143488 219584 143540
rect 220268 143488 220320 143540
rect 220084 143420 220136 143472
rect 240784 143488 240836 143540
rect 214012 143216 214064 143268
rect 215116 143216 215168 143268
rect 53564 142808 53616 142860
rect 223672 142808 223724 142860
rect 245016 142808 245068 142860
rect 69020 142740 69072 142792
rect 70584 142740 70636 142792
rect 223212 142536 223264 142588
rect 223672 142536 223724 142588
rect 57704 142332 57756 142384
rect 89904 142332 89956 142384
rect 88616 142264 88668 142316
rect 218244 142264 218296 142316
rect 90916 142196 90968 142248
rect 213460 142196 213512 142248
rect 215300 142128 215352 142180
rect 223488 142128 223540 142180
rect 63408 141380 63460 141432
rect 77300 141380 77352 141432
rect 88524 141380 88576 141432
rect 184296 141380 184348 141432
rect 223028 140972 223080 141024
rect 227996 140972 228048 141024
rect 21364 140768 21416 140820
rect 88984 140768 89036 140820
rect 193312 140768 193364 140820
rect 196624 140768 196676 140820
rect 203432 140768 203484 140820
rect 289084 140768 289136 140820
rect 223488 140700 223540 140752
rect 251824 140700 251876 140752
rect 193036 140428 193088 140480
rect 194784 140428 194836 140480
rect 78036 140020 78088 140072
rect 87604 140020 87656 140072
rect 89904 139476 89956 139528
rect 96160 139476 96212 139528
rect 86868 139408 86920 139460
rect 84752 139340 84804 139392
rect 90916 139340 90968 139392
rect 205180 140496 205232 140548
rect 210056 140496 210108 140548
rect 215392 140428 215444 140480
rect 287704 140020 287756 140072
rect 251272 139748 251324 139800
rect 251824 139748 251876 139800
rect 193404 138660 193456 138712
rect 225328 138932 225380 138984
rect 227720 138932 227772 138984
rect 70216 138116 70268 138168
rect 71872 138116 71924 138168
rect 70400 138048 70452 138100
rect 71228 138048 71280 138100
rect 73344 138048 73396 138100
rect 73804 138048 73856 138100
rect 88340 138048 88392 138100
rect 89260 138048 89312 138100
rect 67916 137980 67968 138032
rect 159456 137980 159508 138032
rect 3240 137912 3292 137964
rect 73068 137844 73120 137896
rect 88984 137708 89036 137760
rect 91192 137708 91244 137760
rect 173348 137232 173400 137284
rect 183008 137232 183060 137284
rect 79968 136824 80020 136876
rect 80980 136824 81032 136876
rect 76564 136688 76616 136740
rect 77392 136688 77444 136740
rect 85488 136688 85540 136740
rect 86224 136688 86276 136740
rect 66076 136620 66128 136672
rect 94504 136620 94556 136672
rect 182824 136620 182876 136672
rect 191656 136620 191708 136672
rect 173808 136552 173860 136604
rect 191748 136552 191800 136604
rect 54484 135940 54536 135992
rect 90824 135940 90876 135992
rect 91284 135940 91336 135992
rect 64788 135872 64840 135924
rect 69664 135872 69716 135924
rect 70308 135872 70360 135924
rect 161480 135872 161532 135924
rect 226524 135872 226576 135924
rect 239404 135872 239456 135924
rect 243636 135872 243688 135924
rect 304264 135872 304316 135924
rect 226524 135600 226576 135652
rect 230480 135600 230532 135652
rect 160744 135260 160796 135312
rect 191748 135260 191800 135312
rect 94504 135192 94556 135244
rect 192484 135192 192536 135244
rect 232504 135192 232556 135244
rect 249064 135192 249116 135244
rect 96804 135124 96856 135176
rect 188528 135124 188580 135176
rect 93768 134580 93820 134632
rect 95240 134580 95292 134632
rect 247684 134512 247736 134564
rect 298744 134512 298796 134564
rect 96620 133832 96672 133884
rect 102876 133832 102928 133884
rect 188436 133832 188488 133884
rect 191748 133832 191800 133884
rect 226708 133832 226760 133884
rect 229284 133832 229336 133884
rect 226892 133764 226944 133816
rect 227904 133764 227956 133816
rect 268016 133832 268068 133884
rect 103060 133220 103112 133272
rect 160836 133220 160888 133272
rect 56416 133152 56468 133204
rect 66352 133152 66404 133204
rect 110880 133152 110932 133204
rect 187148 133152 187200 133204
rect 50988 132404 51040 132456
rect 66904 132404 66956 132456
rect 96160 132404 96212 132456
rect 191196 132404 191248 132456
rect 226708 132404 226760 132456
rect 229100 132404 229152 132456
rect 96620 132336 96672 132388
rect 148508 132336 148560 132388
rect 187608 131452 187660 131504
rect 192944 131452 192996 131504
rect 165068 131044 165120 131096
rect 182824 131044 182876 131096
rect 225420 131044 225472 131096
rect 273260 131044 273312 131096
rect 226616 130976 226668 131028
rect 256700 130976 256752 131028
rect 96620 130364 96672 130416
rect 170588 130364 170640 130416
rect 96620 130160 96672 130212
rect 102968 130160 103020 130212
rect 127716 129888 127768 129940
rect 133144 129888 133196 129940
rect 186320 129752 186372 129804
rect 191012 129752 191064 129804
rect 159456 129684 159508 129736
rect 185492 129684 185544 129736
rect 185676 129684 185728 129736
rect 227168 129276 227220 129328
rect 227996 129276 228048 129328
rect 104348 129004 104400 129056
rect 191472 129004 191524 129056
rect 192576 129004 192628 129056
rect 230388 129004 230440 129056
rect 249800 129004 249852 129056
rect 187608 128392 187660 128444
rect 189080 128392 189132 128444
rect 191196 128392 191248 128444
rect 226156 128324 226208 128376
rect 299480 128324 299532 128376
rect 48136 128256 48188 128308
rect 66904 128256 66956 128308
rect 97540 128256 97592 128308
rect 127808 128256 127860 128308
rect 163596 128256 163648 128308
rect 191748 128256 191800 128308
rect 226616 128256 226668 128308
rect 231860 128256 231912 128308
rect 233148 128256 233200 128308
rect 227996 127644 228048 127696
rect 267832 127644 267884 127696
rect 97080 127576 97132 127628
rect 183100 127576 183152 127628
rect 233148 127576 233200 127628
rect 331864 127576 331916 127628
rect 57612 126896 57664 126948
rect 66812 126896 66864 126948
rect 97816 126896 97868 126948
rect 110880 126896 110932 126948
rect 226432 126896 226484 126948
rect 255412 126896 255464 126948
rect 63316 126828 63368 126880
rect 66720 126828 66772 126880
rect 226892 126828 226944 126880
rect 227536 126828 227588 126880
rect 230388 126828 230440 126880
rect 126336 126284 126388 126336
rect 141608 126284 141660 126336
rect 108396 126216 108448 126268
rect 191656 126216 191708 126268
rect 193404 126216 193456 126268
rect 98460 125536 98512 125588
rect 152648 125536 152700 125588
rect 166356 125536 166408 125588
rect 186320 125536 186372 125588
rect 226616 125536 226668 125588
rect 259460 125536 259512 125588
rect 115204 124856 115256 124908
rect 127624 124856 127676 124908
rect 60464 124788 60516 124840
rect 66628 124788 66680 124840
rect 57704 124108 57756 124160
rect 66260 124108 66312 124160
rect 97816 124108 97868 124160
rect 147036 124108 147088 124160
rect 180064 124108 180116 124160
rect 191012 124108 191064 124160
rect 226708 124108 226760 124160
rect 233240 124108 233292 124160
rect 288532 124108 288584 124160
rect 582932 124108 582984 124160
rect 97172 124040 97224 124092
rect 135996 124040 136048 124092
rect 226524 123836 226576 123888
rect 229192 123836 229244 123888
rect 162124 123428 162176 123480
rect 173256 123428 173308 123480
rect 97540 122748 97592 122800
rect 153936 122748 153988 122800
rect 226524 122748 226576 122800
rect 236000 122748 236052 122800
rect 181536 122068 181588 122120
rect 181996 122068 182048 122120
rect 191748 122068 191800 122120
rect 226984 122068 227036 122120
rect 309784 122068 309836 122120
rect 54944 121388 54996 121440
rect 66904 121388 66956 121440
rect 96988 121388 97040 121440
rect 103060 121388 103112 121440
rect 185768 121388 185820 121440
rect 191748 121388 191800 121440
rect 226708 121388 226760 121440
rect 240140 121388 240192 121440
rect 61936 121320 61988 121372
rect 66812 121320 66864 121372
rect 110328 120776 110380 120828
rect 142988 120776 143040 120828
rect 108396 120708 108448 120760
rect 124864 120708 124916 120760
rect 131856 120708 131908 120760
rect 187700 120708 187752 120760
rect 239404 120708 239456 120760
rect 282184 120708 282236 120760
rect 96068 120300 96120 120352
rect 98828 120300 98880 120352
rect 187700 120164 187752 120216
rect 188988 120164 189040 120216
rect 191748 120164 191800 120216
rect 53656 120028 53708 120080
rect 66904 120028 66956 120080
rect 97908 120028 97960 120080
rect 123484 120028 123536 120080
rect 181444 120028 181496 120080
rect 191748 120028 191800 120080
rect 64696 119960 64748 120012
rect 66812 119960 66864 120012
rect 109684 118668 109736 118720
rect 173808 118668 173860 118720
rect 174636 118668 174688 118720
rect 57796 118600 57848 118652
rect 66720 118600 66772 118652
rect 97908 118600 97960 118652
rect 173348 118600 173400 118652
rect 181996 118600 182048 118652
rect 184204 118600 184256 118652
rect 181996 117920 182048 117972
rect 191012 117920 191064 117972
rect 227536 117920 227588 117972
rect 353300 117920 353352 117972
rect 99380 117308 99432 117360
rect 100668 117308 100720 117360
rect 108488 117308 108540 117360
rect 226616 117308 226668 117360
rect 252744 117308 252796 117360
rect 64512 117240 64564 117292
rect 66812 117240 66864 117292
rect 97908 117240 97960 117292
rect 177396 117240 177448 117292
rect 182916 117240 182968 117292
rect 191748 117240 191800 117292
rect 61752 117172 61804 117224
rect 66260 117172 66312 117224
rect 97356 117172 97408 117224
rect 155408 117172 155460 117224
rect 188344 117172 188396 117224
rect 191012 117172 191064 117224
rect 226708 116968 226760 117020
rect 230480 116968 230532 117020
rect 231124 116968 231176 117020
rect 230388 116628 230440 116680
rect 262220 116628 262272 116680
rect 231124 116560 231176 116612
rect 281540 116560 281592 116612
rect 304356 116560 304408 116612
rect 226708 115948 226760 116000
rect 229100 115948 229152 116000
rect 230388 115948 230440 116000
rect 55036 115880 55088 115932
rect 66904 115880 66956 115932
rect 97816 115880 97868 115932
rect 99380 115880 99432 115932
rect 180708 115880 180760 115932
rect 190828 115880 190880 115932
rect 64604 115268 64656 115320
rect 66812 115268 66864 115320
rect 233240 115200 233292 115252
rect 277400 115200 277452 115252
rect 97908 114520 97960 114572
rect 169116 114520 169168 114572
rect 226708 114520 226760 114572
rect 233240 114520 233292 114572
rect 8208 114452 8260 114504
rect 59176 114452 59228 114504
rect 66812 114452 66864 114504
rect 226616 114452 226668 114504
rect 242256 114452 242308 114504
rect 250536 114452 250588 114504
rect 63132 114384 63184 114436
rect 66904 114384 66956 114436
rect 97816 113976 97868 114028
rect 101496 113976 101548 114028
rect 235264 113772 235316 113824
rect 242164 113772 242216 113824
rect 97908 113160 97960 113212
rect 173256 113160 173308 113212
rect 188252 113160 188304 113212
rect 191748 113160 191800 113212
rect 52368 112412 52420 112464
rect 66812 112412 66864 112464
rect 157248 112412 157300 112464
rect 191748 112412 191800 112464
rect 97080 111868 97132 111920
rect 100024 111868 100076 111920
rect 98092 111800 98144 111852
rect 100760 111800 100812 111852
rect 156696 111800 156748 111852
rect 157248 111800 157300 111852
rect 226708 111800 226760 111852
rect 231952 111800 232004 111852
rect 324320 111800 324372 111852
rect 3424 111732 3476 111784
rect 21364 111732 21416 111784
rect 96712 111664 96764 111716
rect 98736 111664 98788 111716
rect 239404 111120 239456 111172
rect 252652 111120 252704 111172
rect 41144 111052 41196 111104
rect 57152 111052 57204 111104
rect 101588 111052 101640 111104
rect 114652 111052 114704 111104
rect 227076 111052 227128 111104
rect 227720 111052 227772 111104
rect 242164 111052 242216 111104
rect 188896 110508 188948 110560
rect 191840 110508 191892 110560
rect 57152 110440 57204 110492
rect 57796 110440 57848 110492
rect 66812 110440 66864 110492
rect 97908 110372 97960 110424
rect 102048 110440 102100 110492
rect 186964 110440 187016 110492
rect 187700 110440 187752 110492
rect 191748 110440 191800 110492
rect 227720 110372 227772 110424
rect 228364 110372 228416 110424
rect 233884 110372 233936 110424
rect 100116 109692 100168 109744
rect 111800 109692 111852 109744
rect 160836 109692 160888 109744
rect 188252 109692 188304 109744
rect 236736 109692 236788 109744
rect 258080 109692 258132 109744
rect 50896 109012 50948 109064
rect 57244 109012 57296 109064
rect 66812 109012 66864 109064
rect 123484 109012 123536 109064
rect 156604 108944 156656 108996
rect 189080 108944 189132 108996
rect 226432 108944 226484 108996
rect 245660 108944 245712 108996
rect 97908 108332 97960 108384
rect 107476 108332 107528 108384
rect 108488 108332 108540 108384
rect 155408 108332 155460 108384
rect 44088 108264 44140 108316
rect 63500 108264 63552 108316
rect 101680 108264 101732 108316
rect 187700 108264 187752 108316
rect 231768 108264 231820 108316
rect 269212 108264 269264 108316
rect 63500 107652 63552 107704
rect 64604 107652 64656 107704
rect 66812 107652 66864 107704
rect 226708 107652 226760 107704
rect 230572 107652 230624 107704
rect 231768 107652 231820 107704
rect 171876 107584 171928 107636
rect 191748 107584 191800 107636
rect 226800 107584 226852 107636
rect 282920 107584 282972 107636
rect 7564 106904 7616 106956
rect 34336 106904 34388 106956
rect 60740 106904 60792 106956
rect 97816 106904 97868 106956
rect 180064 106904 180116 106956
rect 282920 106904 282972 106956
rect 342904 106904 342956 106956
rect 96712 106360 96764 106412
rect 98736 106360 98788 106412
rect 60740 106292 60792 106344
rect 61936 106292 61988 106344
rect 66812 106292 66864 106344
rect 109776 106224 109828 106276
rect 191196 106224 191248 106276
rect 46848 105544 46900 105596
rect 65892 105544 65944 105596
rect 66536 105544 66588 105596
rect 158076 105544 158128 105596
rect 190276 105544 190328 105596
rect 191748 105544 191800 105596
rect 226708 105544 226760 105596
rect 267004 105544 267056 105596
rect 112444 105340 112496 105392
rect 113272 105340 113324 105392
rect 53472 104796 53524 104848
rect 66812 104796 66864 104848
rect 96804 104116 96856 104168
rect 112444 104116 112496 104168
rect 130476 104116 130528 104168
rect 152556 104116 152608 104168
rect 233332 104116 233384 104168
rect 235908 104116 235960 104168
rect 305644 104116 305696 104168
rect 96528 103504 96580 103556
rect 183008 103504 183060 103556
rect 226708 103504 226760 103556
rect 233332 103504 233384 103556
rect 63224 103436 63276 103488
rect 66812 103436 66864 103488
rect 164148 103436 164200 103488
rect 193036 103436 193088 103488
rect 98000 102824 98052 102876
rect 166356 102824 166408 102876
rect 94596 102756 94648 102808
rect 164148 102756 164200 102808
rect 233148 102756 233200 102808
rect 278780 102756 278832 102808
rect 321652 102756 321704 102808
rect 182916 102212 182968 102264
rect 191748 102212 191800 102264
rect 226616 102212 226668 102264
rect 231860 102212 231912 102264
rect 233148 102212 233200 102264
rect 226708 102144 226760 102196
rect 237564 102144 237616 102196
rect 97908 102076 97960 102128
rect 129096 102076 129148 102128
rect 226524 102076 226576 102128
rect 266360 102076 266412 102128
rect 129096 101464 129148 101516
rect 162216 101464 162268 101516
rect 55128 101396 55180 101448
rect 66076 101396 66128 101448
rect 66628 101396 66680 101448
rect 98828 101396 98880 101448
rect 162768 101396 162820 101448
rect 191472 101396 191524 101448
rect 191748 101396 191800 101448
rect 186228 100648 186280 100700
rect 191748 100648 191800 100700
rect 178868 100036 178920 100088
rect 191104 100036 191156 100088
rect 57888 99968 57940 100020
rect 64696 99968 64748 100020
rect 66812 99968 66864 100020
rect 97908 99968 97960 100020
rect 101404 99968 101456 100020
rect 184296 99968 184348 100020
rect 226708 99424 226760 99476
rect 229192 99424 229244 99476
rect 245660 99424 245712 99476
rect 97540 99356 97592 99408
rect 133788 99356 133840 99408
rect 226616 99356 226668 99408
rect 320824 99356 320876 99408
rect 60556 99288 60608 99340
rect 66812 99288 66864 99340
rect 227352 98608 227404 98660
rect 236644 98608 236696 98660
rect 245660 98608 245712 98660
rect 277400 98608 277452 98660
rect 97816 98064 97868 98116
rect 106280 98064 106332 98116
rect 97908 97996 97960 98048
rect 152556 97996 152608 98048
rect 187516 97996 187568 98048
rect 190552 97996 190604 98048
rect 159548 97928 159600 97980
rect 190460 97928 190512 97980
rect 226248 97928 226300 97980
rect 237656 97928 237708 97980
rect 96712 97724 96764 97776
rect 98644 97724 98696 97776
rect 97816 97248 97868 97300
rect 129740 97248 129792 97300
rect 3424 96636 3476 96688
rect 61384 96636 61436 96688
rect 226708 96568 226760 96620
rect 262312 96568 262364 96620
rect 59084 95888 59136 95940
rect 66444 95888 66496 95940
rect 226892 95888 226944 95940
rect 273352 95888 273404 95940
rect 97080 95276 97132 95328
rect 100024 95276 100076 95328
rect 97908 95208 97960 95260
rect 188344 95208 188396 95260
rect 61844 95140 61896 95192
rect 66812 95140 66864 95192
rect 67548 95140 67600 95192
rect 68284 95140 68336 95192
rect 99012 94528 99064 94580
rect 166448 94528 166500 94580
rect 191472 94528 191524 94580
rect 191748 94528 191800 94580
rect 95516 94460 95568 94512
rect 177948 94460 178000 94512
rect 191840 94460 191892 94512
rect 170496 93848 170548 93900
rect 193404 93848 193456 93900
rect 67548 93780 67600 93832
rect 67916 93780 67968 93832
rect 97908 93780 97960 93832
rect 106372 93780 106424 93832
rect 186964 93780 187016 93832
rect 193220 93780 193272 93832
rect 191840 93372 191892 93424
rect 199108 93372 199160 93424
rect 221648 93372 221700 93424
rect 225144 93372 225196 93424
rect 193404 93304 193456 93356
rect 193772 93304 193824 93356
rect 168288 93168 168340 93220
rect 183560 93168 183612 93220
rect 190460 93168 190512 93220
rect 249156 93168 249208 93220
rect 264980 93168 265032 93220
rect 107476 93100 107528 93152
rect 170496 93100 170548 93152
rect 207664 93100 207716 93152
rect 225052 93100 225104 93152
rect 258816 93100 258868 93152
rect 316040 93100 316092 93152
rect 67640 92828 67692 92880
rect 68468 92828 68520 92880
rect 95240 92760 95292 92812
rect 71734 92692 71786 92744
rect 87558 92692 87610 92744
rect 93814 92692 93866 92744
rect 94688 92692 94740 92744
rect 59268 92556 59320 92608
rect 66996 92556 67048 92608
rect 67272 92556 67324 92608
rect 71780 92556 71832 92608
rect 74540 92556 74592 92608
rect 75782 92556 75834 92608
rect 81624 92556 81676 92608
rect 82590 92556 82642 92608
rect 86960 92556 87012 92608
rect 88110 92556 88162 92608
rect 89904 92556 89956 92608
rect 90686 92556 90738 92608
rect 94504 92488 94556 92540
rect 122840 92488 122892 92540
rect 56508 92420 56560 92472
rect 72792 92420 72844 92472
rect 75460 92420 75512 92472
rect 95884 92420 95936 92472
rect 184296 92420 184348 92472
rect 226616 92420 226668 92472
rect 60648 92352 60700 92404
rect 81440 92352 81492 92404
rect 92388 92352 92440 92404
rect 103520 92352 103572 92404
rect 205640 92352 205692 92404
rect 225236 92352 225288 92404
rect 193220 92080 193272 92132
rect 193772 92080 193824 92132
rect 112444 91740 112496 91792
rect 205640 91740 205692 91792
rect 245016 91740 245068 91792
rect 258724 91740 258776 91792
rect 104348 91060 104400 91112
rect 111064 91060 111116 91112
rect 63408 90992 63460 91044
rect 73712 90992 73764 91044
rect 112444 90992 112496 91044
rect 113180 90992 113232 91044
rect 179328 90992 179380 91044
rect 194692 90992 194744 91044
rect 195244 90992 195296 91044
rect 217324 90992 217376 91044
rect 296720 90992 296772 91044
rect 66168 90924 66220 90976
rect 70308 90924 70360 90976
rect 78956 90312 79008 90364
rect 96712 90312 96764 90364
rect 97264 90312 97316 90364
rect 105544 90312 105596 90364
rect 212908 90312 212960 90364
rect 242164 90312 242216 90364
rect 271144 90312 271196 90364
rect 70308 90244 70360 90296
rect 71044 90244 71096 90296
rect 223764 90244 223816 90296
rect 224868 90244 224920 90296
rect 204352 89768 204404 89820
rect 205548 89768 205600 89820
rect 124864 89700 124916 89752
rect 125600 89700 125652 89752
rect 204904 89700 204956 89752
rect 207940 89700 207992 89752
rect 67548 89632 67600 89684
rect 99012 89632 99064 89684
rect 61660 89564 61712 89616
rect 74816 89564 74868 89616
rect 89260 89564 89312 89616
rect 118700 89564 118752 89616
rect 217692 89632 217744 89684
rect 219992 89632 220044 89684
rect 277492 89632 277544 89684
rect 278688 89632 278740 89684
rect 125416 89564 125468 89616
rect 218244 89564 218296 89616
rect 278688 88952 278740 89004
rect 582380 88952 582432 89004
rect 52276 88272 52328 88324
rect 79416 88272 79468 88324
rect 87604 88272 87656 88324
rect 88156 88272 88208 88324
rect 121460 88272 121512 88324
rect 215392 88272 215444 88324
rect 73712 88204 73764 88256
rect 95516 88204 95568 88256
rect 205640 88204 205692 88256
rect 226432 88204 226484 88256
rect 100116 87592 100168 87644
rect 125416 87592 125468 87644
rect 164976 87592 165028 87644
rect 165528 87592 165580 87644
rect 206836 87592 206888 87644
rect 227536 87592 227588 87644
rect 241520 87592 241572 87644
rect 80060 86912 80112 86964
rect 165528 86912 165580 86964
rect 184664 86912 184716 86964
rect 199384 86912 199436 86964
rect 212908 86912 212960 86964
rect 213828 86912 213880 86964
rect 235264 86912 235316 86964
rect 259368 86912 259420 86964
rect 276664 86912 276716 86964
rect 580172 86912 580224 86964
rect 67364 86844 67416 86896
rect 98828 86844 98880 86896
rect 199476 86232 199528 86284
rect 244280 86232 244332 86284
rect 3148 85484 3200 85536
rect 57244 85484 57296 85536
rect 160836 85484 160888 85536
rect 220636 85484 220688 85536
rect 263692 85484 263744 85536
rect 69204 85416 69256 85468
rect 107476 85416 107528 85468
rect 108120 85416 108172 85468
rect 204996 85416 205048 85468
rect 242808 85416 242860 85468
rect 243544 85416 243596 85468
rect 206836 84804 206888 84856
rect 220084 84804 220136 84856
rect 216036 84192 216088 84244
rect 242808 84192 242860 84244
rect 67824 84124 67876 84176
rect 94596 84124 94648 84176
rect 104164 84124 104216 84176
rect 213920 84124 213972 84176
rect 70400 84056 70452 84108
rect 169668 84056 169720 84108
rect 195980 84056 196032 84108
rect 209872 84056 209924 84108
rect 210424 84056 210476 84108
rect 275008 84056 275060 84108
rect 275008 83444 275060 83496
rect 322940 83444 322992 83496
rect 195980 82832 196032 82884
rect 196624 82832 196676 82884
rect 75920 82764 75972 82816
rect 102784 82764 102836 82816
rect 115296 82764 115348 82816
rect 224960 82764 225012 82816
rect 84200 82696 84252 82748
rect 105544 82696 105596 82748
rect 155408 82696 155460 82748
rect 252744 82696 252796 82748
rect 252744 81404 252796 81456
rect 253204 81404 253256 81456
rect 80152 81336 80204 81388
rect 112444 81336 112496 81388
rect 183008 81336 183060 81388
rect 233332 81336 233384 81388
rect 89720 81268 89772 81320
rect 100116 81268 100168 81320
rect 173808 81268 173860 81320
rect 204904 81268 204956 81320
rect 262128 80044 262180 80096
rect 263600 80044 263652 80096
rect 81716 79976 81768 80028
rect 112536 79976 112588 80028
rect 169116 79976 169168 80028
rect 230480 79976 230532 80028
rect 204168 79908 204220 79960
rect 237380 79908 237432 79960
rect 203524 79500 203576 79552
rect 204168 79500 204220 79552
rect 90364 79296 90416 79348
rect 134616 79296 134668 79348
rect 64696 78616 64748 78668
rect 191564 78616 191616 78668
rect 248420 78616 248472 78668
rect 249156 78616 249208 78668
rect 82820 78548 82872 78600
rect 181260 78548 181312 78600
rect 190184 77936 190236 77988
rect 214656 77936 214708 77988
rect 88340 77188 88392 77240
rect 121552 77188 121604 77240
rect 133788 77188 133840 77240
rect 229192 77188 229244 77240
rect 3148 76508 3200 76560
rect 95332 76508 95384 76560
rect 200212 76508 200264 76560
rect 245660 76508 245712 76560
rect 121552 76440 121604 76492
rect 122104 76440 122156 76492
rect 57796 75828 57848 75880
rect 188896 75828 188948 75880
rect 263600 75828 263652 75880
rect 65616 75760 65668 75812
rect 66076 75760 66128 75812
rect 182916 75760 182968 75812
rect 81624 74468 81676 74520
rect 106464 74468 106516 74520
rect 210424 74468 210476 74520
rect 212632 74468 212684 74520
rect 269764 74468 269816 74520
rect 57888 73788 57940 73840
rect 185584 73788 185636 73840
rect 212632 73176 212684 73228
rect 213184 73176 213236 73228
rect 86960 73108 87012 73160
rect 215300 73108 215352 73160
rect 162216 73040 162268 73092
rect 237564 73040 237616 73092
rect 215300 71748 215352 71800
rect 215944 71748 215996 71800
rect 237564 71748 237616 71800
rect 238024 71748 238076 71800
rect 61936 71680 61988 71732
rect 178868 71680 178920 71732
rect 180064 71680 180116 71732
rect 228364 71680 228416 71732
rect 124864 71612 124916 71664
rect 218060 71612 218112 71664
rect 218336 71612 218388 71664
rect 88248 71000 88300 71052
rect 111156 71000 111208 71052
rect 218336 71000 218388 71052
rect 351920 71000 351972 71052
rect 94504 70320 94556 70372
rect 222292 70320 222344 70372
rect 222844 70320 222896 70372
rect 71688 69640 71740 69692
rect 171784 69640 171836 69692
rect 193128 69640 193180 69692
rect 270500 69640 270552 69692
rect 69204 68960 69256 69012
rect 194784 68960 194836 69012
rect 195336 68960 195388 69012
rect 89628 68280 89680 68332
rect 163504 68280 163556 68332
rect 192852 68280 192904 68332
rect 281540 68280 281592 68332
rect 71872 67532 71924 67584
rect 197360 67532 197412 67584
rect 198004 67532 198056 67584
rect 201500 67532 201552 67584
rect 202144 67532 202196 67584
rect 293960 67532 294012 67584
rect 166356 67464 166408 67516
rect 231860 67464 231912 67516
rect 100024 66172 100076 66224
rect 241520 66172 241572 66224
rect 75828 65492 75880 65544
rect 177304 65492 177356 65544
rect 187608 65492 187660 65544
rect 214564 65492 214616 65544
rect 85580 64812 85632 64864
rect 118792 64812 118844 64864
rect 213184 64812 213236 64864
rect 152556 64744 152608 64796
rect 227720 64744 227772 64796
rect 106188 64132 106240 64184
rect 126336 64132 126388 64184
rect 227720 63520 227772 63572
rect 228364 63520 228416 63572
rect 193312 63452 193364 63504
rect 295432 63452 295484 63504
rect 122104 63384 122156 63436
rect 217324 63384 217376 63436
rect 85488 62840 85540 62892
rect 115204 62840 115256 62892
rect 81348 62772 81400 62824
rect 130476 62772 130528 62824
rect 88156 62024 88208 62076
rect 216036 62024 216088 62076
rect 71044 61956 71096 62008
rect 194692 61956 194744 62008
rect 195336 61956 195388 62008
rect 285680 61956 285732 62008
rect 286600 61956 286652 62008
rect 286600 61344 286652 61396
rect 345020 61344 345072 61396
rect 194692 60732 194744 60784
rect 195244 60732 195296 60784
rect 67272 60664 67324 60716
rect 183560 60664 183612 60716
rect 184296 60664 184348 60716
rect 97264 60596 97316 60648
rect 204352 60596 204404 60648
rect 204352 60188 204404 60240
rect 204996 60188 205048 60240
rect 193220 59984 193272 60036
rect 264980 59984 265032 60036
rect 3056 59304 3108 59356
rect 51724 59304 51776 59356
rect 67640 59304 67692 59356
rect 193312 59304 193364 59356
rect 193864 59304 193916 59356
rect 112444 59236 112496 59288
rect 207112 59304 207164 59356
rect 207664 59304 207716 59356
rect 200120 59168 200172 59220
rect 289820 59304 289872 59356
rect 93768 57876 93820 57928
rect 222200 57876 222252 57928
rect 222936 57876 222988 57928
rect 73804 57808 73856 57860
rect 200120 57808 200172 57860
rect 200764 57808 200816 57860
rect 74540 56516 74592 56568
rect 202144 56516 202196 56568
rect 198004 56448 198056 56500
rect 247040 56448 247092 56500
rect 247592 56448 247644 56500
rect 247592 55836 247644 55888
rect 342260 55836 342312 55888
rect 103336 54544 103388 54596
rect 133236 54544 133288 54596
rect 73068 54476 73120 54528
rect 145564 54476 145616 54528
rect 184296 54476 184348 54528
rect 320180 54476 320232 54528
rect 97264 53048 97316 53100
rect 141516 53048 141568 53100
rect 214656 53048 214708 53100
rect 286324 53048 286376 53100
rect 61936 51688 61988 51740
rect 144184 51688 144236 51740
rect 186964 51688 187016 51740
rect 580172 51688 580224 51740
rect 3976 50328 4028 50380
rect 142896 50328 142948 50380
rect 182824 50328 182876 50380
rect 335360 50328 335412 50380
rect 59268 48968 59320 49020
rect 151176 48968 151228 49020
rect 193036 48968 193088 49020
rect 310520 48968 310572 49020
rect 65524 47540 65576 47592
rect 149704 47540 149756 47592
rect 181996 47540 182048 47592
rect 226984 47540 227036 47592
rect 119896 46248 119948 46300
rect 153844 46248 153896 46300
rect 3332 46180 3384 46232
rect 65616 46180 65668 46232
rect 67548 46180 67600 46232
rect 129004 46180 129056 46232
rect 217324 46180 217376 46232
rect 291936 46180 291988 46232
rect 190276 44820 190328 44872
rect 288440 44820 288492 44872
rect 77208 43392 77260 43444
rect 146944 43392 146996 43444
rect 191656 43392 191708 43444
rect 305736 43392 305788 43444
rect 79324 42032 79376 42084
rect 137376 42032 137428 42084
rect 305644 42032 305696 42084
rect 329840 42032 329892 42084
rect 99288 40672 99340 40724
rect 162124 40672 162176 40724
rect 239404 40672 239456 40724
rect 349804 40672 349856 40724
rect 82728 39312 82780 39364
rect 167644 39312 167696 39364
rect 199384 39312 199436 39364
rect 233884 39312 233936 39364
rect 244924 37952 244976 38004
rect 258816 37952 258868 38004
rect 68928 37884 68980 37936
rect 174544 37884 174596 37936
rect 184204 37884 184256 37936
rect 249800 37884 249852 37936
rect 67732 36524 67784 36576
rect 125600 36524 125652 36576
rect 214564 36524 214616 36576
rect 327080 36524 327132 36576
rect 75184 35164 75236 35216
rect 155316 35164 155368 35216
rect 222936 35164 222988 35216
rect 301504 35164 301556 35216
rect 55128 33736 55180 33788
rect 140044 33736 140096 33788
rect 200764 33736 200816 33788
rect 340972 33736 341024 33788
rect 3516 33056 3568 33108
rect 54484 33056 54536 33108
rect 64788 32376 64840 32428
rect 175924 32376 175976 32428
rect 44088 31016 44140 31068
rect 169024 31016 169076 31068
rect 195244 31016 195296 31068
rect 311900 31016 311952 31068
rect 46848 29588 46900 29640
rect 166264 29588 166316 29640
rect 193864 29588 193916 29640
rect 291200 29588 291252 29640
rect 291844 29588 291896 29640
rect 325700 29588 325752 29640
rect 86776 28228 86828 28280
rect 164884 28228 164936 28280
rect 213184 28228 213236 28280
rect 287060 28228 287112 28280
rect 93768 26868 93820 26920
rect 157984 26868 158036 26920
rect 56508 25508 56560 25560
rect 135904 25508 135956 25560
rect 209688 25508 209740 25560
rect 278780 25508 278832 25560
rect 66168 24080 66220 24132
rect 138664 24080 138716 24132
rect 207664 24080 207716 24132
rect 246304 24080 246356 24132
rect 78588 22720 78640 22772
rect 178684 22720 178736 22772
rect 213828 22720 213880 22772
rect 334072 22720 334124 22772
rect 74448 21360 74500 21412
rect 108396 21360 108448 21412
rect 111616 21360 111668 21412
rect 127716 21360 127768 21412
rect 204168 21360 204220 21412
rect 324412 21360 324464 21412
rect 3424 20612 3476 20664
rect 93124 20612 93176 20664
rect 242808 20000 242860 20052
rect 284392 20000 284444 20052
rect 91008 19932 91060 19984
rect 141424 19932 141476 19984
rect 185676 19932 185728 19984
rect 242992 19932 243044 19984
rect 50988 18572 51040 18624
rect 170404 18572 170456 18624
rect 222844 18572 222896 18624
rect 339500 18572 339552 18624
rect 228364 17212 228416 17264
rect 331220 17212 331272 17264
rect 240784 15852 240836 15904
rect 253480 15852 253532 15904
rect 253204 15172 253256 15224
rect 256700 15172 256752 15224
rect 95056 14424 95108 14476
rect 152464 14424 152516 14476
rect 204996 14424 205048 14476
rect 344560 14424 344612 14476
rect 70216 13064 70268 13116
rect 142804 13064 142856 13116
rect 249064 13064 249116 13116
rect 302884 13064 302936 13116
rect 84108 11704 84160 11756
rect 131764 11704 131816 11756
rect 215944 11704 215996 11756
rect 266544 11704 266596 11756
rect 79692 10276 79744 10328
rect 148416 10276 148468 10328
rect 202144 10276 202196 10328
rect 321560 10276 321612 10328
rect 99840 8984 99892 9036
rect 173164 8984 173216 9036
rect 572 8916 624 8968
rect 101404 8916 101456 8968
rect 196624 8916 196676 8968
rect 258264 8916 258316 8968
rect 320824 8916 320876 8968
rect 332692 8916 332744 8968
rect 250536 7624 250588 7676
rect 261760 7624 261812 7676
rect 267004 7624 267056 7676
rect 276020 7624 276072 7676
rect 59636 7556 59688 7608
rect 155224 7556 155276 7608
rect 191748 7556 191800 7608
rect 249800 7556 249852 7608
rect 258724 7556 258776 7608
rect 269120 7556 269172 7608
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 52552 6128 52604 6180
rect 159364 6128 159416 6180
rect 224868 6128 224920 6180
rect 254676 6128 254728 6180
rect 271144 6128 271196 6180
rect 297272 6128 297324 6180
rect 305736 5516 305788 5568
rect 309048 5516 309100 5568
rect 349804 5516 349856 5568
rect 351644 5516 351696 5568
rect 96252 4836 96304 4888
rect 151084 4836 151136 4888
rect 1676 4768 1728 4820
rect 97264 4768 97316 4820
rect 204904 4768 204956 4820
rect 274824 4768 274876 4820
rect 331864 4496 331916 4548
rect 337476 4496 337528 4548
rect 238024 4360 238076 4412
rect 239312 4360 239364 4412
rect 134524 4156 134576 4208
rect 136456 4156 136508 4208
rect 342996 4088 343048 4140
rect 346952 4088 347004 4140
rect 233884 4020 233936 4072
rect 240508 4020 240560 4072
rect 44272 3884 44324 3936
rect 47584 3884 47636 3936
rect 304356 3748 304408 3800
rect 307944 3748 307996 3800
rect 27712 3612 27764 3664
rect 32404 3612 32456 3664
rect 60832 3544 60884 3596
rect 61936 3544 61988 3596
rect 101036 3544 101088 3596
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 19432 3476 19484 3528
rect 20628 3476 20680 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 44088 3476 44140 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 64328 3476 64380 3528
rect 64788 3476 64840 3528
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 69112 3476 69164 3528
rect 70216 3476 70268 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 73804 3476 73856 3528
rect 74448 3476 74500 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 80888 3476 80940 3528
rect 81348 3476 81400 3528
rect 82084 3476 82136 3528
rect 82728 3476 82780 3528
rect 83280 3476 83332 3528
rect 84108 3476 84160 3528
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 85672 3476 85724 3528
rect 86776 3476 86828 3528
rect 89168 3476 89220 3528
rect 89628 3476 89680 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 92756 3476 92808 3528
rect 93768 3476 93820 3528
rect 93952 3476 94004 3528
rect 95056 3476 95108 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 102232 3476 102284 3528
rect 103244 3476 103296 3528
rect 114008 3544 114060 3596
rect 114468 3544 114520 3596
rect 115204 3544 115256 3596
rect 115848 3544 115900 3596
rect 116400 3544 116452 3596
rect 117228 3544 117280 3596
rect 117596 3544 117648 3596
rect 118608 3544 118660 3596
rect 122288 3544 122340 3596
rect 122748 3544 122800 3596
rect 126244 3544 126296 3596
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 128268 3476 128320 3528
rect 129372 3476 129424 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 147128 3476 147180 3528
rect 147588 3476 147640 3528
rect 258816 3476 258868 3528
rect 260656 3476 260708 3528
rect 269120 3476 269172 3528
rect 272432 3476 272484 3528
rect 281448 3476 281500 3528
rect 286600 3476 286652 3528
rect 291936 3476 291988 3528
rect 294880 3476 294932 3528
rect 301504 3476 301556 3528
rect 303160 3476 303212 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 327080 3476 327132 3528
rect 328000 3476 328052 3528
rect 340144 3476 340196 3528
rect 342168 3476 342220 3528
rect 582196 3476 582248 3528
rect 583116 3476 583168 3528
rect 15936 3408 15988 3460
rect 43444 3408 43496 3460
rect 63224 3408 63276 3460
rect 75184 3408 75236 3460
rect 77392 3408 77444 3460
rect 90272 3408 90324 3460
rect 91560 3408 91612 3460
rect 104348 3408 104400 3460
rect 105728 3408 105780 3460
rect 106188 3408 106240 3460
rect 106924 3408 106976 3460
rect 107568 3408 107620 3460
rect 109316 3408 109368 3460
rect 110328 3408 110380 3460
rect 110512 3408 110564 3460
rect 111708 3408 111760 3460
rect 108120 3340 108172 3392
rect 137284 3408 137336 3460
rect 220084 3408 220136 3460
rect 242900 3408 242952 3460
rect 260104 3408 260156 3460
rect 267740 3408 267792 3460
rect 304264 3408 304316 3460
rect 310244 3408 310296 3460
rect 327724 3408 327776 3460
rect 329196 3408 329248 3460
rect 341524 3408 341576 3460
rect 350448 3408 350500 3460
rect 287704 3340 287756 3392
rect 290188 3340 290240 3392
rect 20628 3272 20680 3324
rect 25504 3272 25556 3324
rect 249800 3272 249852 3324
rect 251180 3272 251232 3324
rect 298744 3272 298796 3324
rect 301964 3272 302016 3324
rect 317328 3272 317380 3324
rect 321652 3272 321704 3324
rect 76196 3204 76248 3256
rect 77208 3204 77260 3256
rect 289084 3204 289136 3256
rect 292580 3204 292632 3256
rect 349252 3136 349304 3188
rect 351920 3136 351972 3188
rect 299664 3068 299716 3120
rect 302240 3068 302292 3120
rect 11152 3000 11204 3052
rect 15844 3000 15896 3052
rect 118792 3000 118844 3052
rect 119804 3000 119856 3052
rect 309784 3000 309836 3052
rect 315028 3000 315080 3052
rect 348056 3000 348108 3052
rect 353300 3000 353352 3052
rect 581000 3000 581052 3052
rect 582564 3000 582616 3052
rect 246304 2932 246356 2984
rect 247592 2932 247644 2984
rect 282184 2932 282236 2984
rect 283104 2932 283156 2984
rect 299480 2184 299532 2236
rect 300768 2184 300820 2236
rect 51356 2116 51408 2168
rect 79324 2116 79376 2168
rect 7656 2048 7708 2100
rect 65432 2048 65484 2100
rect 140044 2048 140096 2100
rect 160744 2048 160796 2100
rect 226984 2048 227036 2100
rect 280712 2048 280764 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702914 8156 703520
rect 8116 702908 8168 702914
rect 8116 702850 8168 702856
rect 24320 702846 24348 703520
rect 24308 702840 24360 702846
rect 24308 702782 24360 702788
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 11704 683188 11756 683194
rect 11704 683130 11756 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3148 580984 3200 580990
rect 3148 580926 3200 580932
rect 3160 580009 3188 580926
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3436 576842 3464 632023
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618662 3556 619103
rect 3516 618656 3568 618662
rect 3516 618598 3568 618604
rect 7564 618656 7616 618662
rect 7564 618598 7616 618604
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 576836 3476 576842
rect 3424 576778 3476 576784
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 2778 553888 2834 553897
rect 2778 553823 2780 553832
rect 2832 553823 2834 553832
rect 2780 553794 2832 553800
rect 3436 540258 3464 566879
rect 4804 553852 4856 553858
rect 4804 553794 4856 553800
rect 3424 540252 3476 540258
rect 3424 540194 3476 540200
rect 4816 538218 4844 553794
rect 4804 538212 4856 538218
rect 4804 538154 4856 538160
rect 7576 536790 7604 618598
rect 11716 543726 11744 683130
rect 14464 670744 14516 670750
rect 14464 670686 14516 670692
rect 11704 543720 11756 543726
rect 11704 543662 11756 543668
rect 14476 541686 14504 670686
rect 40052 587178 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 69664 702772 69716 702778
rect 69664 702714 69716 702720
rect 67640 702568 67692 702574
rect 67640 702510 67692 702516
rect 67548 588600 67600 588606
rect 67548 588542 67600 588548
rect 40040 587172 40092 587178
rect 40040 587114 40092 587120
rect 52368 585200 52420 585206
rect 52368 585142 52420 585148
rect 41326 582584 41382 582593
rect 41326 582519 41382 582528
rect 14464 541680 14516 541686
rect 14464 541622 14516 541628
rect 11704 538280 11756 538286
rect 11704 538222 11756 538228
rect 7564 536784 7616 536790
rect 7564 536726 7616 536732
rect 3516 530596 3568 530602
rect 3516 530538 3568 530544
rect 3528 527921 3556 530538
rect 3514 527912 3570 527921
rect 3514 527847 3570 527856
rect 3424 526448 3476 526454
rect 3424 526390 3476 526396
rect 3436 501809 3464 526390
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 11716 476134 11744 538222
rect 21364 514820 21416 514826
rect 21364 514762 21416 514768
rect 8208 476128 8260 476134
rect 8208 476070 8260 476076
rect 11704 476128 11756 476134
rect 11704 476070 11756 476076
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 475250 3464 475623
rect 8220 475250 8248 476070
rect 3424 475244 3476 475250
rect 3424 475186 3476 475192
rect 7564 475244 7616 475250
rect 7564 475186 7616 475192
rect 8208 475244 8260 475250
rect 8208 475186 8260 475192
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3240 449812 3292 449818
rect 3240 449754 3292 449760
rect 3252 449585 3280 449754
rect 3238 449576 3294 449585
rect 3238 449511 3294 449520
rect 3424 443012 3476 443018
rect 3424 442954 3476 442960
rect 3436 423609 3464 442954
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 4804 397520 4856 397526
rect 3422 397488 3478 397497
rect 4804 397462 4856 397468
rect 3422 397423 3478 397432
rect 3436 376718 3464 397423
rect 3516 382288 3568 382294
rect 3516 382230 3568 382236
rect 3424 376712 3476 376718
rect 3424 376654 3476 376660
rect 3528 371385 3556 382230
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 4816 358494 4844 397462
rect 7576 387802 7604 475186
rect 11704 462392 11756 462398
rect 11704 462334 11756 462340
rect 7656 409896 7708 409902
rect 7656 409838 7708 409844
rect 7668 389337 7696 409838
rect 7654 389328 7710 389337
rect 7654 389263 7710 389272
rect 11716 389162 11744 462334
rect 21376 441561 21404 514762
rect 21362 441552 21418 441561
rect 21362 441487 21418 441496
rect 15844 434784 15896 434790
rect 15844 434726 15896 434732
rect 11704 389156 11756 389162
rect 11704 389098 11756 389104
rect 7564 387796 7616 387802
rect 7564 387738 7616 387744
rect 2780 358488 2832 358494
rect 2778 358456 2780 358465
rect 4804 358488 4856 358494
rect 2832 358456 2834 358465
rect 4804 358430 4856 358436
rect 2778 358391 2834 358400
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 11704 345092 11756 345098
rect 11704 345034 11756 345040
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 4080 307834 4108 319223
rect 4068 307828 4120 307834
rect 4068 307770 4120 307776
rect 7564 307828 7616 307834
rect 7564 307770 7616 307776
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 279682 3464 306167
rect 4066 297392 4122 297401
rect 4066 297327 4122 297336
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 3424 279676 3476 279682
rect 3424 279618 3476 279624
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 2780 255196 2832 255202
rect 2780 255138 2832 255144
rect 2792 254153 2820 255138
rect 2778 254144 2834 254153
rect 2778 254079 2834 254088
rect 3424 241120 3476 241126
rect 3422 241088 3424 241097
rect 3476 241088 3478 241097
rect 3422 241023 3478 241032
rect 3424 215008 3476 215014
rect 3422 214976 3424 214985
rect 3476 214976 3478 214985
rect 3422 214911 3478 214920
rect 3240 202156 3292 202162
rect 3240 202098 3292 202104
rect 3252 201929 3280 202098
rect 3238 201920 3294 201929
rect 3238 201855 3294 201864
rect 3424 188896 3476 188902
rect 3422 188864 3424 188873
rect 3476 188864 3478 188873
rect 3422 188799 3478 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3146 149832 3202 149841
rect 3146 149767 3202 149776
rect 3160 145761 3188 149767
rect 3436 147014 3464 162823
rect 3424 147008 3476 147014
rect 3424 146950 3476 146956
rect 3146 145752 3202 145761
rect 3146 145687 3202 145696
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3436 96694 3464 97543
rect 3424 96688 3476 96694
rect 3424 96630 3476 96636
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3148 76560 3200 76566
rect 3148 76502 3200 76508
rect 3160 71641 3188 76502
rect 3146 71632 3202 71641
rect 3146 71567 3202 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3976 50380 4028 50386
rect 3976 50322 4028 50328
rect 3332 46232 3384 46238
rect 3332 46174 3384 46180
rect 3344 45529 3372 46174
rect 3330 45520 3386 45529
rect 3330 45455 3386 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 572 8968 624 8974
rect 572 8910 624 8916
rect 584 480 612 8910
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 3988 3534 4016 50322
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 2884 480 2912 3470
rect 4080 480 4108 297327
rect 4804 280220 4856 280226
rect 4804 280162 4856 280168
rect 4816 255202 4844 280162
rect 7576 279478 7604 307770
rect 9588 306400 9640 306406
rect 9588 306342 9640 306348
rect 7656 279676 7708 279682
rect 7656 279618 7708 279624
rect 7564 279472 7616 279478
rect 7564 279414 7616 279420
rect 7564 261520 7616 261526
rect 7564 261462 7616 261468
rect 4804 255196 4856 255202
rect 4804 255138 4856 255144
rect 5446 221504 5502 221513
rect 5446 221439 5502 221448
rect 5460 6914 5488 221439
rect 7576 215014 7604 261462
rect 7668 253230 7696 279618
rect 7748 262268 7800 262274
rect 7748 262210 7800 262216
rect 7656 253224 7708 253230
rect 7656 253166 7708 253172
rect 7760 241126 7788 262210
rect 7748 241120 7800 241126
rect 7748 241062 7800 241068
rect 7656 231872 7708 231878
rect 7656 231814 7708 231820
rect 7564 215008 7616 215014
rect 7564 214950 7616 214956
rect 6826 203552 6882 203561
rect 6826 203487 6882 203496
rect 6840 6914 6868 203487
rect 7668 188902 7696 231814
rect 8208 215008 8260 215014
rect 8208 214950 8260 214956
rect 7656 188896 7708 188902
rect 7656 188838 7708 188844
rect 8220 114510 8248 214950
rect 8208 114504 8260 114510
rect 8208 114446 8260 114452
rect 7564 106956 7616 106962
rect 7564 106898 7616 106904
rect 5276 6886 5488 6914
rect 6472 6886 6868 6914
rect 5276 480 5304 6886
rect 6472 480 6500 6886
rect 7576 6662 7604 106898
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 9600 3534 9628 306342
rect 11716 288425 11744 345034
rect 13726 332616 13782 332625
rect 13726 332551 13782 332560
rect 11702 288416 11758 288425
rect 11702 288351 11758 288360
rect 12348 180124 12400 180130
rect 12348 180066 12400 180072
rect 10966 156632 11022 156641
rect 10966 156567 11022 156576
rect 10980 3534 11008 156567
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7668 480 7696 2042
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 480 11192 2994
rect 12360 480 12388 180066
rect 13740 6914 13768 332551
rect 15856 319462 15884 434726
rect 41340 417489 41368 582519
rect 50988 582412 51040 582418
rect 50988 582354 51040 582360
rect 48136 560312 48188 560318
rect 48136 560254 48188 560260
rect 42800 541680 42852 541686
rect 42800 541622 42852 541628
rect 42812 541006 42840 541622
rect 42800 541000 42852 541006
rect 42800 540942 42852 540948
rect 43996 541000 44048 541006
rect 43996 540942 44048 540948
rect 41326 417480 41382 417489
rect 41326 417415 41382 417424
rect 39948 411324 40000 411330
rect 39948 411266 40000 411272
rect 37188 343664 37240 343670
rect 37188 343606 37240 343612
rect 31666 335472 31722 335481
rect 31666 335407 31722 335416
rect 22006 329896 22062 329905
rect 22006 329831 22062 329840
rect 15844 319456 15896 319462
rect 15844 319398 15896 319404
rect 17866 307864 17922 307873
rect 17866 307799 17922 307808
rect 15844 302252 15896 302258
rect 15844 302194 15896 302200
rect 14464 292596 14516 292602
rect 14464 292538 14516 292544
rect 14476 241369 14504 292538
rect 14462 241360 14518 241369
rect 14462 241295 14518 241304
rect 15106 236600 15162 236609
rect 15106 236535 15162 236544
rect 15120 6914 15148 236535
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 15856 3058 15884 302194
rect 17880 3534 17908 307799
rect 19248 294636 19300 294642
rect 19248 294578 19300 294584
rect 19260 3534 19288 294578
rect 20626 218648 20682 218657
rect 20626 218583 20682 218592
rect 20640 3534 20668 218583
rect 21364 140820 21416 140826
rect 21364 140762 21416 140768
rect 21376 111790 21404 140762
rect 21364 111784 21416 111790
rect 21364 111726 21416 111732
rect 22020 6914 22048 329831
rect 25502 322960 25558 322969
rect 25502 322895 25558 322904
rect 23386 311944 23442 311953
rect 23386 311879 23442 311888
rect 23400 6914 23428 311879
rect 24766 186960 24822 186969
rect 24766 186895 24822 186904
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15948 480 15976 3402
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 19444 480 19472 3470
rect 20628 3324 20680 3330
rect 20628 3266 20680 3272
rect 20640 480 20668 3266
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 186895
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3470
rect 25516 3330 25544 322895
rect 30286 310584 30342 310593
rect 30286 310519 30342 310528
rect 26146 299568 26202 299577
rect 26146 299503 26202 299512
rect 26160 3534 26188 299503
rect 28906 235240 28962 235249
rect 28906 235175 28962 235184
rect 27528 192500 27580 192506
rect 27528 192442 27580 192448
rect 27540 3534 27568 192442
rect 27712 3664 27764 3670
rect 27712 3606 27764 3612
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 25504 3324 25556 3330
rect 25504 3266 25556 3272
rect 26528 480 26556 3470
rect 27724 480 27752 3606
rect 28920 480 28948 235175
rect 30300 6914 30328 310519
rect 31680 6914 31708 335407
rect 35806 334112 35862 334121
rect 35806 334047 35862 334056
rect 34426 331256 34482 331265
rect 34426 331191 34482 331200
rect 32402 312080 32458 312089
rect 32402 312015 32458 312024
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 32416 3670 32444 312015
rect 33784 290488 33836 290494
rect 33784 290430 33836 290436
rect 33796 267714 33824 290430
rect 33784 267708 33836 267714
rect 33784 267650 33836 267656
rect 34334 251832 34390 251841
rect 34334 251767 34390 251776
rect 33046 217288 33102 217297
rect 33046 217223 33102 217232
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 33060 3534 33088 217223
rect 34348 106962 34376 251767
rect 34336 106956 34388 106962
rect 34336 106898 34388 106904
rect 34440 3534 34468 331191
rect 35820 3534 35848 334047
rect 37096 279472 37148 279478
rect 37096 279414 37148 279420
rect 37108 155242 37136 279414
rect 37096 155236 37148 155242
rect 37096 155178 37148 155184
rect 37094 44840 37150 44849
rect 37094 44775 37150 44784
rect 37108 3534 37136 44775
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 36004 480 36032 3470
rect 37200 480 37228 343606
rect 38566 325816 38622 325825
rect 38566 325751 38622 325760
rect 38580 6914 38608 325751
rect 39960 260166 39988 411266
rect 41236 406428 41288 406434
rect 41236 406370 41288 406376
rect 39948 260160 40000 260166
rect 39948 260102 40000 260108
rect 41144 258732 41196 258738
rect 41144 258674 41196 258680
rect 39946 233880 40002 233889
rect 39946 233815 40002 233824
rect 39960 6914 39988 233815
rect 41156 111110 41184 258674
rect 41248 256018 41276 406370
rect 44008 386374 44036 540942
rect 48148 477562 48176 560254
rect 48228 533384 48280 533390
rect 48228 533326 48280 533332
rect 48136 477556 48188 477562
rect 48136 477498 48188 477504
rect 44088 439000 44140 439006
rect 44088 438942 44140 438948
rect 43996 386368 44048 386374
rect 43996 386310 44048 386316
rect 42708 336796 42760 336802
rect 42708 336738 42760 336744
rect 41326 313440 41382 313449
rect 41326 313375 41382 313384
rect 41236 256012 41288 256018
rect 41236 255954 41288 255960
rect 41144 111104 41196 111110
rect 41144 111046 41196 111052
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3534 41368 313375
rect 42720 3534 42748 336738
rect 43442 301336 43498 301345
rect 43442 301271 43498 301280
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 43456 3466 43484 301271
rect 44100 282198 44128 438942
rect 48148 437510 48176 477498
rect 48136 437504 48188 437510
rect 48136 437446 48188 437452
rect 46848 412684 46900 412690
rect 46848 412626 46900 412632
rect 45376 366376 45428 366382
rect 45376 366318 45428 366324
rect 44088 282192 44140 282198
rect 44088 282134 44140 282140
rect 44088 257372 44140 257378
rect 44088 257314 44140 257320
rect 44100 186318 44128 257314
rect 45388 238066 45416 366318
rect 45466 298752 45522 298761
rect 45466 298687 45522 298696
rect 45376 238060 45428 238066
rect 45376 238002 45428 238008
rect 44088 186312 44140 186318
rect 44088 186254 44140 186260
rect 44100 108322 44128 186254
rect 44088 108316 44140 108322
rect 44088 108258 44140 108264
rect 44088 31068 44140 31074
rect 44088 31010 44140 31016
rect 44100 3534 44128 31010
rect 44272 3936 44324 3942
rect 44272 3878 44324 3884
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 44284 480 44312 3878
rect 45480 480 45508 298687
rect 46860 258806 46888 412626
rect 48136 407176 48188 407182
rect 48136 407118 48188 407124
rect 48148 378049 48176 407118
rect 48240 389094 48268 533326
rect 50896 529236 50948 529242
rect 50896 529178 50948 529184
rect 49608 422952 49660 422958
rect 49608 422894 49660 422900
rect 48228 389088 48280 389094
rect 48228 389030 48280 389036
rect 48134 378040 48190 378049
rect 48134 377975 48190 377984
rect 47582 340912 47638 340921
rect 47582 340847 47638 340856
rect 46848 258800 46900 258806
rect 46848 258742 46900 258748
rect 46848 253972 46900 253978
rect 46848 253914 46900 253920
rect 46756 238060 46808 238066
rect 46756 238002 46808 238008
rect 46768 90817 46796 238002
rect 46860 105602 46888 253914
rect 46848 105596 46900 105602
rect 46848 105538 46900 105544
rect 46754 90808 46810 90817
rect 46754 90743 46810 90752
rect 46848 29640 46900 29646
rect 46848 29582 46900 29588
rect 46860 6914 46888 29582
rect 46676 6886 46888 6914
rect 46676 480 46704 6886
rect 47596 3942 47624 340847
rect 48148 255270 48176 377975
rect 48226 339552 48282 339561
rect 48226 339487 48282 339496
rect 48136 255264 48188 255270
rect 48136 255206 48188 255212
rect 48148 253978 48176 255206
rect 48136 253972 48188 253978
rect 48136 253914 48188 253920
rect 48136 155236 48188 155242
rect 48136 155178 48188 155184
rect 48148 154630 48176 155178
rect 48136 154624 48188 154630
rect 48136 154566 48188 154572
rect 48148 128314 48176 154566
rect 48136 128308 48188 128314
rect 48136 128250 48188 128256
rect 48240 6914 48268 339487
rect 49620 266529 49648 422894
rect 50804 411256 50856 411262
rect 50804 411198 50856 411204
rect 50816 379409 50844 411198
rect 50908 396030 50936 529178
rect 51000 442241 51028 582354
rect 52276 563100 52328 563106
rect 52276 563042 52328 563048
rect 52288 445058 52316 563042
rect 52276 445052 52328 445058
rect 52276 444994 52328 445000
rect 50986 442232 51042 442241
rect 50986 442167 51042 442176
rect 50988 437504 51040 437510
rect 50988 437446 51040 437452
rect 50896 396024 50948 396030
rect 50896 395966 50948 395972
rect 50802 379400 50858 379409
rect 50802 379335 50858 379344
rect 49606 266520 49662 266529
rect 49606 266455 49662 266464
rect 49620 215966 49648 266455
rect 50816 258058 50844 379335
rect 51000 284345 51028 437446
rect 52184 436144 52236 436150
rect 52184 436086 52236 436092
rect 51448 389156 51500 389162
rect 51448 389098 51500 389104
rect 51460 388385 51488 389098
rect 51446 388376 51502 388385
rect 51446 388311 51502 388320
rect 52196 311137 52224 436086
rect 52276 421592 52328 421598
rect 52276 421534 52328 421540
rect 52182 311128 52238 311137
rect 52182 311063 52238 311072
rect 52182 285968 52238 285977
rect 52182 285903 52238 285912
rect 50986 284336 51042 284345
rect 50986 284271 51042 284280
rect 50896 260228 50948 260234
rect 50896 260170 50948 260176
rect 50804 258052 50856 258058
rect 50804 257994 50856 258000
rect 50816 257378 50844 257994
rect 50804 257372 50856 257378
rect 50804 257314 50856 257320
rect 49608 215960 49660 215966
rect 49608 215902 49660 215908
rect 49608 195288 49660 195294
rect 49608 195230 49660 195236
rect 47872 6886 48268 6914
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 47872 480 47900 6886
rect 49620 3534 49648 195230
rect 50908 109070 50936 260170
rect 51000 132462 51028 284271
rect 52196 138689 52224 285903
rect 52288 265062 52316 421534
rect 52380 389162 52408 585142
rect 62028 581120 62080 581126
rect 62028 581062 62080 581068
rect 60648 581052 60700 581058
rect 60648 580994 60700 581000
rect 53656 571396 53708 571402
rect 53656 571338 53708 571344
rect 53668 447914 53696 571338
rect 55036 570648 55088 570654
rect 55036 570590 55088 570596
rect 53748 549296 53800 549302
rect 53748 549238 53800 549244
rect 53656 447908 53708 447914
rect 53656 447850 53708 447856
rect 53656 414044 53708 414050
rect 53656 413986 53708 413992
rect 53380 396772 53432 396778
rect 53380 396714 53432 396720
rect 52368 389156 52420 389162
rect 52368 389098 52420 389104
rect 52366 311128 52422 311137
rect 52366 311063 52422 311072
rect 52380 277370 52408 311063
rect 52368 277364 52420 277370
rect 52368 277306 52420 277312
rect 53288 269136 53340 269142
rect 53288 269078 53340 269084
rect 52276 265056 52328 265062
rect 52276 264998 52328 265004
rect 52368 261588 52420 261594
rect 52368 261530 52420 261536
rect 52276 199436 52328 199442
rect 52276 199378 52328 199384
rect 52182 138680 52238 138689
rect 52182 138615 52238 138624
rect 51722 136776 51778 136785
rect 51722 136711 51778 136720
rect 50988 132456 51040 132462
rect 50988 132398 51040 132404
rect 50896 109064 50948 109070
rect 50896 109006 50948 109012
rect 51736 59362 51764 136711
rect 52288 88330 52316 199378
rect 52380 112470 52408 261530
rect 53300 139505 53328 269078
rect 53392 248470 53420 396714
rect 53564 284504 53616 284510
rect 53564 284446 53616 284452
rect 53472 256012 53524 256018
rect 53472 255954 53524 255960
rect 53380 248464 53432 248470
rect 53380 248406 53432 248412
rect 53484 198626 53512 255954
rect 53472 198620 53524 198626
rect 53472 198562 53524 198568
rect 53286 139496 53342 139505
rect 53286 139431 53342 139440
rect 52368 112464 52420 112470
rect 52368 112406 52420 112412
rect 53484 104854 53512 198562
rect 53576 142866 53604 284446
rect 53668 264246 53696 413986
rect 53760 389230 53788 549238
rect 54944 423700 54996 423706
rect 54944 423642 54996 423648
rect 53840 407108 53892 407114
rect 53840 407050 53892 407056
rect 53852 406434 53880 407050
rect 53840 406428 53892 406434
rect 53840 406370 53892 406376
rect 53748 389224 53800 389230
rect 53748 389166 53800 389172
rect 54758 270736 54814 270745
rect 54758 270671 54814 270680
rect 53656 264240 53708 264246
rect 53656 264182 53708 264188
rect 54772 171134 54800 270671
rect 54956 267782 54984 423642
rect 55048 407114 55076 570590
rect 59268 570036 59320 570042
rect 59268 569978 59320 569984
rect 57704 565888 57756 565894
rect 57704 565830 57756 565836
rect 56508 564460 56560 564466
rect 56508 564402 56560 564408
rect 55128 546508 55180 546514
rect 55128 546450 55180 546456
rect 55036 407108 55088 407114
rect 55036 407050 55088 407056
rect 55036 403028 55088 403034
rect 55036 402970 55088 402976
rect 54944 267776 54996 267782
rect 54944 267718 54996 267724
rect 54864 265062 54892 265093
rect 54852 265056 54904 265062
rect 54850 265024 54852 265033
rect 54904 265024 54906 265033
rect 54850 264959 54906 264968
rect 54864 201482 54892 264959
rect 55048 251870 55076 402970
rect 55140 382129 55168 546450
rect 56416 392012 56468 392018
rect 56416 391954 56468 391960
rect 55126 382120 55182 382129
rect 55126 382055 55182 382064
rect 56428 359514 56456 391954
rect 56520 385014 56548 564402
rect 57612 434104 57664 434110
rect 57612 434046 57664 434052
rect 56508 385008 56560 385014
rect 56508 384950 56560 384956
rect 56416 359508 56468 359514
rect 56416 359450 56468 359456
rect 56428 354674 56456 359450
rect 56428 354646 56548 354674
rect 56416 282940 56468 282946
rect 56416 282882 56468 282888
rect 55036 251864 55088 251870
rect 55036 251806 55088 251812
rect 55126 226944 55182 226953
rect 55126 226879 55182 226888
rect 54852 201476 54904 201482
rect 54852 201418 54904 201424
rect 55036 201476 55088 201482
rect 55036 201418 55088 201424
rect 54772 171106 54984 171134
rect 54956 160721 54984 171106
rect 54942 160712 54998 160721
rect 54942 160647 54998 160656
rect 53748 148368 53800 148374
rect 53748 148310 53800 148316
rect 53564 142860 53616 142866
rect 53564 142802 53616 142808
rect 53654 139496 53710 139505
rect 53654 139431 53710 139440
rect 53668 120086 53696 139431
rect 53656 120080 53708 120086
rect 53656 120022 53708 120028
rect 53472 104848 53524 104854
rect 53472 104790 53524 104796
rect 52276 88324 52328 88330
rect 52276 88266 52328 88272
rect 51724 59356 51776 59362
rect 51724 59298 51776 59304
rect 50988 18624 51040 18630
rect 50988 18566 51040 18572
rect 51000 3534 51028 18566
rect 52552 6180 52604 6186
rect 52552 6122 52604 6128
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51356 2168 51408 2174
rect 51356 2110 51408 2116
rect 51368 480 51396 2110
rect 52564 480 52592 6122
rect 53760 480 53788 148310
rect 54484 135992 54536 135998
rect 54484 135934 54536 135940
rect 54496 33114 54524 135934
rect 54956 121446 54984 160647
rect 55048 149122 55076 201418
rect 55036 149116 55088 149122
rect 55036 149058 55088 149064
rect 54944 121440 54996 121446
rect 54944 121382 54996 121388
rect 55048 115938 55076 149058
rect 55036 115932 55088 115938
rect 55036 115874 55088 115880
rect 55140 101454 55168 226879
rect 56428 171834 56456 282882
rect 56520 244254 56548 354646
rect 57624 310486 57652 434046
rect 57716 411262 57744 565830
rect 57888 558952 57940 558958
rect 57888 558894 57940 558900
rect 57796 425740 57848 425746
rect 57796 425682 57848 425688
rect 57704 411256 57756 411262
rect 57704 411198 57756 411204
rect 57612 310480 57664 310486
rect 57612 310422 57664 310428
rect 57520 309936 57572 309942
rect 57520 309878 57572 309884
rect 57244 270496 57296 270502
rect 57244 270438 57296 270444
rect 57256 269142 57284 270438
rect 57244 269136 57296 269142
rect 57244 269078 57296 269084
rect 56508 244248 56560 244254
rect 56508 244190 56560 244196
rect 56506 239456 56562 239465
rect 56506 239391 56562 239400
rect 56520 211138 56548 239391
rect 57532 238377 57560 309878
rect 57704 275324 57756 275330
rect 57704 275266 57756 275272
rect 57518 238368 57574 238377
rect 57518 238303 57574 238312
rect 56508 211132 56560 211138
rect 56508 211074 56560 211080
rect 56416 171828 56468 171834
rect 56416 171770 56468 171776
rect 56428 133210 56456 171770
rect 56416 133204 56468 133210
rect 56416 133146 56468 133152
rect 55128 101448 55180 101454
rect 55128 101390 55180 101396
rect 56520 92478 56548 211074
rect 57716 142390 57744 275266
rect 57808 270502 57836 425682
rect 57900 399537 57928 558894
rect 59176 545148 59228 545154
rect 59176 545090 59228 545096
rect 59084 518220 59136 518226
rect 59084 518162 59136 518168
rect 58898 430672 58954 430681
rect 58898 430607 58954 430616
rect 57886 399528 57942 399537
rect 57886 399463 57942 399472
rect 57888 310480 57940 310486
rect 57888 310422 57940 310428
rect 57900 309806 57928 310422
rect 57888 309800 57940 309806
rect 57888 309742 57940 309748
rect 57900 276010 57928 309742
rect 57888 276004 57940 276010
rect 57888 275946 57940 275952
rect 58912 273358 58940 430607
rect 59096 408474 59124 518162
rect 59188 476066 59216 545090
rect 59176 476060 59228 476066
rect 59176 476002 59228 476008
rect 59280 449954 59308 569978
rect 60464 452668 60516 452674
rect 60464 452610 60516 452616
rect 59268 449948 59320 449954
rect 59268 449890 59320 449896
rect 59176 445868 59228 445874
rect 59176 445810 59228 445816
rect 59188 418334 59216 445810
rect 59280 418810 59308 449890
rect 60476 420918 60504 452610
rect 60556 445052 60608 445058
rect 60556 444994 60608 445000
rect 60568 444446 60596 444994
rect 60556 444440 60608 444446
rect 60556 444382 60608 444388
rect 60464 420912 60516 420918
rect 60464 420854 60516 420860
rect 59268 418804 59320 418810
rect 59268 418746 59320 418752
rect 59176 418328 59228 418334
rect 59176 418270 59228 418276
rect 59084 408468 59136 408474
rect 59084 408410 59136 408416
rect 59082 385656 59138 385665
rect 59082 385591 59138 385600
rect 58992 293276 59044 293282
rect 58992 293218 59044 293224
rect 58900 273352 58952 273358
rect 58900 273294 58952 273300
rect 57796 270496 57848 270502
rect 57796 270438 57848 270444
rect 57796 267776 57848 267782
rect 57796 267718 57848 267724
rect 57808 146946 57836 267718
rect 57888 248464 57940 248470
rect 57888 248406 57940 248412
rect 57796 146940 57848 146946
rect 57796 146882 57848 146888
rect 57704 142384 57756 142390
rect 57704 142326 57756 142332
rect 57610 138816 57666 138825
rect 57610 138751 57666 138760
rect 57624 126954 57652 138751
rect 57612 126948 57664 126954
rect 57612 126890 57664 126896
rect 57716 124166 57744 142326
rect 57704 124160 57756 124166
rect 57704 124102 57756 124108
rect 57808 118658 57836 146882
rect 57796 118652 57848 118658
rect 57796 118594 57848 118600
rect 57152 111104 57204 111110
rect 57152 111046 57204 111052
rect 57164 110498 57192 111046
rect 57152 110492 57204 110498
rect 57152 110434 57204 110440
rect 57796 110492 57848 110498
rect 57796 110434 57848 110440
rect 57244 109064 57296 109070
rect 57244 109006 57296 109012
rect 56508 92472 56560 92478
rect 56508 92414 56560 92420
rect 57256 85542 57284 109006
rect 57244 85536 57296 85542
rect 57244 85478 57296 85484
rect 57808 75886 57836 110434
rect 57900 100026 57928 248406
rect 58900 244316 58952 244322
rect 58900 244258 58952 244264
rect 58912 211818 58940 244258
rect 59004 241534 59032 293218
rect 58992 241528 59044 241534
rect 58992 241470 59044 241476
rect 59096 237386 59124 385591
rect 59188 263702 59216 418270
rect 60568 380254 60596 444382
rect 60660 434110 60688 580994
rect 61936 557592 61988 557598
rect 61936 557534 61988 557540
rect 61842 534712 61898 534721
rect 61842 534647 61898 534656
rect 60648 434104 60700 434110
rect 60648 434046 60700 434052
rect 61658 429312 61714 429321
rect 61658 429247 61714 429256
rect 60648 400240 60700 400246
rect 60648 400182 60700 400188
rect 60556 380248 60608 380254
rect 60556 380190 60608 380196
rect 60464 304292 60516 304298
rect 60464 304234 60516 304240
rect 60476 279478 60504 304234
rect 60660 287054 60688 400182
rect 60568 287026 60688 287054
rect 60568 283393 60596 287026
rect 60554 283384 60610 283393
rect 60554 283319 60610 283328
rect 60464 279472 60516 279478
rect 60464 279414 60516 279420
rect 59176 263696 59228 263702
rect 59176 263638 59228 263644
rect 59084 237380 59136 237386
rect 59084 237322 59136 237328
rect 58900 211812 58952 211818
rect 58900 211754 58952 211760
rect 58912 209774 58940 211754
rect 58912 209746 59124 209774
rect 57888 100020 57940 100026
rect 57888 99962 57940 99968
rect 59096 95946 59124 209746
rect 59188 143721 59216 263638
rect 60464 260160 60516 260166
rect 60464 260102 60516 260108
rect 60476 258233 60504 260102
rect 60462 258224 60518 258233
rect 60462 258159 60518 258168
rect 60004 256012 60056 256018
rect 60004 255954 60056 255960
rect 60016 254590 60044 255954
rect 60004 254584 60056 254590
rect 60004 254526 60056 254532
rect 59268 241596 59320 241602
rect 59268 241538 59320 241544
rect 59174 143712 59230 143721
rect 59174 143647 59230 143656
rect 59188 114510 59216 143647
rect 59176 114504 59228 114510
rect 59176 114446 59228 114452
rect 59084 95940 59136 95946
rect 59084 95882 59136 95888
rect 59280 92614 59308 241538
rect 60476 233209 60504 258159
rect 60568 250782 60596 283319
rect 60648 273352 60700 273358
rect 60648 273294 60700 273300
rect 60556 250776 60608 250782
rect 60556 250718 60608 250724
rect 60556 247104 60608 247110
rect 60556 247046 60608 247052
rect 60462 233200 60518 233209
rect 60462 233135 60518 233144
rect 60568 187746 60596 247046
rect 60556 187740 60608 187746
rect 60556 187682 60608 187688
rect 60464 164212 60516 164218
rect 60464 164154 60516 164160
rect 60476 163538 60504 164154
rect 60464 163532 60516 163538
rect 60464 163474 60516 163480
rect 60476 124846 60504 163474
rect 60464 124840 60516 124846
rect 60464 124782 60516 124788
rect 60568 99346 60596 187682
rect 60660 164218 60688 273294
rect 61672 271998 61700 429247
rect 61750 414352 61806 414361
rect 61750 414287 61806 414296
rect 61764 290465 61792 414287
rect 61856 393446 61884 534647
rect 61948 522306 61976 557534
rect 61936 522300 61988 522306
rect 61936 522242 61988 522248
rect 62040 460970 62068 581062
rect 65982 580000 66038 580009
rect 65982 579935 66038 579944
rect 64696 568608 64748 568614
rect 64696 568550 64748 568556
rect 63316 553444 63368 553450
rect 63316 553386 63368 553392
rect 62028 460964 62080 460970
rect 62028 460906 62080 460912
rect 61934 436248 61990 436257
rect 61934 436183 61990 436192
rect 61844 393440 61896 393446
rect 61844 393382 61896 393388
rect 61750 290456 61806 290465
rect 61750 290391 61806 290400
rect 61660 271992 61712 271998
rect 61660 271934 61712 271940
rect 61764 261594 61792 290391
rect 61844 289128 61896 289134
rect 61844 289070 61896 289076
rect 61016 261588 61068 261594
rect 61016 261530 61068 261536
rect 61752 261588 61804 261594
rect 61752 261530 61804 261536
rect 61028 260953 61056 261530
rect 61014 260944 61070 260953
rect 61014 260879 61070 260888
rect 61752 242956 61804 242962
rect 61752 242898 61804 242904
rect 61764 209774 61792 242898
rect 61856 233918 61884 289070
rect 61948 287026 61976 436183
rect 62040 422278 62068 460906
rect 63224 441652 63276 441658
rect 63224 441594 63276 441600
rect 62028 422272 62080 422278
rect 62028 422214 62080 422220
rect 62040 421598 62068 422214
rect 62028 421592 62080 421598
rect 62028 421534 62080 421540
rect 63236 415070 63264 441594
rect 63328 416770 63356 553386
rect 64708 527882 64736 568550
rect 65890 567624 65946 567633
rect 65890 567559 65946 567568
rect 65904 538801 65932 567559
rect 65890 538792 65946 538801
rect 65890 538727 65946 538736
rect 64788 532024 64840 532030
rect 64788 531966 64840 531972
rect 64696 527876 64748 527882
rect 64696 527818 64748 527824
rect 64800 462398 64828 531966
rect 65996 490618 66024 579935
rect 67178 578640 67234 578649
rect 67178 578575 67234 578584
rect 66718 573200 66774 573209
rect 66718 573135 66774 573144
rect 66732 570654 66760 573135
rect 66810 571840 66866 571849
rect 66810 571775 66866 571784
rect 66824 571402 66852 571775
rect 66812 571396 66864 571402
rect 66812 571338 66864 571344
rect 66720 570648 66772 570654
rect 66720 570590 66772 570596
rect 66902 570208 66958 570217
rect 66902 570143 66958 570152
rect 66916 570042 66944 570143
rect 66904 570036 66956 570042
rect 66904 569978 66956 569984
rect 66534 568984 66590 568993
rect 66534 568919 66590 568928
rect 66548 568614 66576 568919
rect 66536 568608 66588 568614
rect 66536 568550 66588 568556
rect 66902 564768 66958 564777
rect 66902 564703 66958 564712
rect 66916 564466 66944 564703
rect 66904 564460 66956 564466
rect 66904 564402 66956 564408
rect 66902 563408 66958 563417
rect 66902 563343 66958 563352
rect 66916 563106 66944 563343
rect 66904 563100 66956 563106
rect 66904 563042 66956 563048
rect 66166 562048 66222 562057
rect 66166 561983 66222 561992
rect 66074 544096 66130 544105
rect 66074 544031 66130 544040
rect 65984 490612 66036 490618
rect 65984 490554 66036 490560
rect 64788 462392 64840 462398
rect 64788 462334 64840 462340
rect 64696 448588 64748 448594
rect 64696 448530 64748 448536
rect 64604 431996 64656 432002
rect 64604 431938 64656 431944
rect 63408 426488 63460 426494
rect 63408 426430 63460 426436
rect 63316 416764 63368 416770
rect 63316 416706 63368 416712
rect 63224 415064 63276 415070
rect 63224 415006 63276 415012
rect 62764 408536 62816 408542
rect 62764 408478 62816 408484
rect 62776 292574 62804 408478
rect 63316 397520 63368 397526
rect 63316 397462 63368 397468
rect 63328 365702 63356 397462
rect 63316 365696 63368 365702
rect 63316 365638 63368 365644
rect 62776 292546 63172 292574
rect 63144 289105 63172 292546
rect 63130 289096 63186 289105
rect 63130 289031 63186 289040
rect 61936 287020 61988 287026
rect 61936 286962 61988 286968
rect 61936 271992 61988 271998
rect 61936 271934 61988 271940
rect 61844 233912 61896 233918
rect 61844 233854 61896 233860
rect 61764 209746 61884 209774
rect 61856 196625 61884 209746
rect 61842 196616 61898 196625
rect 61842 196551 61898 196560
rect 60648 164212 60700 164218
rect 60648 164154 60700 164160
rect 61660 153876 61712 153882
rect 61660 153818 61712 153824
rect 60648 152584 60700 152590
rect 60648 152526 60700 152532
rect 60556 99340 60608 99346
rect 60556 99282 60608 99288
rect 59268 92608 59320 92614
rect 59268 92550 59320 92556
rect 60660 92410 60688 152526
rect 60740 106956 60792 106962
rect 60740 106898 60792 106904
rect 60752 106350 60780 106898
rect 60740 106344 60792 106350
rect 60740 106286 60792 106292
rect 61384 96688 61436 96694
rect 61384 96630 61436 96636
rect 60648 92404 60700 92410
rect 60648 92346 60700 92352
rect 61396 79937 61424 96630
rect 61672 89622 61700 153818
rect 61752 150476 61804 150482
rect 61752 150418 61804 150424
rect 61764 117230 61792 150418
rect 61752 117224 61804 117230
rect 61752 117166 61804 117172
rect 61856 95198 61884 196551
rect 61948 157418 61976 271934
rect 62028 266416 62080 266422
rect 62028 266358 62080 266364
rect 61936 157412 61988 157418
rect 61936 157354 61988 157360
rect 61948 121378 61976 157354
rect 62040 150482 62068 266358
rect 63144 255474 63172 289031
rect 63224 283008 63276 283014
rect 63224 282950 63276 282956
rect 63132 255468 63184 255474
rect 63132 255410 63184 255416
rect 63038 252784 63094 252793
rect 63038 252719 63094 252728
rect 63052 151814 63080 252719
rect 63236 231130 63264 282950
rect 63316 276072 63368 276078
rect 63316 276014 63368 276020
rect 63224 231124 63276 231130
rect 63224 231066 63276 231072
rect 63328 165646 63356 276014
rect 63420 270638 63448 426430
rect 64616 401674 64644 431938
rect 64708 418130 64736 448530
rect 64800 422958 64828 462334
rect 65984 443556 66036 443562
rect 65984 443498 66036 443504
rect 65996 438190 66024 443498
rect 66088 439657 66116 544031
rect 66074 439648 66130 439657
rect 66074 439583 66130 439592
rect 65984 438184 66036 438190
rect 65984 438126 66036 438132
rect 65996 425241 66024 438126
rect 66074 430400 66130 430409
rect 66074 430335 66130 430344
rect 65982 425232 66038 425241
rect 65982 425167 66038 425176
rect 64788 422952 64840 422958
rect 64788 422894 64840 422900
rect 64788 420300 64840 420306
rect 64788 420242 64840 420248
rect 64696 418124 64748 418130
rect 64696 418066 64748 418072
rect 64696 404388 64748 404394
rect 64696 404330 64748 404336
rect 64604 401668 64656 401674
rect 64604 401610 64656 401616
rect 63500 282192 63552 282198
rect 63500 282134 63552 282140
rect 63512 281654 63540 282134
rect 63500 281648 63552 281654
rect 63500 281590 63552 281596
rect 64604 281648 64656 281654
rect 64604 281590 64656 281596
rect 64616 278730 64644 281590
rect 64604 278724 64656 278730
rect 64604 278666 64656 278672
rect 63408 270632 63460 270638
rect 63408 270574 63460 270580
rect 64604 270632 64656 270638
rect 64604 270574 64656 270580
rect 64512 258800 64564 258806
rect 64512 258742 64564 258748
rect 64524 235278 64552 258742
rect 64512 235272 64564 235278
rect 64512 235214 64564 235220
rect 64616 171134 64644 270574
rect 64708 252793 64736 404330
rect 64800 266422 64828 420242
rect 65890 399528 65946 399537
rect 65890 399463 65946 399472
rect 65904 398857 65932 399463
rect 65890 398848 65946 398857
rect 65890 398783 65946 398792
rect 65904 373969 65932 398783
rect 65890 373960 65946 373969
rect 65890 373895 65946 373904
rect 65800 291848 65852 291854
rect 65800 291790 65852 291796
rect 65706 273184 65762 273193
rect 65706 273119 65762 273128
rect 64788 266416 64840 266422
rect 64788 266358 64840 266364
rect 64788 264988 64840 264994
rect 64788 264930 64840 264936
rect 64694 252784 64750 252793
rect 64694 252719 64750 252728
rect 64616 171106 64736 171134
rect 63316 165640 63368 165646
rect 63316 165582 63368 165588
rect 63052 151786 63264 151814
rect 62028 150476 62080 150482
rect 62028 150418 62080 150424
rect 63132 143608 63184 143614
rect 63132 143550 63184 143556
rect 61936 121372 61988 121378
rect 61936 121314 61988 121320
rect 63144 114442 63172 143550
rect 63236 139641 63264 151786
rect 63222 139632 63278 139641
rect 63222 139567 63278 139576
rect 63132 114436 63184 114442
rect 63132 114378 63184 114384
rect 61936 106344 61988 106350
rect 61936 106286 61988 106292
rect 61844 95192 61896 95198
rect 61844 95134 61896 95140
rect 61660 89616 61712 89622
rect 61660 89558 61712 89564
rect 61382 79928 61438 79937
rect 61382 79863 61438 79872
rect 57796 75880 57848 75886
rect 57796 75822 57848 75828
rect 57888 73840 57940 73846
rect 57888 73782 57940 73788
rect 55128 33788 55180 33794
rect 55128 33730 55180 33736
rect 54484 33108 54536 33114
rect 54484 33050 54536 33056
rect 55140 6914 55168 33730
rect 56508 25560 56560 25566
rect 56508 25502 56560 25508
rect 54956 6886 55168 6914
rect 54956 480 54984 6886
rect 56520 3534 56548 25502
rect 57900 3534 57928 73782
rect 61948 71738 61976 106286
rect 63236 103494 63264 139567
rect 63328 126886 63356 165582
rect 64708 158778 64736 171106
rect 64696 158772 64748 158778
rect 64696 158714 64748 158720
rect 64604 152516 64656 152522
rect 64604 152458 64656 152464
rect 64510 151056 64566 151065
rect 64510 150991 64566 151000
rect 63408 141432 63460 141438
rect 63408 141374 63460 141380
rect 63316 126880 63368 126886
rect 63316 126822 63368 126828
rect 63224 103488 63276 103494
rect 63224 103430 63276 103436
rect 63420 91050 63448 141374
rect 64524 117298 64552 150991
rect 64512 117292 64564 117298
rect 64512 117234 64564 117240
rect 64616 115326 64644 152458
rect 64708 120018 64736 158714
rect 64800 152522 64828 264930
rect 65720 171134 65748 273119
rect 65812 260234 65840 291790
rect 65996 287609 66024 425167
rect 65982 287600 66038 287609
rect 65982 287535 66038 287544
rect 65984 287020 66036 287026
rect 65984 286962 66036 286968
rect 65996 286249 66024 286962
rect 65982 286240 66038 286249
rect 65982 286175 66038 286184
rect 65892 262268 65944 262274
rect 65892 262210 65944 262216
rect 65800 260228 65852 260234
rect 65800 260170 65852 260176
rect 65904 228410 65932 262210
rect 65996 240106 66024 286175
rect 66088 273193 66116 430335
rect 66180 384946 66208 561983
rect 66810 560688 66866 560697
rect 66810 560623 66866 560632
rect 66824 560318 66852 560623
rect 66812 560312 66864 560318
rect 66812 560254 66864 560260
rect 66810 559328 66866 559337
rect 66810 559263 66866 559272
rect 66824 558958 66852 559263
rect 66812 558952 66864 558958
rect 66812 558894 66864 558900
rect 66810 557968 66866 557977
rect 66810 557903 66866 557912
rect 66824 557598 66852 557903
rect 66812 557592 66864 557598
rect 66812 557534 66864 557540
rect 66902 553616 66958 553625
rect 66902 553551 66958 553560
rect 66916 553450 66944 553551
rect 66904 553444 66956 553450
rect 66904 553386 66956 553392
rect 66718 549536 66774 549545
rect 66718 549471 66774 549480
rect 66732 549302 66760 549471
rect 66720 549296 66772 549302
rect 66720 549238 66772 549244
rect 66810 546816 66866 546825
rect 66810 546751 66866 546760
rect 66824 546514 66852 546751
rect 66812 546508 66864 546514
rect 66812 546450 66864 546456
rect 66810 545456 66866 545465
rect 66810 545391 66866 545400
rect 66824 545154 66852 545391
rect 66812 545148 66864 545154
rect 66812 545090 66864 545096
rect 66626 541376 66682 541385
rect 66626 541311 66682 541320
rect 66640 541006 66668 541311
rect 66628 541000 66680 541006
rect 66628 540942 66680 540948
rect 67088 440904 67140 440910
rect 67088 440846 67140 440852
rect 66812 434104 66864 434110
rect 66812 434046 66864 434052
rect 66824 433401 66852 434046
rect 66810 433392 66866 433401
rect 66810 433327 66866 433336
rect 67100 428233 67128 440846
rect 67086 428224 67142 428233
rect 67086 428159 67142 428168
rect 66994 427408 67050 427417
rect 66994 427343 67050 427352
rect 67008 426494 67036 427343
rect 66996 426488 67048 426494
rect 66996 426430 67048 426436
rect 66626 424144 66682 424153
rect 66626 424079 66682 424088
rect 66640 423706 66668 424079
rect 66628 423700 66680 423706
rect 66628 423642 66680 423648
rect 66810 423328 66866 423337
rect 66810 423263 66866 423272
rect 66824 422958 66852 423263
rect 66812 422952 66864 422958
rect 66812 422894 66864 422900
rect 66628 422272 66680 422278
rect 66628 422214 66680 422220
rect 67086 422240 67142 422249
rect 66640 421161 66668 422214
rect 67086 422175 67142 422184
rect 66626 421152 66682 421161
rect 66626 421087 66682 421096
rect 66812 420912 66864 420918
rect 66812 420854 66864 420860
rect 66824 420073 66852 420854
rect 67100 420306 67128 422175
rect 67088 420300 67140 420306
rect 67088 420242 67140 420248
rect 66810 420064 66866 420073
rect 66810 419999 66866 420008
rect 66810 418976 66866 418985
rect 66810 418911 66866 418920
rect 66824 418334 66852 418911
rect 66812 418328 66864 418334
rect 66812 418270 66864 418276
rect 67086 418160 67142 418169
rect 67086 418095 67088 418104
rect 67140 418095 67142 418104
rect 67088 418066 67140 418072
rect 66260 416764 66312 416770
rect 66260 416706 66312 416712
rect 66272 415993 66300 416706
rect 66258 415984 66314 415993
rect 66258 415919 66314 415928
rect 66272 414361 66300 415919
rect 66904 415064 66956 415070
rect 66904 415006 66956 415012
rect 66810 414896 66866 414905
rect 66810 414831 66866 414840
rect 66258 414352 66314 414361
rect 66258 414287 66314 414296
rect 66824 414050 66852 414831
rect 66916 414089 66944 415006
rect 66902 414080 66958 414089
rect 66812 414044 66864 414050
rect 66902 414015 66958 414024
rect 66812 413986 66864 413992
rect 66258 412992 66314 413001
rect 66258 412927 66314 412936
rect 66272 412690 66300 412927
rect 66260 412684 66312 412690
rect 66260 412626 66312 412632
rect 66258 411904 66314 411913
rect 66258 411839 66314 411848
rect 66272 411330 66300 411839
rect 66260 411324 66312 411330
rect 66260 411266 66312 411272
rect 66628 411256 66680 411262
rect 66628 411198 66680 411204
rect 66640 410825 66668 411198
rect 66626 410816 66682 410825
rect 66626 410751 66682 410760
rect 66810 408912 66866 408921
rect 66810 408847 66866 408856
rect 66824 408542 66852 408847
rect 66812 408536 66864 408542
rect 66812 408478 66864 408484
rect 66902 407824 66958 407833
rect 66902 407759 66958 407768
rect 66916 407182 66944 407759
rect 66904 407176 66956 407182
rect 66904 407118 66956 407124
rect 66812 407108 66864 407114
rect 66812 407050 66864 407056
rect 66824 406745 66852 407050
rect 66810 406736 66866 406745
rect 66810 406671 66866 406680
rect 66810 404560 66866 404569
rect 66810 404495 66866 404504
rect 66824 404394 66852 404495
rect 66812 404388 66864 404394
rect 66812 404330 66864 404336
rect 66810 403744 66866 403753
rect 66810 403679 66866 403688
rect 66824 403034 66852 403679
rect 66812 403028 66864 403034
rect 66812 402970 66864 402976
rect 67192 402665 67220 578575
rect 67454 577280 67510 577289
rect 67454 577215 67510 577224
rect 67362 555248 67418 555257
rect 67362 555183 67418 555192
rect 67270 552256 67326 552265
rect 67270 552191 67326 552200
rect 67284 539102 67312 552191
rect 67272 539096 67324 539102
rect 67272 539038 67324 539044
rect 67376 530670 67404 555183
rect 67364 530664 67416 530670
rect 67364 530606 67416 530612
rect 67468 441614 67496 577215
rect 67560 575385 67588 588542
rect 67546 575376 67602 575385
rect 67546 575311 67602 575320
rect 67652 566681 67680 702510
rect 69676 581074 69704 702714
rect 71688 700324 71740 700330
rect 71688 700266 71740 700272
rect 71700 588606 71728 700266
rect 71792 596329 71820 702986
rect 86224 702840 86276 702846
rect 86224 702782 86276 702788
rect 84108 702636 84160 702642
rect 84108 702578 84160 702584
rect 79968 702500 80020 702506
rect 79968 702442 80020 702448
rect 74540 656940 74592 656946
rect 74540 656882 74592 656888
rect 71778 596320 71834 596329
rect 71778 596255 71834 596264
rect 74552 596174 74580 656882
rect 74552 596146 74672 596174
rect 71688 588600 71740 588606
rect 71688 588542 71740 588548
rect 69940 582412 69992 582418
rect 69940 582354 69992 582360
rect 73528 582412 73580 582418
rect 73528 582354 73580 582360
rect 69032 581058 69704 581074
rect 69020 581052 69704 581058
rect 69072 581046 69704 581052
rect 69952 581074 69980 582354
rect 73540 581074 73568 582354
rect 74262 581224 74318 581233
rect 74262 581159 74318 581168
rect 74276 581074 74304 581159
rect 69952 581046 70288 581074
rect 73232 581046 73568 581074
rect 74152 581046 74304 581074
rect 74644 581074 74672 596146
rect 79980 589898 80008 702442
rect 84120 592686 84148 702578
rect 81440 592680 81492 592686
rect 81440 592622 81492 592628
rect 84108 592680 84160 592686
rect 84108 592622 84160 592628
rect 79324 589892 79376 589898
rect 79324 589834 79376 589840
rect 79968 589892 80020 589898
rect 79968 589834 80020 589840
rect 78128 585812 78180 585818
rect 78128 585754 78180 585760
rect 76288 583772 76340 583778
rect 76288 583714 76340 583720
rect 75366 581088 75422 581097
rect 74644 581046 75366 581074
rect 76300 581074 76328 583714
rect 77208 582820 77260 582826
rect 77208 582762 77260 582768
rect 77220 581074 77248 582762
rect 78140 581074 78168 585754
rect 79336 582826 79364 589834
rect 79980 589354 80008 589834
rect 79968 589348 80020 589354
rect 79968 589290 80020 589296
rect 79324 582820 79376 582826
rect 79324 582762 79376 582768
rect 79048 582480 79100 582486
rect 79048 582422 79100 582428
rect 80702 582448 80758 582457
rect 79060 581074 79088 582422
rect 80702 582383 80758 582392
rect 75992 581046 76328 581074
rect 76912 581046 77248 581074
rect 77832 581046 78168 581074
rect 78752 581046 79088 581074
rect 80244 581052 80296 581058
rect 75366 581023 75422 581032
rect 69020 580994 69072 581000
rect 80244 580994 80296 581000
rect 80256 580938 80284 580994
rect 80716 580938 80744 582383
rect 81452 581346 81480 592622
rect 82728 586560 82780 586566
rect 82728 586502 82780 586508
rect 81452 581318 81526 581346
rect 81498 581060 81526 581318
rect 82740 581074 82768 586502
rect 84292 585200 84344 585206
rect 84292 585142 84344 585148
rect 83002 582584 83058 582593
rect 83002 582519 83058 582528
rect 82432 581046 82768 581074
rect 83016 581074 83044 582519
rect 84304 581074 84332 585142
rect 85486 583944 85542 583953
rect 85486 583879 85542 583888
rect 85500 581074 85528 583879
rect 86236 582554 86264 702782
rect 89180 702434 89208 703520
rect 102048 703044 102100 703050
rect 102048 702986 102100 702992
rect 96620 702908 96672 702914
rect 96620 702850 96672 702856
rect 90364 702704 90416 702710
rect 90364 702646 90416 702652
rect 88352 702406 89208 702434
rect 88352 585818 88380 702406
rect 90376 596174 90404 702646
rect 93124 605872 93176 605878
rect 93124 605814 93176 605820
rect 90376 596146 90588 596174
rect 88340 585812 88392 585818
rect 88340 585754 88392 585760
rect 87512 585200 87564 585206
rect 87512 585142 87564 585148
rect 86224 582548 86276 582554
rect 86224 582490 86276 582496
rect 86236 581346 86264 582490
rect 86868 582480 86920 582486
rect 86868 582422 86920 582428
rect 86236 581318 86310 581346
rect 83016 581046 83352 581074
rect 84304 581046 84456 581074
rect 85376 581046 85528 581074
rect 86282 581060 86310 581318
rect 80256 580910 80744 580938
rect 71502 580816 71558 580825
rect 71208 580774 71502 580802
rect 72422 580816 72478 580825
rect 72128 580774 72422 580802
rect 71502 580751 71558 580760
rect 79874 580816 79930 580825
rect 79672 580774 79874 580802
rect 72422 580751 72478 580760
rect 79874 580751 79930 580760
rect 86880 580718 86908 582422
rect 87524 581074 87552 585142
rect 88246 582584 88302 582593
rect 88246 582519 88302 582528
rect 88260 581074 88288 582519
rect 90560 581126 90588 596146
rect 93136 584458 93164 605814
rect 93124 584452 93176 584458
rect 93124 584394 93176 584400
rect 92110 583808 92166 583817
rect 92110 583743 92166 583752
rect 90548 581120 90600 581126
rect 87216 581046 87552 581074
rect 88136 581046 88288 581074
rect 89976 581058 90312 581074
rect 92124 581074 92152 583743
rect 95884 582412 95936 582418
rect 95884 582354 95936 582360
rect 90600 581068 90896 581074
rect 90548 581062 90896 581068
rect 89976 581052 90324 581058
rect 89976 581046 90272 581052
rect 90560 581046 90896 581062
rect 91816 581046 92152 581074
rect 90272 580994 90324 581000
rect 88706 580816 88762 580825
rect 92386 580816 92442 580825
rect 88762 580774 89056 580802
rect 88706 580751 88762 580760
rect 92442 580774 92736 580802
rect 93656 580774 93808 580802
rect 92386 580751 92442 580760
rect 93780 580718 93808 580774
rect 86868 580712 86920 580718
rect 86868 580654 86920 580660
rect 93768 580712 93820 580718
rect 93768 580654 93820 580660
rect 94576 580366 94728 580394
rect 67732 576836 67784 576842
rect 67732 576778 67784 576784
rect 67744 575929 67772 576778
rect 67730 575920 67786 575929
rect 67730 575855 67786 575864
rect 67638 566672 67694 566681
rect 67638 566607 67694 566616
rect 67652 565894 67680 566607
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67640 543720 67692 543726
rect 67640 543662 67692 543668
rect 67652 463078 67680 543662
rect 67744 479505 67772 575855
rect 94700 573374 94728 580366
rect 95238 574832 95294 574841
rect 95238 574767 95294 574776
rect 94688 573368 94740 573374
rect 94688 573310 94740 573316
rect 94686 563680 94742 563689
rect 94686 563615 94742 563624
rect 67822 556608 67878 556617
rect 67822 556543 67878 556552
rect 67836 534750 67864 556543
rect 68650 548312 68706 548321
rect 68650 548247 68706 548256
rect 68376 543720 68428 543726
rect 68376 543662 68428 543668
rect 68388 543357 68416 543662
rect 68664 543561 68692 548247
rect 68650 543552 68706 543561
rect 68650 543487 68706 543496
rect 68374 543348 68430 543357
rect 68374 543283 68430 543292
rect 69400 539850 69736 539866
rect 69388 539844 69736 539850
rect 69440 539838 69736 539844
rect 91008 539844 91060 539850
rect 69388 539786 69440 539792
rect 91008 539786 91060 539792
rect 68816 539158 68968 539186
rect 68940 536178 68968 539158
rect 68928 536172 68980 536178
rect 68928 536114 68980 536120
rect 67824 534744 67876 534750
rect 67824 534686 67876 534692
rect 69400 528554 69428 539786
rect 70306 539744 70362 539753
rect 70306 539679 70308 539688
rect 70360 539679 70362 539688
rect 76564 539708 76616 539714
rect 70308 539650 70360 539656
rect 76564 539650 76616 539656
rect 70656 539158 70716 539186
rect 70688 538218 70716 539158
rect 70872 539158 71576 539186
rect 71792 539158 72496 539186
rect 73416 539158 73476 539186
rect 70676 538212 70728 538218
rect 70676 538154 70728 538160
rect 70688 536858 70716 538154
rect 70676 536852 70728 536858
rect 70676 536794 70728 536800
rect 70872 528554 70900 539158
rect 71044 536852 71096 536858
rect 71044 536794 71096 536800
rect 69032 528526 69428 528554
rect 70504 528526 70900 528554
rect 69032 484362 69060 528526
rect 67824 484356 67876 484362
rect 67824 484298 67876 484304
rect 69020 484356 69072 484362
rect 69020 484298 69072 484304
rect 67730 479496 67786 479505
rect 67730 479431 67786 479440
rect 67640 463072 67692 463078
rect 67640 463014 67692 463020
rect 67376 441586 67496 441614
rect 67376 440298 67404 441586
rect 67364 440292 67416 440298
rect 67364 440234 67416 440240
rect 67272 435396 67324 435402
rect 67272 435338 67324 435344
rect 67284 427417 67312 435338
rect 67270 427408 67326 427417
rect 67270 427343 67326 427352
rect 67270 426320 67326 426329
rect 67270 426255 67326 426264
rect 67284 425746 67312 426255
rect 67272 425740 67324 425746
rect 67272 425682 67324 425688
rect 67376 405657 67404 440234
rect 67546 432576 67602 432585
rect 67546 432511 67602 432520
rect 67560 432002 67588 432511
rect 67548 431996 67600 432002
rect 67548 431938 67600 431944
rect 67548 428392 67600 428398
rect 67548 428334 67600 428340
rect 67560 426329 67588 428334
rect 67546 426320 67602 426329
rect 67546 426255 67602 426264
rect 67640 418804 67692 418810
rect 67640 418746 67692 418752
rect 67454 418160 67510 418169
rect 67454 418095 67510 418104
rect 67362 405648 67418 405657
rect 67362 405583 67418 405592
rect 67178 402656 67234 402665
rect 67178 402591 67234 402600
rect 67192 401713 67220 402591
rect 67178 401704 67234 401713
rect 66260 401668 66312 401674
rect 67178 401639 67234 401648
rect 66260 401610 66312 401616
rect 66168 384940 66220 384946
rect 66168 384882 66220 384888
rect 66272 292574 66300 401610
rect 66718 401568 66774 401577
rect 66718 401503 66774 401512
rect 66732 400246 66760 401503
rect 66720 400240 66772 400246
rect 66720 400182 66772 400188
rect 66810 399664 66866 399673
rect 66810 399599 66866 399608
rect 66824 396778 66852 399599
rect 67180 397520 67232 397526
rect 67178 397488 67180 397497
rect 67232 397488 67234 397497
rect 67178 397423 67234 397432
rect 66812 396772 66864 396778
rect 66812 396714 66864 396720
rect 67180 396024 67232 396030
rect 67180 395966 67232 395972
rect 67192 395321 67220 395966
rect 67178 395312 67234 395321
rect 67178 395247 67234 395256
rect 67364 393304 67416 393310
rect 67364 393246 67416 393252
rect 66810 392320 66866 392329
rect 66810 392255 66866 392264
rect 66824 392018 66852 392255
rect 66812 392012 66864 392018
rect 66812 391954 66864 391960
rect 67376 387297 67404 393246
rect 67362 387288 67418 387297
rect 67362 387223 67418 387232
rect 67468 347818 67496 418095
rect 67652 417081 67680 418746
rect 67638 417072 67694 417081
rect 67638 417007 67694 417016
rect 67546 400480 67602 400489
rect 67546 400415 67602 400424
rect 67560 379438 67588 400415
rect 67836 396409 67864 484298
rect 70308 469872 70360 469878
rect 70308 469814 70360 469820
rect 69662 466576 69718 466585
rect 69662 466511 69718 466520
rect 69676 439006 69704 466511
rect 70320 445641 70348 469814
rect 69754 445632 69810 445641
rect 69754 445567 69810 445576
rect 70306 445632 70362 445641
rect 70306 445567 70362 445576
rect 69664 439000 69716 439006
rect 69664 438942 69716 438948
rect 68284 438932 68336 438938
rect 68284 438874 68336 438880
rect 68006 434752 68062 434761
rect 68006 434687 68062 434696
rect 67822 396400 67878 396409
rect 67822 396335 67878 396344
rect 67652 393446 67680 393477
rect 67640 393440 67692 393446
rect 67638 393408 67640 393417
rect 67692 393408 67694 393417
rect 67638 393343 67694 393352
rect 67652 393310 67680 393343
rect 67640 393304 67692 393310
rect 67640 393246 67692 393252
rect 67732 390584 67784 390590
rect 67732 390526 67784 390532
rect 67548 379432 67600 379438
rect 67548 379374 67600 379380
rect 67456 347812 67508 347818
rect 67456 347754 67508 347760
rect 66272 292546 66484 292574
rect 66166 287600 66222 287609
rect 66166 287535 66222 287544
rect 66180 287201 66208 287535
rect 66166 287192 66222 287201
rect 66166 287127 66222 287136
rect 66074 273184 66130 273193
rect 66074 273119 66130 273128
rect 66180 269113 66208 287127
rect 66258 282976 66314 282985
rect 66258 282911 66260 282920
rect 66312 282911 66314 282920
rect 66260 282882 66312 282888
rect 66456 275330 66484 292546
rect 67364 284368 67416 284374
rect 67364 284310 67416 284316
rect 67376 279721 67404 284310
rect 67362 279712 67418 279721
rect 67362 279647 67418 279656
rect 66812 279472 66864 279478
rect 66812 279414 66864 279420
rect 66824 278905 66852 279414
rect 66810 278896 66866 278905
rect 66810 278831 66866 278840
rect 66812 278724 66864 278730
rect 66812 278666 66864 278672
rect 66824 278089 66852 278666
rect 66810 278080 66866 278089
rect 66810 278015 66866 278024
rect 66812 277364 66864 277370
rect 66812 277306 66864 277312
rect 66824 276457 66852 277306
rect 66810 276448 66866 276457
rect 66810 276383 66866 276392
rect 66812 276004 66864 276010
rect 66812 275946 66864 275952
rect 66824 275641 66852 275946
rect 66810 275632 66866 275641
rect 66810 275567 66866 275576
rect 66444 275324 66496 275330
rect 66444 275266 66496 275272
rect 66720 275324 66772 275330
rect 66720 275266 66772 275272
rect 66732 274825 66760 275266
rect 66718 274816 66774 274825
rect 66718 274751 66774 274760
rect 66810 274000 66866 274009
rect 66810 273935 66866 273944
rect 66824 273358 66852 273935
rect 66812 273352 66864 273358
rect 66812 273294 66864 273300
rect 66810 272368 66866 272377
rect 66810 272303 66866 272312
rect 66824 271998 66852 272303
rect 66812 271992 66864 271998
rect 66812 271934 66864 271940
rect 66810 270736 66866 270745
rect 66810 270671 66866 270680
rect 66824 270638 66852 270671
rect 66812 270632 66864 270638
rect 66812 270574 66864 270580
rect 66628 270496 66680 270502
rect 66628 270438 66680 270444
rect 66640 269929 66668 270438
rect 66626 269920 66682 269929
rect 66626 269855 66682 269864
rect 66166 269104 66222 269113
rect 66166 269039 66222 269048
rect 66810 268288 66866 268297
rect 66810 268223 66866 268232
rect 66824 267782 66852 268223
rect 66812 267776 66864 267782
rect 66812 267718 66864 267724
rect 66810 266656 66866 266665
rect 66810 266591 66866 266600
rect 66824 266422 66852 266591
rect 66812 266416 66864 266422
rect 66812 266358 66864 266364
rect 66534 265024 66590 265033
rect 66534 264959 66536 264968
rect 66588 264959 66590 264968
rect 66536 264930 66588 264936
rect 66260 264240 66312 264246
rect 66260 264182 66312 264188
rect 66810 264208 66866 264217
rect 66272 260953 66300 264182
rect 66810 264143 66866 264152
rect 66824 263702 66852 264143
rect 66812 263696 66864 263702
rect 66812 263638 66864 263644
rect 67468 263401 67496 347754
rect 67546 289232 67602 289241
rect 67546 289167 67602 289176
rect 67560 282169 67588 289167
rect 67638 282840 67694 282849
rect 67638 282775 67694 282784
rect 67546 282160 67602 282169
rect 67546 282095 67602 282104
rect 67548 280220 67600 280226
rect 67548 280162 67600 280168
rect 67086 263392 67142 263401
rect 67086 263327 67142 263336
rect 67454 263392 67510 263401
rect 67454 263327 67510 263336
rect 66534 262576 66590 262585
rect 66534 262511 66590 262520
rect 66548 262274 66576 262511
rect 66536 262268 66588 262274
rect 66536 262210 66588 262216
rect 67100 261526 67128 263327
rect 67088 261520 67140 261526
rect 67088 261462 67140 261468
rect 66258 260944 66314 260953
rect 66258 260879 66314 260888
rect 66272 258738 66300 260879
rect 66536 260228 66588 260234
rect 66536 260170 66588 260176
rect 66548 260137 66576 260170
rect 66534 260128 66590 260137
rect 66534 260063 66590 260072
rect 66352 258800 66404 258806
rect 66352 258742 66404 258748
rect 66260 258732 66312 258738
rect 66260 258674 66312 258680
rect 66364 257990 66392 258742
rect 66444 258052 66496 258058
rect 66444 257994 66496 258000
rect 66352 257984 66404 257990
rect 66352 257926 66404 257932
rect 66456 257689 66484 257994
rect 66442 257680 66498 257689
rect 66442 257615 66498 257624
rect 66534 256728 66590 256737
rect 66534 256663 66590 256672
rect 66260 255468 66312 255474
rect 66260 255410 66312 255416
rect 66272 255377 66300 255410
rect 66258 255368 66314 255377
rect 66258 255303 66314 255312
rect 66076 251864 66128 251870
rect 66548 251841 66576 256663
rect 66812 255264 66864 255270
rect 66810 255232 66812 255241
rect 66864 255232 66866 255241
rect 66810 255167 66866 255176
rect 66812 254584 66864 254590
rect 66812 254526 66864 254532
rect 66824 254425 66852 254526
rect 66810 254416 66866 254425
rect 66810 254351 66866 254360
rect 66994 253600 67050 253609
rect 66994 253535 67050 253544
rect 67008 253230 67036 253535
rect 66996 253224 67048 253230
rect 66996 253166 67048 253172
rect 67364 253224 67416 253230
rect 67364 253166 67416 253172
rect 66626 251968 66682 251977
rect 66626 251903 66682 251912
rect 66640 251870 66668 251903
rect 66628 251864 66680 251870
rect 66076 251806 66128 251812
rect 66534 251832 66590 251841
rect 65984 240100 66036 240106
rect 65984 240042 66036 240048
rect 65892 228404 65944 228410
rect 65892 228346 65944 228352
rect 65720 171106 66024 171134
rect 65996 156670 66024 171106
rect 65984 156664 66036 156670
rect 65984 156606 66036 156612
rect 65892 153332 65944 153338
rect 65892 153274 65944 153280
rect 64788 152516 64840 152522
rect 64788 152458 64840 152464
rect 64788 135924 64840 135930
rect 64788 135866 64840 135872
rect 64696 120012 64748 120018
rect 64696 119954 64748 119960
rect 64604 115320 64656 115326
rect 64604 115262 64656 115268
rect 63500 108316 63552 108322
rect 63500 108258 63552 108264
rect 63512 107710 63540 108258
rect 63500 107704 63552 107710
rect 63500 107646 63552 107652
rect 64604 107704 64656 107710
rect 64604 107646 64656 107652
rect 63408 91044 63460 91050
rect 63408 90986 63460 90992
rect 64616 88233 64644 107646
rect 64696 100020 64748 100026
rect 64696 99962 64748 99968
rect 64602 88224 64658 88233
rect 64602 88159 64658 88168
rect 64708 78674 64736 99962
rect 64800 94489 64828 135866
rect 65904 130665 65932 153274
rect 65890 130656 65946 130665
rect 65890 130591 65946 130600
rect 65996 122233 66024 156606
rect 66088 136678 66116 251806
rect 66628 251806 66680 251812
rect 66534 251767 66590 251776
rect 66812 250776 66864 250782
rect 66812 250718 66864 250724
rect 66824 250345 66852 250718
rect 66810 250336 66866 250345
rect 66810 250271 66866 250280
rect 66810 248704 66866 248713
rect 66810 248639 66866 248648
rect 66824 248470 66852 248639
rect 66812 248464 66864 248470
rect 66812 248406 66864 248412
rect 66534 247888 66590 247897
rect 66534 247823 66590 247832
rect 66548 247110 66576 247823
rect 66536 247104 66588 247110
rect 66536 247046 66588 247052
rect 66810 245440 66866 245449
rect 66810 245375 66866 245384
rect 66824 244322 66852 245375
rect 66812 244316 66864 244322
rect 66812 244258 66864 244264
rect 66720 244248 66772 244254
rect 66720 244190 66772 244196
rect 66732 243001 66760 244190
rect 66902 243808 66958 243817
rect 66902 243743 66958 243752
rect 66718 242992 66774 243001
rect 66916 242962 66944 243743
rect 66718 242927 66774 242936
rect 66904 242956 66956 242962
rect 66904 242898 66956 242904
rect 66810 242176 66866 242185
rect 66810 242111 66866 242120
rect 66824 241602 66852 242111
rect 66812 241596 66864 241602
rect 66812 241538 66864 241544
rect 67376 238241 67404 253166
rect 67454 246256 67510 246265
rect 67454 246191 67510 246200
rect 67362 238232 67418 238241
rect 67362 238167 67418 238176
rect 67376 144974 67404 238167
rect 67468 231742 67496 246191
rect 67456 231736 67508 231742
rect 67456 231678 67508 231684
rect 67364 144968 67416 144974
rect 67364 144910 67416 144916
rect 66166 140856 66222 140865
rect 66166 140791 66222 140800
rect 66076 136672 66128 136678
rect 66076 136614 66128 136620
rect 65982 122224 66038 122233
rect 65982 122159 66038 122168
rect 65982 108624 66038 108633
rect 65982 108559 66038 108568
rect 65892 105596 65944 105602
rect 65892 105538 65944 105544
rect 64786 94480 64842 94489
rect 64786 94415 64842 94424
rect 65904 84153 65932 105538
rect 65890 84144 65946 84153
rect 65890 84079 65946 84088
rect 64696 78668 64748 78674
rect 64696 78610 64748 78616
rect 65996 77081 66024 108559
rect 66088 102649 66116 136614
rect 66074 102640 66130 102649
rect 66074 102575 66130 102584
rect 66076 101448 66128 101454
rect 66076 101390 66128 101396
rect 65982 77072 66038 77081
rect 65982 77007 66038 77016
rect 66088 75818 66116 101390
rect 66180 90982 66208 140791
rect 66352 133204 66404 133210
rect 66352 133146 66404 133152
rect 66364 131209 66392 133146
rect 66904 132456 66956 132462
rect 66904 132398 66956 132404
rect 66916 132025 66944 132398
rect 66902 132016 66958 132025
rect 66902 131951 66958 131960
rect 66350 131200 66406 131209
rect 66350 131135 66406 131144
rect 66904 128308 66956 128314
rect 66904 128250 66956 128256
rect 66916 127673 66944 128250
rect 66902 127664 66958 127673
rect 66902 127599 66958 127608
rect 66812 126948 66864 126954
rect 66812 126890 66864 126896
rect 66720 126880 66772 126886
rect 66824 126857 66852 126890
rect 66720 126822 66772 126828
rect 66810 126848 66866 126857
rect 66732 126041 66760 126822
rect 66810 126783 66866 126792
rect 66718 126032 66774 126041
rect 66718 125967 66774 125976
rect 66628 124840 66680 124846
rect 66628 124782 66680 124788
rect 66260 124160 66312 124166
rect 66260 124102 66312 124108
rect 66272 123865 66300 124102
rect 66258 123856 66314 123865
rect 66258 123791 66314 123800
rect 66640 123049 66668 124782
rect 66626 123040 66682 123049
rect 66626 122975 66682 122984
rect 66904 121440 66956 121446
rect 66810 121408 66866 121417
rect 66904 121382 66956 121388
rect 66810 121343 66812 121352
rect 66864 121343 66866 121352
rect 66812 121314 66864 121320
rect 66916 120601 66944 121382
rect 66902 120592 66958 120601
rect 66902 120527 66958 120536
rect 66904 120080 66956 120086
rect 66810 120048 66866 120057
rect 66904 120022 66956 120028
rect 66810 119983 66812 119992
rect 66864 119983 66866 119992
rect 66812 119954 66864 119960
rect 66916 119241 66944 120022
rect 66902 119232 66958 119241
rect 66902 119167 66958 119176
rect 66720 118652 66772 118658
rect 66720 118594 66772 118600
rect 66732 117609 66760 118594
rect 66718 117600 66774 117609
rect 66718 117535 66774 117544
rect 66812 117292 66864 117298
rect 66812 117234 66864 117240
rect 66260 117224 66312 117230
rect 66260 117166 66312 117172
rect 66272 116249 66300 117166
rect 66824 117065 66852 117234
rect 66810 117056 66866 117065
rect 66810 116991 66866 117000
rect 66258 116240 66314 116249
rect 66258 116175 66314 116184
rect 66904 115932 66956 115938
rect 66904 115874 66956 115880
rect 66916 115433 66944 115874
rect 66902 115424 66958 115433
rect 66902 115359 66958 115368
rect 66812 115320 66864 115326
rect 66812 115262 66864 115268
rect 66824 114617 66852 115262
rect 66810 114608 66866 114617
rect 66810 114543 66866 114552
rect 66812 114504 66864 114510
rect 66812 114446 66864 114452
rect 66824 113801 66852 114446
rect 66904 114436 66956 114442
rect 66904 114378 66956 114384
rect 66810 113792 66866 113801
rect 66810 113727 66866 113736
rect 66916 113257 66944 114378
rect 66902 113248 66958 113257
rect 66902 113183 66958 113192
rect 66812 112464 66864 112470
rect 66812 112406 66864 112412
rect 66824 111625 66852 112406
rect 66810 111616 66866 111625
rect 66810 111551 66866 111560
rect 66810 110800 66866 110809
rect 66810 110735 66866 110744
rect 66824 110498 66852 110735
rect 66812 110492 66864 110498
rect 66812 110434 66864 110440
rect 66810 110256 66866 110265
rect 66810 110191 66866 110200
rect 66824 109070 66852 110191
rect 66812 109064 66864 109070
rect 66812 109006 66864 109012
rect 66810 107808 66866 107817
rect 66810 107743 66866 107752
rect 66824 107710 66852 107743
rect 66812 107704 66864 107710
rect 66812 107646 66864 107652
rect 66810 106992 66866 107001
rect 66810 106927 66866 106936
rect 66824 106350 66852 106927
rect 66812 106344 66864 106350
rect 66812 106286 66864 106292
rect 66534 105632 66590 105641
rect 66534 105567 66536 105576
rect 66588 105567 66590 105576
rect 66536 105538 66588 105544
rect 66812 104848 66864 104854
rect 66810 104816 66812 104825
rect 66864 104816 66866 104825
rect 66810 104751 66866 104760
rect 67376 104009 67404 144910
rect 67362 104000 67418 104009
rect 67362 103935 67418 103944
rect 66812 103488 66864 103494
rect 66812 103430 66864 103436
rect 66824 103193 66852 103430
rect 66810 103184 66866 103193
rect 66810 103119 66866 103128
rect 66626 101824 66682 101833
rect 66626 101759 66682 101768
rect 66640 101454 66668 101759
rect 66628 101448 66680 101454
rect 66628 101390 66680 101396
rect 67362 100192 67418 100201
rect 67362 100127 67418 100136
rect 66812 100020 66864 100026
rect 66812 99962 66864 99968
rect 66824 99657 66852 99962
rect 66810 99648 66866 99657
rect 66810 99583 66866 99592
rect 66812 99340 66864 99346
rect 66812 99282 66864 99288
rect 66824 98841 66852 99282
rect 66810 98832 66866 98841
rect 66810 98767 66866 98776
rect 66442 96384 66498 96393
rect 66442 96319 66498 96328
rect 66456 95946 66484 96319
rect 66444 95940 66496 95946
rect 66444 95882 66496 95888
rect 66812 95192 66864 95198
rect 66812 95134 66864 95140
rect 66824 95033 66852 95134
rect 66810 95024 66866 95033
rect 66810 94959 66866 94968
rect 66994 93392 67050 93401
rect 66994 93327 67050 93336
rect 67008 92614 67036 93327
rect 66996 92608 67048 92614
rect 66996 92550 67048 92556
rect 67272 92608 67324 92614
rect 67272 92550 67324 92556
rect 66168 90976 66220 90982
rect 66168 90918 66220 90924
rect 65616 75812 65668 75818
rect 65616 75754 65668 75760
rect 66076 75812 66128 75818
rect 66076 75754 66128 75760
rect 62026 72448 62082 72457
rect 62026 72383 62082 72392
rect 61936 71732 61988 71738
rect 61936 71674 61988 71680
rect 61936 51740 61988 51746
rect 61936 51682 61988 51688
rect 59268 49020 59320 49026
rect 59268 48962 59320 48968
rect 59280 3534 59308 48962
rect 61948 16574 61976 51682
rect 61856 16546 61976 16574
rect 59636 7608 59688 7614
rect 59636 7550 59688 7556
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 7550
rect 60832 3596 60884 3602
rect 60832 3538 60884 3544
rect 60844 480 60872 3538
rect 61856 3482 61884 16546
rect 62040 6914 62068 72383
rect 65524 47592 65576 47598
rect 65524 47534 65576 47540
rect 64788 32428 64840 32434
rect 64788 32370 64840 32376
rect 61948 6886 62068 6914
rect 61948 3602 61976 6886
rect 61936 3596 61988 3602
rect 61936 3538 61988 3544
rect 64800 3534 64828 32370
rect 65536 6914 65564 47534
rect 65628 46238 65656 75754
rect 67284 60722 67312 92550
rect 67376 86902 67404 100127
rect 67468 97209 67496 231678
rect 67560 129849 67588 280162
rect 67652 277273 67680 282775
rect 67638 277264 67694 277273
rect 67638 277199 67694 277208
rect 67652 276078 67680 277199
rect 67640 276072 67692 276078
rect 67640 276014 67692 276020
rect 67744 242554 67772 390526
rect 67836 371249 67864 396335
rect 67914 395312 67970 395321
rect 67914 395247 67970 395256
rect 67928 372609 67956 395247
rect 67914 372600 67970 372609
rect 67914 372535 67970 372544
rect 67822 371240 67878 371249
rect 67822 371175 67878 371184
rect 68020 282985 68048 434687
rect 68296 428398 68324 438874
rect 68928 437164 68980 437170
rect 68928 437106 68980 437112
rect 68940 436150 68968 437106
rect 69676 436370 69704 438942
rect 69768 437170 69796 445567
rect 70504 443562 70532 528526
rect 71056 497486 71084 536794
rect 71792 525094 71820 539158
rect 71872 539096 71924 539102
rect 71872 539038 71924 539044
rect 71780 525088 71832 525094
rect 71780 525030 71832 525036
rect 71044 497480 71096 497486
rect 71044 497422 71096 497428
rect 71042 453112 71098 453121
rect 71042 453047 71098 453056
rect 70492 443556 70544 443562
rect 70492 443498 70544 443504
rect 70400 442264 70452 442270
rect 70400 442206 70452 442212
rect 70412 441614 70440 442206
rect 70412 441586 70624 441614
rect 69756 437164 69808 437170
rect 69756 437106 69808 437112
rect 69676 436342 69796 436370
rect 68928 436144 68980 436150
rect 68928 436086 68980 436092
rect 69664 436144 69716 436150
rect 69664 436086 69716 436092
rect 68940 434194 68968 436086
rect 69202 434344 69258 434353
rect 69676 434330 69704 436086
rect 69258 434302 69704 434330
rect 69768 434330 69796 436342
rect 70596 434790 70624 441586
rect 71056 436150 71084 453047
rect 71136 445800 71188 445806
rect 71136 445742 71188 445748
rect 71044 436144 71096 436150
rect 71044 436086 71096 436092
rect 70584 434784 70636 434790
rect 70584 434726 70636 434732
rect 70596 434330 70624 434726
rect 69768 434302 70288 434330
rect 70596 434302 71024 434330
rect 69202 434279 69258 434288
rect 68816 434166 68968 434194
rect 71148 433702 71176 445742
rect 71688 437436 71740 437442
rect 71688 437378 71740 437384
rect 71226 434888 71282 434897
rect 71226 434823 71282 434832
rect 71240 434625 71268 434823
rect 71226 434616 71282 434625
rect 71226 434551 71282 434560
rect 71700 434330 71728 437378
rect 71884 436121 71912 539038
rect 73448 538214 73476 539158
rect 73632 539158 74336 539186
rect 74552 539158 75256 539186
rect 75932 539158 76176 539186
rect 73448 538186 73568 538214
rect 73540 536790 73568 538186
rect 73528 536784 73580 536790
rect 73528 536726 73580 536732
rect 73540 536110 73568 536726
rect 73528 536104 73580 536110
rect 73528 536046 73580 536052
rect 73632 528554 73660 539158
rect 73172 528526 73660 528554
rect 73172 493338 73200 528526
rect 73160 493332 73212 493338
rect 73160 493274 73212 493280
rect 72424 455524 72476 455530
rect 72424 455466 72476 455472
rect 72436 437442 72464 455466
rect 73804 449880 73856 449886
rect 73804 449822 73856 449828
rect 72424 437436 72476 437442
rect 72424 437378 72476 437384
rect 71870 436112 71926 436121
rect 71870 436047 71926 436056
rect 72698 436112 72754 436121
rect 72698 436047 72754 436056
rect 72606 435296 72662 435305
rect 72606 435231 72662 435240
rect 72620 434330 72648 435231
rect 71576 434302 71728 434330
rect 72312 434302 72648 434330
rect 72712 434330 72740 436047
rect 73816 434761 73844 449822
rect 74552 448594 74580 539158
rect 75932 459649 75960 539158
rect 75918 459640 75974 459649
rect 75918 459575 75974 459584
rect 76576 458833 76604 539650
rect 86592 539640 86644 539646
rect 76746 539608 76802 539617
rect 76802 539566 77096 539594
rect 86592 539582 86644 539588
rect 76746 539543 76802 539552
rect 76760 533390 76788 539543
rect 78016 539158 78352 539186
rect 77944 536104 77996 536110
rect 77944 536046 77996 536052
rect 76748 533384 76800 533390
rect 76748 533326 76800 533332
rect 77956 487830 77984 536046
rect 78324 533390 78352 539158
rect 78692 539158 78936 539186
rect 80040 539158 80100 539186
rect 78312 533384 78364 533390
rect 78312 533326 78364 533332
rect 77944 487824 77996 487830
rect 77944 487766 77996 487772
rect 77300 482316 77352 482322
rect 77300 482258 77352 482264
rect 77208 458856 77260 458862
rect 76562 458824 76618 458833
rect 77208 458798 77260 458804
rect 76562 458759 76618 458768
rect 76564 454096 76616 454102
rect 76564 454038 76616 454044
rect 74540 448588 74592 448594
rect 74540 448530 74592 448536
rect 75828 448588 75880 448594
rect 75828 448530 75880 448536
rect 75840 447846 75868 448530
rect 75828 447840 75880 447846
rect 75828 447782 75880 447788
rect 74816 437504 74868 437510
rect 74816 437446 74868 437452
rect 74080 436484 74132 436490
rect 74080 436426 74132 436432
rect 73802 434752 73858 434761
rect 73802 434687 73858 434696
rect 74092 434330 74120 436426
rect 74170 434752 74226 434761
rect 74170 434687 74226 434696
rect 72712 434302 73048 434330
rect 73784 434302 74120 434330
rect 74184 434330 74212 434687
rect 74828 434330 74856 437446
rect 76576 436490 76604 454038
rect 77220 441614 77248 458798
rect 76944 441586 77248 441614
rect 76564 436484 76616 436490
rect 76564 436426 76616 436432
rect 75828 436144 75880 436150
rect 75828 436086 75880 436092
rect 75840 435441 75868 436086
rect 75826 435432 75882 435441
rect 75826 435367 75882 435376
rect 76378 434344 76434 434353
rect 74184 434302 74336 434330
rect 74828 434302 75072 434330
rect 76944 434330 76972 441586
rect 77312 434602 77340 482258
rect 78692 461650 78720 539158
rect 80072 536110 80100 539158
rect 80164 539158 80960 539186
rect 81452 539158 81880 539186
rect 82800 539158 82860 539186
rect 80060 536104 80112 536110
rect 80060 536046 80112 536052
rect 80164 528554 80192 539158
rect 80704 536172 80756 536178
rect 80704 536114 80756 536120
rect 80072 528526 80192 528554
rect 80072 463010 80100 528526
rect 80716 486470 80744 536114
rect 80704 486464 80756 486470
rect 80704 486406 80756 486412
rect 81452 472569 81480 539158
rect 82832 536178 82860 539158
rect 82924 539158 83720 539186
rect 84212 539158 84640 539186
rect 85560 539158 85620 539186
rect 82820 536172 82872 536178
rect 82820 536114 82872 536120
rect 82924 528554 82952 539158
rect 83464 534744 83516 534750
rect 83464 534686 83516 534692
rect 82832 528526 82952 528554
rect 81438 472560 81494 472569
rect 81438 472495 81494 472504
rect 81348 463072 81400 463078
rect 81348 463014 81400 463020
rect 80060 463004 80112 463010
rect 80060 462946 80112 462952
rect 78680 461644 78732 461650
rect 78680 461586 78732 461592
rect 81360 459610 81388 463014
rect 81348 459604 81400 459610
rect 81348 459546 81400 459552
rect 78680 456816 78732 456822
rect 78680 456758 78732 456764
rect 77390 454064 77446 454073
rect 77390 453999 77446 454008
rect 77404 441614 77432 453999
rect 78692 441614 78720 456758
rect 77404 441586 78168 441614
rect 78692 441586 78904 441614
rect 76434 434302 76972 434330
rect 77266 434574 77340 434602
rect 76378 434279 76434 434288
rect 77114 433800 77170 433809
rect 77266 433786 77294 434574
rect 78140 434330 78168 441586
rect 78876 434330 78904 441586
rect 80980 437368 81032 437374
rect 80980 437310 81032 437316
rect 80992 436257 81020 437310
rect 80978 436248 81034 436257
rect 80978 436183 81034 436192
rect 80428 436144 80480 436150
rect 80334 436112 80390 436121
rect 80428 436086 80480 436092
rect 80334 436047 80390 436056
rect 80348 434330 80376 436047
rect 78140 434302 78568 434330
rect 78876 434302 79304 434330
rect 80040 434302 80376 434330
rect 80440 434330 80468 436086
rect 80992 434330 81020 436183
rect 81360 436121 81388 459546
rect 82832 455394 82860 528526
rect 82820 455388 82872 455394
rect 82820 455330 82872 455336
rect 82728 451988 82780 451994
rect 82728 451930 82780 451936
rect 82740 441614 82768 451930
rect 82464 441586 82768 441614
rect 81346 436112 81402 436121
rect 81346 436047 81402 436056
rect 81898 434344 81954 434353
rect 80440 434302 80592 434330
rect 80992 434302 81328 434330
rect 82464 434330 82492 441586
rect 82818 439648 82874 439657
rect 82818 439583 82874 439592
rect 82832 437442 82860 439583
rect 83476 439006 83504 534686
rect 84212 529242 84240 539158
rect 84200 529236 84252 529242
rect 84200 529178 84252 529184
rect 85592 494766 85620 539158
rect 85684 539158 86480 539186
rect 85684 522442 85712 539158
rect 86604 528554 86632 539582
rect 86236 528526 86632 528554
rect 86972 539158 87400 539186
rect 88320 539158 88472 539186
rect 85672 522436 85724 522442
rect 85672 522378 85724 522384
rect 85672 522300 85724 522306
rect 85672 522242 85724 522248
rect 85580 494760 85632 494766
rect 85580 494702 85632 494708
rect 85580 476808 85632 476814
rect 85580 476750 85632 476756
rect 85488 469260 85540 469266
rect 85488 469202 85540 469208
rect 85500 441614 85528 469202
rect 85224 441586 85528 441614
rect 83464 439000 83516 439006
rect 83464 438942 83516 438948
rect 83740 439000 83792 439006
rect 83740 438942 83792 438948
rect 82820 437436 82872 437442
rect 82820 437378 82872 437384
rect 83094 436112 83150 436121
rect 83094 436047 83150 436056
rect 83108 434353 83136 436047
rect 83094 434344 83150 434353
rect 81954 434302 82492 434330
rect 82800 434302 83094 434330
rect 81898 434279 81954 434288
rect 83752 434330 83780 438942
rect 83924 437436 83976 437442
rect 83924 437378 83976 437384
rect 83536 434302 83780 434330
rect 83094 434279 83150 434288
rect 83108 434219 83136 434279
rect 83830 434072 83886 434081
rect 83936 434058 83964 437378
rect 84658 434344 84714 434353
rect 85224 434330 85252 441586
rect 85592 436370 85620 476750
rect 85684 441614 85712 522242
rect 86236 469266 86264 528526
rect 86224 469260 86276 469266
rect 86224 469202 86276 469208
rect 86222 449984 86278 449993
rect 86222 449919 86278 449928
rect 85684 441586 85896 441614
rect 85592 436342 85712 436370
rect 84714 434302 85252 434330
rect 84658 434279 84714 434288
rect 83886 434030 84088 434058
rect 83830 434007 83886 434016
rect 85684 433922 85712 436342
rect 85868 434353 85896 441586
rect 86236 437374 86264 449919
rect 86972 446457 87000 539158
rect 87604 536172 87656 536178
rect 87604 536114 87656 536120
rect 87616 460902 87644 536114
rect 88444 534857 88472 539158
rect 88536 539158 89240 539186
rect 90160 539158 90404 539186
rect 88430 534848 88486 534857
rect 88430 534783 88486 534792
rect 88536 528554 88564 539158
rect 90376 536761 90404 539158
rect 90362 536752 90418 536761
rect 90362 536687 90418 536696
rect 88984 535492 89036 535498
rect 88984 535434 89036 535440
rect 88352 528526 88564 528554
rect 88352 461553 88380 528526
rect 88996 482322 89024 535434
rect 88984 482316 89036 482322
rect 88984 482258 89036 482264
rect 88338 461544 88394 461553
rect 88338 461479 88394 461488
rect 87604 460896 87656 460902
rect 87604 460838 87656 460844
rect 90376 458862 90404 536687
rect 90914 476776 90970 476785
rect 90914 476711 90970 476720
rect 90928 473414 90956 476711
rect 90916 473408 90968 473414
rect 90916 473350 90968 473356
rect 90364 458856 90416 458862
rect 90364 458798 90416 458804
rect 87604 451920 87656 451926
rect 87604 451862 87656 451868
rect 86958 446448 87014 446457
rect 86958 446383 87014 446392
rect 87616 437442 87644 451862
rect 88522 449984 88578 449993
rect 88522 449919 88578 449928
rect 88248 445052 88300 445058
rect 88248 444994 88300 445000
rect 87604 437436 87656 437442
rect 87604 437378 87656 437384
rect 86224 437368 86276 437374
rect 86224 437310 86276 437316
rect 88260 436354 88288 444994
rect 88536 444446 88564 449919
rect 88524 444440 88576 444446
rect 88524 444382 88576 444388
rect 88536 441614 88564 444382
rect 88536 441586 88656 441614
rect 87328 436348 87380 436354
rect 87328 436290 87380 436296
rect 88248 436348 88300 436354
rect 88248 436290 88300 436296
rect 85854 434344 85910 434353
rect 87340 434330 87368 436290
rect 85910 434302 86296 434330
rect 87032 434302 87368 434330
rect 88628 434330 88656 441586
rect 90928 437442 90956 473350
rect 91020 445058 91048 539786
rect 94318 539744 94374 539753
rect 94318 539679 94374 539688
rect 94332 539646 94360 539679
rect 94320 539640 94372 539646
rect 94320 539582 94372 539588
rect 91112 539158 91264 539186
rect 91572 539158 92184 539186
rect 93104 539158 93440 539186
rect 94024 539158 94544 539186
rect 91112 535498 91140 539158
rect 91100 535492 91152 535498
rect 91100 535434 91152 535440
rect 91572 528554 91600 539158
rect 93412 536178 93440 539158
rect 93950 538928 94006 538937
rect 93950 538863 94006 538872
rect 93964 538286 93992 538863
rect 93952 538280 94004 538286
rect 93952 538222 94004 538228
rect 93400 536172 93452 536178
rect 93400 536114 93452 536120
rect 93124 536104 93176 536110
rect 93124 536046 93176 536052
rect 91204 528526 91600 528554
rect 91204 469878 91232 528526
rect 92572 490612 92624 490618
rect 92572 490554 92624 490560
rect 91192 469872 91244 469878
rect 91192 469814 91244 469820
rect 91744 461644 91796 461650
rect 91744 461586 91796 461592
rect 91008 445052 91060 445058
rect 91008 444994 91060 445000
rect 90916 437436 90968 437442
rect 90916 437378 90968 437384
rect 91756 436762 91784 461586
rect 91744 436756 91796 436762
rect 91744 436698 91796 436704
rect 92584 434602 92612 490554
rect 93136 480962 93164 536046
rect 94516 526454 94544 539158
rect 94504 526448 94556 526454
rect 94504 526390 94556 526396
rect 93124 480956 93176 480962
rect 93124 480898 93176 480904
rect 94516 473346 94544 526390
rect 94700 520985 94728 563615
rect 95148 525836 95200 525842
rect 95148 525778 95200 525784
rect 94686 520976 94742 520985
rect 94686 520911 94742 520920
rect 94504 473340 94556 473346
rect 94504 473282 94556 473288
rect 95056 473340 95108 473346
rect 95056 473282 95108 473288
rect 95068 472054 95096 473282
rect 95056 472048 95108 472054
rect 95056 471990 95108 471996
rect 93860 467900 93912 467906
rect 93860 467842 93912 467848
rect 93872 434602 93900 467842
rect 95068 437646 95096 471990
rect 95160 467906 95188 525778
rect 95252 476814 95280 574767
rect 95896 567866 95924 582354
rect 95884 567860 95936 567866
rect 95884 567802 95936 567808
rect 95330 567216 95386 567225
rect 95330 567151 95386 567160
rect 95344 523705 95372 567151
rect 96632 556986 96660 702850
rect 96712 587172 96764 587178
rect 96712 587114 96764 587120
rect 96724 576854 96752 587114
rect 97264 584452 97316 584458
rect 97264 584394 97316 584400
rect 97170 578912 97226 578921
rect 97170 578847 97226 578856
rect 97184 578270 97212 578847
rect 97172 578264 97224 578270
rect 97172 578206 97224 578212
rect 96724 576826 96936 576854
rect 96710 565856 96766 565865
rect 96710 565791 96766 565800
rect 96724 557534 96752 565791
rect 96802 562320 96858 562329
rect 96802 562255 96858 562264
rect 96816 561746 96844 562255
rect 96804 561740 96856 561746
rect 96804 561682 96856 561688
rect 96802 560960 96858 560969
rect 96802 560895 96858 560904
rect 96816 560318 96844 560895
rect 96804 560312 96856 560318
rect 96804 560254 96856 560260
rect 96908 558793 96936 576826
rect 96986 573472 97042 573481
rect 96986 573407 97042 573416
rect 97000 572762 97028 573407
rect 96988 572756 97040 572762
rect 96988 572698 97040 572704
rect 97276 570722 97304 584394
rect 101402 583944 101458 583953
rect 101402 583879 101458 583888
rect 97906 577552 97962 577561
rect 97962 577510 98040 577538
rect 97906 577487 97962 577496
rect 98012 576910 98040 577510
rect 98000 576904 98052 576910
rect 98000 576846 98052 576852
rect 97908 576768 97960 576774
rect 97906 576736 97908 576745
rect 97960 576736 97962 576745
rect 97906 576671 97962 576680
rect 97538 572112 97594 572121
rect 97538 572047 97594 572056
rect 97552 571402 97580 572047
rect 97540 571396 97592 571402
rect 97540 571338 97592 571344
rect 97264 570716 97316 570722
rect 97264 570658 97316 570664
rect 97276 569265 97304 570658
rect 97906 570072 97962 570081
rect 97906 570007 97962 570016
rect 97920 569974 97948 570007
rect 97908 569968 97960 569974
rect 97908 569910 97960 569916
rect 97262 569256 97318 569265
rect 97262 569191 97318 569200
rect 97078 559600 97134 559609
rect 97078 559535 97134 559544
rect 97092 559026 97120 559535
rect 97080 559020 97132 559026
rect 97080 558962 97132 558968
rect 96894 558784 96950 558793
rect 96894 558719 96950 558728
rect 97906 558784 97962 558793
rect 97906 558719 97962 558728
rect 97920 558210 97948 558719
rect 97908 558204 97960 558210
rect 97908 558146 97960 558152
rect 96724 557506 96844 557534
rect 96620 556980 96672 556986
rect 96620 556922 96672 556928
rect 96618 556880 96674 556889
rect 96618 556815 96674 556824
rect 95422 552528 95478 552537
rect 95422 552463 95478 552472
rect 95436 525842 95464 552463
rect 96632 551886 96660 556815
rect 96710 555520 96766 555529
rect 96710 555455 96766 555464
rect 96724 554810 96752 555455
rect 96712 554804 96764 554810
rect 96712 554746 96764 554752
rect 96816 554690 96844 557506
rect 97080 556980 97132 556986
rect 97080 556922 97132 556928
rect 96724 554662 96844 554690
rect 96620 551880 96672 551886
rect 96620 551822 96672 551828
rect 96724 547874 96752 554662
rect 96894 554160 96950 554169
rect 96894 554095 96950 554104
rect 96908 551970 96936 554095
rect 96986 552800 97042 552809
rect 96986 552735 97042 552744
rect 97000 552090 97028 552735
rect 97092 552537 97120 556922
rect 97078 552528 97134 552537
rect 97078 552463 97134 552472
rect 96988 552084 97040 552090
rect 96988 552026 97040 552032
rect 96908 551942 97028 551970
rect 96896 551880 96948 551886
rect 96896 551822 96948 551828
rect 96724 547846 96844 547874
rect 96710 545728 96766 545737
rect 96710 545663 96766 545672
rect 96618 541648 96674 541657
rect 96618 541583 96674 541592
rect 96632 541006 96660 541583
rect 96620 541000 96672 541006
rect 96620 540942 96672 540948
rect 95424 525836 95476 525842
rect 95424 525778 95476 525784
rect 95330 523696 95386 523705
rect 95330 523631 95386 523640
rect 95240 476808 95292 476814
rect 95240 476750 95292 476756
rect 96724 468489 96752 545663
rect 96816 539850 96844 547846
rect 96804 539844 96856 539850
rect 96804 539786 96856 539792
rect 96908 532030 96936 551822
rect 96896 532024 96948 532030
rect 96896 531966 96948 531972
rect 96710 468480 96766 468489
rect 96710 468415 96766 468424
rect 95148 467900 95200 467906
rect 95148 467842 95200 467848
rect 95240 458312 95292 458318
rect 95240 458254 95292 458260
rect 95056 437640 95108 437646
rect 95056 437582 95108 437588
rect 94228 437436 94280 437442
rect 94228 437378 94280 437384
rect 92538 434574 92612 434602
rect 93826 434574 93900 434602
rect 88628 434302 89056 434330
rect 85854 434279 85910 434288
rect 85868 434219 85896 434279
rect 92538 434194 92566 434574
rect 93826 434316 93854 434574
rect 94240 434330 94268 437378
rect 95252 434602 95280 458254
rect 95330 442232 95386 442241
rect 95330 442167 95386 442176
rect 95344 441614 95372 442167
rect 97000 441614 97028 551942
rect 97446 549400 97502 549409
rect 97446 549335 97448 549344
rect 97500 549335 97502 549344
rect 97448 549306 97500 549312
rect 97078 544368 97134 544377
rect 97078 544303 97134 544312
rect 97092 543794 97120 544303
rect 97080 543788 97132 543794
rect 97080 543730 97132 543736
rect 97078 543008 97134 543017
rect 97078 542943 97134 542952
rect 97092 542434 97120 542943
rect 97080 542428 97132 542434
rect 97080 542370 97132 542376
rect 98012 530602 98040 576846
rect 100852 572756 100904 572762
rect 100852 572698 100904 572704
rect 99380 571396 99432 571402
rect 99380 571338 99432 571344
rect 98736 570716 98788 570722
rect 98736 570658 98788 570664
rect 98644 536172 98696 536178
rect 98644 536114 98696 536120
rect 98000 530596 98052 530602
rect 98000 530538 98052 530544
rect 98000 455456 98052 455462
rect 98000 455398 98052 455404
rect 95344 441586 95648 441614
rect 95620 436801 95648 441586
rect 96908 441586 97028 441614
rect 95606 436792 95662 436801
rect 95606 436727 95662 436736
rect 95252 434574 95326 434602
rect 94240 434302 94576 434330
rect 95298 434316 95326 434574
rect 95620 434330 95648 436727
rect 96908 436121 96936 441586
rect 96988 437640 97040 437646
rect 96988 437582 97040 437588
rect 96894 436112 96950 436121
rect 96894 436047 96950 436056
rect 96250 434344 96306 434353
rect 95620 434302 96250 434330
rect 96908 434330 96936 436047
rect 96600 434302 96936 434330
rect 97000 434330 97028 437582
rect 98012 434602 98040 455398
rect 98656 438161 98684 536114
rect 98748 478174 98776 570658
rect 99392 569265 99420 571338
rect 99378 569256 99434 569265
rect 99378 569191 99434 569200
rect 100024 559020 100076 559026
rect 100024 558962 100076 558968
rect 99472 486464 99524 486470
rect 99472 486406 99524 486412
rect 98736 478168 98788 478174
rect 98736 478110 98788 478116
rect 99484 441614 99512 486406
rect 100036 442241 100064 558962
rect 100760 549364 100812 549370
rect 100760 549306 100812 549312
rect 100772 449818 100800 549306
rect 100864 518226 100892 572698
rect 100852 518220 100904 518226
rect 100852 518162 100904 518168
rect 101416 450566 101444 583879
rect 102060 576774 102088 702986
rect 105464 700330 105492 703520
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 124220 589348 124272 589354
rect 124220 589290 124272 589296
rect 123484 586560 123536 586566
rect 123484 586502 123536 586508
rect 112444 585812 112496 585818
rect 112444 585754 112496 585760
rect 121736 585812 121788 585818
rect 121736 585754 121788 585760
rect 108304 583772 108356 583778
rect 108304 583714 108356 583720
rect 104162 582584 104218 582593
rect 104162 582519 104218 582528
rect 106924 582548 106976 582554
rect 102784 580304 102836 580310
rect 102784 580246 102836 580252
rect 102048 576768 102100 576774
rect 102048 576710 102100 576716
rect 102060 576162 102088 576710
rect 102048 576156 102100 576162
rect 102048 576098 102100 576104
rect 102796 471306 102824 580246
rect 102876 487824 102928 487830
rect 102876 487766 102928 487772
rect 102140 471300 102192 471306
rect 102140 471242 102192 471248
rect 102784 471300 102836 471306
rect 102784 471242 102836 471248
rect 101404 450560 101456 450566
rect 101404 450502 101456 450508
rect 100760 449812 100812 449818
rect 100760 449754 100812 449760
rect 100772 448633 100800 449754
rect 100758 448624 100814 448633
rect 100758 448559 100814 448568
rect 100022 442232 100078 442241
rect 100022 442167 100078 442176
rect 99484 441586 99696 441614
rect 98642 438152 98698 438161
rect 98642 438087 98698 438096
rect 98012 434574 98086 434602
rect 97000 434302 97336 434330
rect 98058 434316 98086 434574
rect 99668 434330 99696 441586
rect 101218 436248 101274 436257
rect 101218 436183 101274 436192
rect 100390 434344 100446 434353
rect 99668 434302 100390 434330
rect 96250 434279 96306 434288
rect 101232 434330 101260 436183
rect 102152 434330 102180 471242
rect 102888 437442 102916 487766
rect 102876 437436 102928 437442
rect 102876 437378 102928 437384
rect 102888 434330 102916 437378
rect 103888 435464 103940 435470
rect 103888 435406 103940 435412
rect 103900 434330 103928 435406
rect 101232 434302 101568 434330
rect 102152 434302 102304 434330
rect 102888 434302 103040 434330
rect 103592 434302 103928 434330
rect 100390 434279 100446 434288
rect 92846 434208 92902 434217
rect 92538 434180 92846 434194
rect 92552 434166 92846 434180
rect 92846 434143 92902 434152
rect 85854 434072 85910 434081
rect 104176 434042 104204 582519
rect 106924 582490 106976 582496
rect 104256 581052 104308 581058
rect 104256 580994 104308 581000
rect 104268 474774 104296 580994
rect 105544 522436 105596 522442
rect 105544 522378 105596 522384
rect 104256 474768 104308 474774
rect 104256 474710 104308 474716
rect 104268 441561 104296 474710
rect 105556 469878 105584 522378
rect 106936 483682 106964 582490
rect 106924 483676 106976 483682
rect 106924 483618 106976 483624
rect 105544 469872 105596 469878
rect 105544 469814 105596 469820
rect 105556 469266 105584 469814
rect 104900 469260 104952 469266
rect 104900 469202 104952 469208
rect 105544 469260 105596 469266
rect 105544 469202 105596 469208
rect 104912 441614 104940 469202
rect 106924 447908 106976 447914
rect 106924 447850 106976 447856
rect 104912 441586 105400 441614
rect 104254 441552 104310 441561
rect 104254 441487 104310 441496
rect 104268 434602 104296 441487
rect 104440 436756 104492 436762
rect 104440 436698 104492 436704
rect 104452 435470 104480 436698
rect 104440 435464 104492 435470
rect 104440 435406 104492 435412
rect 104898 434616 104954 434625
rect 104268 434574 104342 434602
rect 104314 434316 104342 434574
rect 104898 434551 104954 434560
rect 104912 434330 104940 434551
rect 105372 434330 105400 441586
rect 106936 437345 106964 447850
rect 107660 443828 107712 443834
rect 107660 443770 107712 443776
rect 106922 437336 106978 437345
rect 106922 437271 106978 437280
rect 106936 434330 106964 437271
rect 104912 434302 105064 434330
rect 105372 434302 105800 434330
rect 106352 434302 106964 434330
rect 107672 434330 107700 443770
rect 108316 436150 108344 583714
rect 109684 569968 109736 569974
rect 109684 569910 109736 569916
rect 108396 543788 108448 543794
rect 108396 543730 108448 543736
rect 108408 443834 108436 543730
rect 109696 463593 109724 569910
rect 111064 567860 111116 567866
rect 111064 567802 111116 567808
rect 111076 478922 111104 567802
rect 111156 533384 111208 533390
rect 111156 533326 111208 533332
rect 110420 478916 110472 478922
rect 110420 478858 110472 478864
rect 111064 478916 111116 478922
rect 111064 478858 111116 478864
rect 109776 476128 109828 476134
rect 109776 476070 109828 476076
rect 109682 463584 109738 463593
rect 109682 463519 109738 463528
rect 109040 460896 109092 460902
rect 109040 460838 109092 460844
rect 109052 460222 109080 460838
rect 109788 460222 109816 476070
rect 110326 463584 110382 463593
rect 110326 463519 110382 463528
rect 110340 462369 110368 463519
rect 110326 462360 110382 462369
rect 110326 462295 110382 462304
rect 109040 460216 109092 460222
rect 109040 460158 109092 460164
rect 109776 460216 109828 460222
rect 109776 460158 109828 460164
rect 108396 443828 108448 443834
rect 108396 443770 108448 443776
rect 109052 441614 109080 460158
rect 110340 442377 110368 462295
rect 110326 442368 110382 442377
rect 110326 442303 110382 442312
rect 110432 441614 110460 478858
rect 111168 468518 111196 533326
rect 111156 468512 111208 468518
rect 111156 468454 111208 468460
rect 111708 458244 111760 458250
rect 111708 458186 111760 458192
rect 111720 455394 111748 458186
rect 111708 455388 111760 455394
rect 111708 455330 111760 455336
rect 112456 447914 112484 585754
rect 121748 585206 121776 585754
rect 121460 585200 121512 585206
rect 121460 585142 121512 585148
rect 121736 585200 121788 585206
rect 121736 585142 121788 585148
rect 119342 583808 119398 583817
rect 119342 583743 119398 583752
rect 113180 561740 113232 561746
rect 113180 561682 113232 561688
rect 112536 552084 112588 552090
rect 112536 552026 112588 552032
rect 112548 466478 112576 552026
rect 112536 466472 112588 466478
rect 112536 466414 112588 466420
rect 112444 447908 112496 447914
rect 112444 447850 112496 447856
rect 112548 444378 112576 466414
rect 112720 455388 112772 455394
rect 112720 455330 112772 455336
rect 111892 444372 111944 444378
rect 111892 444314 111944 444320
rect 112536 444372 112588 444378
rect 112536 444314 112588 444320
rect 111904 443018 111932 444314
rect 111892 443012 111944 443018
rect 111892 442954 111944 442960
rect 111904 441614 111932 442954
rect 109052 441586 109448 441614
rect 110432 441586 110920 441614
rect 111904 441586 112208 441614
rect 108304 436144 108356 436150
rect 108304 436086 108356 436092
rect 108316 434330 108344 436086
rect 109420 434330 109448 441586
rect 110786 437064 110842 437073
rect 110786 436999 110842 437008
rect 110800 434330 110828 436999
rect 107672 434302 107824 434330
rect 108316 434302 108560 434330
rect 109420 434302 109848 434330
rect 110584 434302 110828 434330
rect 110892 434330 110920 441586
rect 112180 434330 112208 441586
rect 110892 434302 111320 434330
rect 112180 434302 112608 434330
rect 85854 434007 85910 434016
rect 104164 434036 104216 434042
rect 85868 433922 85896 434007
rect 104164 433978 104216 433984
rect 85560 433894 85896 433922
rect 97722 433936 97778 433945
rect 97722 433871 97778 433880
rect 101126 433936 101182 433945
rect 101126 433871 101182 433880
rect 105358 433936 105414 433945
rect 105358 433871 105414 433880
rect 110142 433936 110198 433945
rect 110142 433871 110198 433880
rect 77170 433772 77294 433786
rect 77170 433758 77280 433772
rect 77114 433735 77170 433744
rect 68376 433696 68428 433702
rect 68376 433638 68428 433644
rect 71136 433696 71188 433702
rect 97736 433673 97764 433871
rect 101140 433673 101168 433871
rect 105372 433673 105400 433871
rect 110156 433673 110184 433871
rect 112352 433696 112404 433702
rect 71136 433638 71188 433644
rect 75458 433664 75514 433673
rect 68388 431905 68416 433638
rect 77482 433664 77538 433673
rect 75514 433622 75808 433650
rect 75458 433599 75514 433608
rect 87234 433664 87290 433673
rect 77538 433622 77832 433650
rect 77482 433599 77538 433608
rect 87970 433664 88026 433673
rect 87290 433622 87584 433650
rect 87234 433599 87290 433608
rect 89626 433664 89682 433673
rect 88026 433622 88320 433650
rect 87970 433599 88026 433608
rect 90086 433664 90142 433673
rect 89682 433622 89792 433650
rect 89626 433599 89682 433608
rect 91282 433664 91338 433673
rect 90142 433622 90344 433650
rect 91080 433622 91282 433650
rect 90086 433599 90142 433608
rect 91282 433599 91338 433608
rect 91558 433664 91614 433673
rect 92938 433664 92994 433673
rect 91614 433622 91816 433650
rect 91558 433599 91614 433608
rect 97722 433664 97778 433673
rect 92994 433622 93288 433650
rect 92938 433599 92994 433608
rect 97722 433599 97778 433608
rect 98366 433664 98422 433673
rect 99194 433664 99250 433673
rect 98422 433622 98808 433650
rect 98366 433599 98422 433608
rect 100666 433664 100722 433673
rect 99250 433622 99544 433650
rect 99194 433599 99250 433608
rect 101126 433664 101182 433673
rect 100722 433622 100832 433650
rect 100666 433599 100722 433608
rect 101126 433599 101182 433608
rect 105358 433664 105414 433673
rect 105358 433599 105414 433608
rect 106738 433664 106794 433673
rect 109038 433664 109094 433673
rect 106794 433622 107088 433650
rect 106738 433599 106794 433608
rect 110142 433664 110198 433673
rect 109094 433622 109296 433650
rect 109038 433599 109094 433608
rect 112056 433644 112352 433650
rect 112056 433638 112404 433644
rect 112056 433622 112392 433638
rect 110142 433599 110198 433608
rect 68652 433288 68704 433294
rect 68652 433230 68704 433236
rect 68664 433129 68692 433230
rect 68650 433120 68706 433129
rect 68650 433055 68706 433064
rect 68374 431896 68430 431905
rect 68374 431831 68430 431840
rect 112732 429865 112760 455330
rect 112718 429856 112774 429865
rect 112718 429791 112774 429800
rect 68284 428392 68336 428398
rect 68284 428334 68336 428340
rect 112718 418432 112774 418441
rect 112718 418367 112774 418376
rect 112732 418130 112760 418367
rect 112720 418124 112772 418130
rect 112720 418066 112772 418072
rect 70398 390960 70454 390969
rect 71686 390960 71742 390969
rect 71576 390918 71686 390946
rect 70398 390895 70454 390904
rect 71686 390895 71742 390904
rect 73986 390960 74042 390969
rect 111982 390960 112038 390969
rect 74042 390918 74488 390946
rect 73986 390895 74042 390904
rect 68652 390584 68704 390590
rect 68704 390532 68816 390538
rect 68652 390526 68816 390532
rect 68664 390510 68816 390526
rect 69368 390374 69704 390402
rect 69110 390144 69166 390153
rect 69110 390079 69166 390088
rect 69124 389201 69152 390079
rect 69110 389192 69166 389201
rect 69676 389162 69704 390374
rect 70090 390153 70118 390388
rect 70076 390144 70132 390153
rect 70076 390079 70132 390088
rect 69110 389127 69166 389136
rect 69664 389156 69716 389162
rect 68834 303648 68890 303657
rect 68834 303583 68890 303592
rect 68652 285796 68704 285802
rect 68652 285738 68704 285744
rect 68006 282976 68062 282985
rect 68006 282911 68062 282920
rect 68558 276040 68614 276049
rect 68558 275975 68614 275984
rect 68190 258768 68246 258777
rect 68190 258703 68246 258712
rect 68204 257990 68232 258703
rect 68192 257984 68244 257990
rect 68192 257926 68244 257932
rect 67822 249520 67878 249529
rect 67822 249455 67878 249464
rect 67732 242548 67784 242554
rect 67732 242490 67784 242496
rect 67744 238754 67772 242490
rect 67836 241398 67864 249455
rect 68572 241806 68600 275975
rect 68560 241800 68612 241806
rect 68560 241742 68612 241748
rect 67824 241392 67876 241398
rect 67824 241334 67876 241340
rect 68572 240145 68600 241742
rect 68664 240825 68692 285738
rect 68848 282946 68876 303583
rect 69124 283257 69152 389127
rect 69664 389098 69716 389104
rect 69294 316160 69350 316169
rect 69294 316095 69350 316104
rect 69202 284336 69258 284345
rect 69202 284271 69258 284280
rect 69110 283248 69166 283257
rect 69110 283183 69166 283192
rect 69216 283098 69244 284271
rect 69308 283529 69336 316095
rect 70412 285705 70440 390895
rect 73712 390584 73764 390590
rect 73712 390526 73764 390532
rect 70840 390374 71176 390402
rect 72128 390374 72464 390402
rect 71148 387870 71176 390374
rect 72436 389065 72464 390374
rect 72528 390374 72864 390402
rect 73172 390374 73600 390402
rect 72528 389094 72556 390374
rect 72516 389088 72568 389094
rect 72422 389056 72478 389065
rect 72516 389030 72568 389036
rect 73066 389056 73122 389065
rect 72422 388991 72478 389000
rect 71136 387864 71188 387870
rect 71136 387806 71188 387812
rect 71688 387864 71740 387870
rect 71688 387806 71740 387812
rect 71700 363662 71728 387806
rect 72528 380905 72556 389030
rect 73066 388991 73122 389000
rect 73080 383625 73108 388991
rect 73066 383616 73122 383625
rect 73066 383551 73122 383560
rect 72514 380896 72570 380905
rect 72514 380831 72570 380840
rect 73172 380186 73200 390374
rect 73724 389162 73752 390526
rect 73712 389156 73764 389162
rect 73712 389098 73764 389104
rect 74460 388793 74488 390918
rect 111982 390895 112038 390904
rect 91282 390824 91338 390833
rect 91080 390782 91282 390810
rect 91282 390759 91338 390768
rect 107934 390688 107990 390697
rect 80440 390646 80592 390674
rect 74644 390374 75072 390402
rect 75624 390374 75776 390402
rect 74446 388784 74502 388793
rect 74446 388719 74502 388728
rect 73160 380180 73212 380186
rect 73160 380122 73212 380128
rect 72422 373280 72478 373289
rect 72422 373215 72478 373224
rect 71688 363656 71740 363662
rect 71688 363598 71740 363604
rect 71964 318096 72016 318102
rect 71964 318038 72016 318044
rect 71872 289876 71924 289882
rect 71872 289818 71924 289824
rect 70858 285832 70914 285841
rect 70858 285767 70914 285776
rect 70398 285696 70454 285705
rect 70398 285631 70454 285640
rect 70306 284880 70362 284889
rect 70306 284815 70362 284824
rect 69294 283520 69350 283529
rect 70320 283506 70348 284815
rect 70872 284442 70900 285767
rect 71320 285728 71372 285734
rect 71320 285670 71372 285676
rect 71332 284510 71360 285670
rect 71320 284504 71372 284510
rect 71320 284446 71372 284452
rect 70860 284436 70912 284442
rect 70860 284378 70912 284384
rect 69350 283478 69552 283506
rect 70104 283478 70348 283506
rect 69294 283455 69350 283464
rect 69308 283395 69336 283455
rect 70872 283370 70900 284378
rect 71332 283370 71360 284446
rect 71884 283506 71912 289818
rect 71976 283665 72004 318038
rect 72436 285734 72464 373215
rect 74644 367810 74672 390374
rect 74632 367804 74684 367810
rect 74632 367746 74684 367752
rect 75748 355366 75776 390374
rect 75932 390374 76360 390402
rect 77096 390374 77248 390402
rect 77832 390374 78168 390402
rect 78384 390374 78628 390402
rect 75826 386200 75882 386209
rect 75826 386135 75882 386144
rect 75736 355360 75788 355366
rect 75736 355302 75788 355308
rect 75840 320210 75868 386135
rect 75932 372502 75960 390374
rect 77220 386345 77248 390374
rect 78140 387870 78168 390374
rect 78600 389473 78628 390374
rect 79106 390130 79134 390388
rect 79244 390374 79856 390402
rect 79106 390102 79180 390130
rect 78586 389464 78642 389473
rect 78586 389399 78642 389408
rect 79152 389065 79180 390102
rect 79138 389056 79194 389065
rect 79138 388991 79194 389000
rect 78128 387864 78180 387870
rect 78128 387806 78180 387812
rect 78588 387864 78640 387870
rect 78588 387806 78640 387812
rect 77206 386336 77262 386345
rect 77206 386271 77262 386280
rect 77484 380248 77536 380254
rect 77484 380190 77536 380196
rect 75920 372496 75972 372502
rect 75920 372438 75972 372444
rect 75932 366382 75960 372438
rect 75920 366376 75972 366382
rect 75920 366318 75972 366324
rect 75828 320204 75880 320210
rect 75828 320146 75880 320152
rect 75182 317384 75238 317393
rect 75182 317319 75238 317328
rect 73068 301504 73120 301510
rect 73068 301446 73120 301452
rect 73080 287054 73108 301446
rect 72620 287026 73108 287054
rect 72424 285728 72476 285734
rect 72424 285670 72476 285676
rect 71962 283656 72018 283665
rect 71962 283591 72018 283600
rect 71760 283478 71912 283506
rect 70656 283342 70900 283370
rect 71208 283342 71360 283370
rect 69000 283070 69244 283098
rect 72422 282976 72478 282985
rect 68836 282940 68888 282946
rect 72312 282934 72422 282962
rect 72620 282962 72648 287026
rect 73802 286240 73858 286249
rect 73802 286175 73858 286184
rect 73710 285696 73766 285705
rect 73710 285631 73766 285640
rect 73724 283121 73752 285631
rect 73816 283506 73844 286175
rect 75196 285977 75224 317319
rect 75736 286340 75788 286346
rect 75736 286282 75788 286288
rect 74906 285968 74962 285977
rect 74906 285903 74962 285912
rect 75182 285968 75238 285977
rect 75182 285903 75238 285912
rect 74816 285728 74868 285734
rect 74816 285670 74868 285676
rect 74828 283506 74856 285670
rect 73816 283478 73968 283506
rect 74520 283478 74856 283506
rect 74920 283506 74948 285903
rect 75748 283506 75776 286282
rect 75840 285734 75868 320146
rect 75918 320104 75974 320113
rect 75918 320039 75974 320048
rect 75828 285728 75880 285734
rect 75828 285670 75880 285676
rect 75932 284986 75960 320039
rect 77392 295384 77444 295390
rect 77392 295326 77444 295332
rect 77298 292768 77354 292777
rect 77298 292703 77354 292712
rect 76010 292632 76066 292641
rect 76010 292567 76066 292576
rect 75920 284980 75972 284986
rect 75920 284922 75972 284928
rect 74920 283478 75072 283506
rect 75624 283478 75776 283506
rect 76024 283506 76052 292567
rect 76380 284980 76432 284986
rect 76380 284922 76432 284928
rect 76392 283506 76420 284922
rect 77312 283778 77340 292703
rect 77266 283750 77340 283778
rect 76024 283478 76176 283506
rect 76392 283478 76728 283506
rect 77266 283492 77294 283750
rect 77404 283506 77432 295326
rect 77496 289134 77524 380190
rect 78600 377466 78628 387806
rect 78588 377460 78640 377466
rect 78588 377402 78640 377408
rect 79244 373994 79272 390374
rect 79874 389056 79930 389065
rect 79874 388991 79930 389000
rect 80058 389056 80114 389065
rect 80058 388991 80114 389000
rect 79322 387016 79378 387025
rect 79322 386951 79378 386960
rect 78692 373966 79272 373994
rect 78586 322824 78642 322833
rect 78586 322759 78642 322768
rect 78600 296002 78628 322759
rect 78588 295996 78640 296002
rect 78588 295938 78640 295944
rect 78600 295390 78628 295938
rect 78588 295384 78640 295390
rect 78588 295326 78640 295332
rect 78692 293282 78720 373966
rect 78680 293276 78732 293282
rect 78680 293218 78732 293224
rect 77484 289128 77536 289134
rect 77484 289070 77536 289076
rect 78588 287700 78640 287706
rect 78588 287642 78640 287648
rect 78600 283506 78628 287642
rect 79232 285728 79284 285734
rect 79336 285705 79364 386951
rect 79888 382265 79916 388991
rect 79966 388376 80022 388385
rect 79966 388311 80022 388320
rect 79980 387870 80008 388311
rect 79968 387864 80020 387870
rect 79968 387806 80020 387812
rect 79874 382256 79930 382265
rect 79874 382191 79930 382200
rect 79980 354686 80008 387806
rect 79968 354680 80020 354686
rect 79968 354622 80020 354628
rect 79966 318064 80022 318073
rect 79966 317999 80022 318008
rect 79980 289814 80008 317999
rect 80072 309942 80100 388991
rect 80440 385665 80468 390646
rect 111996 390658 112024 390895
rect 107934 390623 107990 390632
rect 111984 390652 112036 390658
rect 96986 390552 97042 390561
rect 93840 390510 93992 390538
rect 80992 390374 81328 390402
rect 81544 390374 81880 390402
rect 82004 390374 82616 390402
rect 83016 390374 83352 390402
rect 83476 390374 84088 390402
rect 84212 390374 84824 390402
rect 85040 390374 85376 390402
rect 85592 390374 86112 390402
rect 80992 389065 81020 390374
rect 80978 389056 81034 389065
rect 80978 388991 81034 389000
rect 81544 387870 81572 390374
rect 81532 387864 81584 387870
rect 81532 387806 81584 387812
rect 80426 385656 80482 385665
rect 80426 385591 80482 385600
rect 82004 373994 82032 390374
rect 83016 389230 83044 390374
rect 83004 389224 83056 389230
rect 83004 389166 83056 389172
rect 83016 388385 83044 389166
rect 83002 388376 83058 388385
rect 83002 388311 83058 388320
rect 83476 387002 83504 390374
rect 82832 386974 83504 387002
rect 82084 385688 82136 385694
rect 82084 385630 82136 385636
rect 81544 373966 82032 373994
rect 81544 354006 81572 373966
rect 81532 354000 81584 354006
rect 81532 353942 81584 353948
rect 80060 309936 80112 309942
rect 80060 309878 80112 309884
rect 81346 309904 81402 309913
rect 81346 309839 81402 309848
rect 81360 292574 81388 309839
rect 81806 297528 81862 297537
rect 81806 297463 81862 297472
rect 80992 292546 81388 292574
rect 79968 289808 80020 289814
rect 79968 289750 80020 289756
rect 79980 285734 80008 289750
rect 80152 289128 80204 289134
rect 80152 289070 80204 289076
rect 79968 285728 80020 285734
rect 79232 285670 79284 285676
rect 79322 285696 79378 285705
rect 79244 283506 79272 285670
rect 79968 285670 80020 285676
rect 79322 285631 79378 285640
rect 77404 283478 77832 283506
rect 78384 283478 78628 283506
rect 78936 283478 79272 283506
rect 79336 283506 79364 285631
rect 79336 283478 79488 283506
rect 72698 283112 72754 283121
rect 73710 283112 73766 283121
rect 72754 283070 72864 283098
rect 72698 283047 72754 283056
rect 73710 283047 73766 283056
rect 76024 283014 76052 283478
rect 80164 283370 80192 289070
rect 80992 285977 81020 292546
rect 81530 286104 81586 286113
rect 81530 286039 81586 286048
rect 80978 285968 81034 285977
rect 80978 285903 81034 285912
rect 80992 283506 81020 285903
rect 81256 285864 81308 285870
rect 81256 285806 81308 285812
rect 80592 283478 81020 283506
rect 81268 283370 81296 285806
rect 80040 283342 80192 283370
rect 81144 283342 81296 283370
rect 81544 283370 81572 286039
rect 81820 283506 81848 297463
rect 82096 286113 82124 385630
rect 82832 366382 82860 386974
rect 83462 384296 83518 384305
rect 83462 384231 83518 384240
rect 82820 366376 82872 366382
rect 82820 366318 82872 366324
rect 82910 313304 82966 313313
rect 82910 313239 82966 313248
rect 82924 306374 82952 313239
rect 82924 306346 83412 306374
rect 83094 291816 83150 291825
rect 83094 291751 83150 291760
rect 82082 286104 82138 286113
rect 82082 286039 82138 286048
rect 83108 283506 83136 291751
rect 83186 286104 83242 286113
rect 83186 286039 83242 286048
rect 81820 283478 82248 283506
rect 82800 283478 83136 283506
rect 83200 283370 83228 286039
rect 83384 285716 83412 306346
rect 83476 285870 83504 384231
rect 84212 358766 84240 390374
rect 85040 378729 85068 390374
rect 85026 378720 85082 378729
rect 85026 378655 85082 378664
rect 85592 361554 85620 390374
rect 86834 390130 86862 390388
rect 87064 390374 87584 390402
rect 87800 390374 88136 390402
rect 88872 390374 89208 390402
rect 86834 390102 86908 390130
rect 86224 387864 86276 387870
rect 86224 387806 86276 387812
rect 86236 385014 86264 387806
rect 86880 387433 86908 390102
rect 86866 387424 86922 387433
rect 86866 387359 86922 387368
rect 86224 385008 86276 385014
rect 86224 384950 86276 384956
rect 86236 362846 86264 384950
rect 86224 362840 86276 362846
rect 86224 362782 86276 362788
rect 85580 361548 85632 361554
rect 85580 361490 85632 361496
rect 84200 358760 84252 358766
rect 84200 358702 84252 358708
rect 86224 322244 86276 322250
rect 86224 322186 86276 322192
rect 84200 308440 84252 308446
rect 84200 308382 84252 308388
rect 84106 293312 84162 293321
rect 84106 293247 84162 293256
rect 84120 286113 84148 293247
rect 84106 286104 84162 286113
rect 84106 286039 84162 286048
rect 83464 285864 83516 285870
rect 83464 285806 83516 285812
rect 83384 285688 83504 285716
rect 83476 283506 83504 285688
rect 84212 283506 84240 308382
rect 86236 291854 86264 322186
rect 86866 319424 86922 319433
rect 86866 319359 86922 319368
rect 86774 309768 86830 309777
rect 86774 309703 86830 309712
rect 86224 291848 86276 291854
rect 86224 291790 86276 291796
rect 86788 291242 86816 309703
rect 85856 291236 85908 291242
rect 85856 291178 85908 291184
rect 86776 291236 86828 291242
rect 86776 291178 86828 291184
rect 85304 285932 85356 285938
rect 85304 285874 85356 285880
rect 85316 283506 85344 285874
rect 85868 283506 85896 291178
rect 86682 283792 86738 283801
rect 86512 283750 86682 283778
rect 86512 283506 86540 283750
rect 86880 283778 86908 319359
rect 87064 317393 87092 390374
rect 87604 387932 87656 387938
rect 87604 387874 87656 387880
rect 87616 384946 87644 387874
rect 87800 387870 87828 390374
rect 87788 387864 87840 387870
rect 87788 387806 87840 387812
rect 89180 384946 89208 390374
rect 89272 390374 89608 390402
rect 89732 390374 90344 390402
rect 91296 390374 91632 390402
rect 92032 390374 92368 390402
rect 92492 390374 93104 390402
rect 89272 386374 89300 390374
rect 89260 386368 89312 386374
rect 89260 386310 89312 386316
rect 87604 384940 87656 384946
rect 87604 384882 87656 384888
rect 89168 384940 89220 384946
rect 89168 384882 89220 384888
rect 87616 375358 87644 384882
rect 88982 382936 89038 382945
rect 88982 382871 89038 382880
rect 87604 375352 87656 375358
rect 87604 375294 87656 375300
rect 88248 375352 88300 375358
rect 88248 375294 88300 375300
rect 88260 342310 88288 375294
rect 88996 345098 89024 382871
rect 89272 373994 89300 386310
rect 89626 385656 89682 385665
rect 89626 385591 89682 385600
rect 89088 373966 89300 373994
rect 89088 367878 89116 373966
rect 89076 367872 89128 367878
rect 89076 367814 89128 367820
rect 88984 345092 89036 345098
rect 88984 345034 89036 345040
rect 88248 342304 88300 342310
rect 88248 342246 88300 342252
rect 88154 318064 88210 318073
rect 88154 317999 88210 318008
rect 87050 317384 87106 317393
rect 87050 317319 87106 317328
rect 87604 316668 87656 316674
rect 87604 316610 87656 316616
rect 86960 294704 87012 294710
rect 86960 294646 87012 294652
rect 86738 283750 86908 283778
rect 86682 283727 86738 283736
rect 86696 283667 86724 283727
rect 83476 283478 83904 283506
rect 84212 283478 84456 283506
rect 85008 283478 85344 283506
rect 85560 283478 85896 283506
rect 86112 283478 86540 283506
rect 86972 283506 87000 294646
rect 87616 290494 87644 316610
rect 87696 302320 87748 302326
rect 87696 302262 87748 302268
rect 87604 290488 87656 290494
rect 87604 290430 87656 290436
rect 87708 285938 87736 302262
rect 88168 287094 88196 317999
rect 88260 316674 88288 342246
rect 88996 318102 89024 345034
rect 88984 318096 89036 318102
rect 88984 318038 89036 318044
rect 88248 316668 88300 316674
rect 88248 316610 88300 316616
rect 88260 316062 88288 316610
rect 88248 316056 88300 316062
rect 88248 315998 88300 316004
rect 88430 304192 88486 304201
rect 88430 304127 88486 304136
rect 87880 287088 87932 287094
rect 87880 287030 87932 287036
rect 88156 287088 88208 287094
rect 88156 287030 88208 287036
rect 87696 285932 87748 285938
rect 87696 285874 87748 285880
rect 87892 283506 87920 287030
rect 88294 283756 88346 283762
rect 88294 283698 88346 283704
rect 88306 283506 88334 283698
rect 86972 283478 87216 283506
rect 87768 283478 87920 283506
rect 88168 283492 88334 283506
rect 88444 283506 88472 304127
rect 89534 293176 89590 293185
rect 89534 293111 89590 293120
rect 89548 283762 89576 293111
rect 89536 283756 89588 283762
rect 89536 283698 89588 283704
rect 89534 283520 89590 283529
rect 88168 283478 88320 283492
rect 88444 283478 88872 283506
rect 89424 283478 89534 283506
rect 81544 283342 81696 283370
rect 83200 283342 83504 283370
rect 83476 283257 83504 283342
rect 88168 283257 88196 283478
rect 89640 283506 89668 385591
rect 89732 289785 89760 390374
rect 91098 387832 91154 387841
rect 91098 387767 91154 387776
rect 91112 385694 91140 387767
rect 91100 385688 91152 385694
rect 91100 385630 91152 385636
rect 91006 383752 91062 383761
rect 91006 383687 91062 383696
rect 89718 289776 89774 289785
rect 89718 289711 89774 289720
rect 90916 286272 90968 286278
rect 90916 286214 90968 286220
rect 90270 286104 90326 286113
rect 90270 286039 90326 286048
rect 90086 283520 90142 283529
rect 89590 283478 89668 283506
rect 89976 283478 90086 283506
rect 89534 283455 89590 283464
rect 90284 283506 90312 286039
rect 90822 285696 90878 285705
rect 90822 285631 90878 285640
rect 90836 283506 90864 285631
rect 90142 283478 90312 283506
rect 90528 283478 90864 283506
rect 90086 283455 90142 283464
rect 89548 283395 89576 283455
rect 90100 283395 90128 283455
rect 90928 283370 90956 286214
rect 91020 286113 91048 383687
rect 91192 297424 91244 297430
rect 91192 297366 91244 297372
rect 91006 286104 91062 286113
rect 91006 286039 91062 286048
rect 91204 283506 91232 297366
rect 91296 291145 91324 390374
rect 92032 387938 92060 390374
rect 92020 387932 92072 387938
rect 92020 387874 92072 387880
rect 92492 376650 92520 390374
rect 93964 387802 93992 390510
rect 101034 390552 101090 390561
rect 97042 390510 97488 390538
rect 96986 390487 97042 390496
rect 94056 390374 94392 390402
rect 93952 387796 94004 387802
rect 93952 387738 94004 387744
rect 92480 376644 92532 376650
rect 92480 376586 92532 376592
rect 94056 370530 94084 390374
rect 95114 390130 95142 390388
rect 95252 390374 95864 390402
rect 96600 390374 96936 390402
rect 95114 390102 95188 390130
rect 94504 387796 94556 387802
rect 94504 387738 94556 387744
rect 94044 370524 94096 370530
rect 94044 370466 94096 370472
rect 94516 359582 94544 387738
rect 94504 359576 94556 359582
rect 94504 359518 94556 359524
rect 95160 351898 95188 390102
rect 95148 351892 95200 351898
rect 95148 351834 95200 351840
rect 93766 329080 93822 329089
rect 93766 329015 93822 329024
rect 92848 298784 92900 298790
rect 92848 298726 92900 298732
rect 91282 291136 91338 291145
rect 91282 291071 91338 291080
rect 92710 283756 92762 283762
rect 92710 283698 92762 283704
rect 91204 283478 91632 283506
rect 92722 283492 92750 283698
rect 92860 283506 92888 298726
rect 93780 293962 93808 329015
rect 95146 319424 95202 319433
rect 95146 319359 95202 319368
rect 94502 316160 94558 316169
rect 94502 316095 94558 316104
rect 93768 293956 93820 293962
rect 93768 293898 93820 293904
rect 93780 283762 93808 293898
rect 94516 286278 94544 316095
rect 95160 292574 95188 319359
rect 94792 292546 95188 292574
rect 94504 286272 94556 286278
rect 94504 286214 94556 286220
rect 93858 285696 93914 285705
rect 93858 285631 93914 285640
rect 93872 285025 93900 285631
rect 93858 285016 93914 285025
rect 93858 284951 93914 284960
rect 93768 283756 93820 283762
rect 93768 283698 93820 283704
rect 94042 283520 94098 283529
rect 92860 283478 93288 283506
rect 94792 283506 94820 292546
rect 95148 291236 95200 291242
rect 95148 291178 95200 291184
rect 95160 283506 95188 291178
rect 95252 288561 95280 390374
rect 96908 388929 96936 390374
rect 97460 389065 97488 390510
rect 100956 390510 101034 390538
rect 99654 390416 99710 390425
rect 97552 390374 97888 390402
rect 98624 390374 98960 390402
rect 99360 390374 99654 390402
rect 97446 389056 97502 389065
rect 97446 388991 97502 389000
rect 96894 388920 96950 388929
rect 96894 388855 96950 388864
rect 97552 373994 97580 390374
rect 97906 389056 97962 389065
rect 97906 388991 97962 389000
rect 97920 382974 97948 388991
rect 98932 387569 98960 390374
rect 100956 390402 100984 390510
rect 101034 390487 101090 390496
rect 105266 390416 105322 390425
rect 100096 390374 100432 390402
rect 100832 390374 100984 390402
rect 99654 390351 99710 390360
rect 98918 387560 98974 387569
rect 98918 387495 98974 387504
rect 99668 386374 99696 390351
rect 100404 387802 100432 390374
rect 100392 387796 100444 387802
rect 100392 387738 100444 387744
rect 99656 386368 99708 386374
rect 99656 386310 99708 386316
rect 100852 386368 100904 386374
rect 100852 386310 100904 386316
rect 100864 385801 100892 386310
rect 100850 385792 100906 385801
rect 100850 385727 100906 385736
rect 100956 385014 100984 390374
rect 101048 390374 101384 390402
rect 100944 385008 100996 385014
rect 100944 384950 100996 384956
rect 97908 382968 97960 382974
rect 97908 382910 97960 382916
rect 101048 382226 101076 390374
rect 102106 390130 102134 390388
rect 102856 390374 103192 390402
rect 102106 390102 102180 390130
rect 101956 385688 102008 385694
rect 101956 385630 102008 385636
rect 101036 382220 101088 382226
rect 101036 382162 101088 382168
rect 101404 381540 101456 381546
rect 101404 381482 101456 381488
rect 96632 373966 97580 373994
rect 96526 309768 96582 309777
rect 96526 309703 96582 309712
rect 96540 292574 96568 309703
rect 96448 292546 96568 292574
rect 95238 288552 95294 288561
rect 95238 288487 95294 288496
rect 95792 287020 95844 287026
rect 95792 286962 95844 286968
rect 95804 283506 95832 286962
rect 96448 285705 96476 292546
rect 96632 289921 96660 373966
rect 100576 373312 100628 373318
rect 100576 373254 100628 373260
rect 97262 325000 97318 325009
rect 97262 324935 97318 324944
rect 96712 293276 96764 293282
rect 96712 293218 96764 293224
rect 96618 289912 96674 289921
rect 96618 289847 96674 289856
rect 96434 285696 96490 285705
rect 96434 285631 96490 285640
rect 96448 283506 96476 285631
rect 94098 283478 94820 283506
rect 94944 283478 95188 283506
rect 95496 283478 95832 283506
rect 96048 283478 96476 283506
rect 96724 283506 96752 293218
rect 97276 287745 97304 324935
rect 98000 319456 98052 319462
rect 98000 319398 98052 319404
rect 97908 304360 97960 304366
rect 97908 304302 97960 304308
rect 97920 288454 97948 304302
rect 97540 288448 97592 288454
rect 97540 288390 97592 288396
rect 97908 288448 97960 288454
rect 97908 288390 97960 288396
rect 97262 287736 97318 287745
rect 97262 287671 97318 287680
rect 97552 287026 97580 288390
rect 97540 287020 97592 287026
rect 97540 286962 97592 286968
rect 97262 286376 97318 286385
rect 97262 286311 97318 286320
rect 96724 283478 97152 283506
rect 94042 283455 94098 283464
rect 97276 283422 97304 286311
rect 96896 283416 96948 283422
rect 90928 283342 91080 283370
rect 96600 283364 96896 283370
rect 96600 283358 96948 283364
rect 97264 283416 97316 283422
rect 97264 283358 97316 283364
rect 96600 283342 96936 283358
rect 83462 283248 83518 283257
rect 83462 283183 83518 283192
rect 88154 283248 88210 283257
rect 92386 283248 92442 283257
rect 92184 283206 92386 283234
rect 88154 283183 88210 283192
rect 92386 283183 92442 283192
rect 86664 283082 86908 283098
rect 86664 283076 86920 283082
rect 86664 283070 86868 283076
rect 86868 283018 86920 283024
rect 76012 283008 76064 283014
rect 73526 282976 73582 282985
rect 72478 282934 72648 282962
rect 73416 282934 73526 282962
rect 72422 282911 72478 282920
rect 94136 283008 94188 283014
rect 76012 282950 76064 282956
rect 93840 282956 94136 282962
rect 97906 282976 97962 282985
rect 93840 282950 94188 282956
rect 93840 282934 94176 282950
rect 97704 282934 97906 282962
rect 73526 282911 73582 282920
rect 97906 282911 97962 282920
rect 68836 282882 68888 282888
rect 68848 281217 68876 282882
rect 98012 282690 98040 319398
rect 100022 297528 100078 297537
rect 100022 297463 100078 297472
rect 98460 290556 98512 290562
rect 98460 290498 98512 290504
rect 98472 283506 98500 290498
rect 98734 284880 98790 284889
rect 98734 284815 98790 284824
rect 98256 283478 98500 283506
rect 98380 282798 98624 282826
rect 98380 282690 98408 282798
rect 98012 282662 98408 282690
rect 68834 281208 68890 281217
rect 68834 281143 68890 281152
rect 68848 280226 68876 281143
rect 68836 280220 68888 280226
rect 68836 280162 68888 280168
rect 98380 277394 98408 282662
rect 98104 277366 98408 277394
rect 98000 243568 98052 243574
rect 98000 243510 98052 243516
rect 68790 242548 68842 242554
rect 68790 242490 68842 242496
rect 68802 242284 68830 242490
rect 69388 241800 69440 241806
rect 70950 241768 71006 241777
rect 69440 241748 69736 241754
rect 69388 241742 69736 241748
rect 69400 241726 69736 241742
rect 70840 241726 70950 241754
rect 83830 241768 83886 241777
rect 83536 241726 83830 241754
rect 70950 241703 71006 241712
rect 83830 241703 83886 241712
rect 86590 241768 86646 241777
rect 90362 241768 90418 241777
rect 86646 241726 86848 241754
rect 90160 241726 90362 241754
rect 86590 241703 86646 241712
rect 90362 241703 90418 241712
rect 91558 241768 91614 241777
rect 95882 241768 95938 241777
rect 91614 241726 92244 241754
rect 91558 241703 91614 241712
rect 85854 241632 85910 241641
rect 69184 241590 69520 241618
rect 68926 241496 68982 241505
rect 68926 241431 68982 241440
rect 68650 240816 68706 240825
rect 68650 240751 68706 240760
rect 68558 240136 68614 240145
rect 68558 240071 68614 240080
rect 67652 238726 67772 238754
rect 67546 129840 67602 129849
rect 67546 129775 67602 129784
rect 67546 128888 67602 128897
rect 67546 128823 67602 128832
rect 67560 125225 67588 128823
rect 67546 125216 67602 125225
rect 67546 125151 67602 125160
rect 67546 109440 67602 109449
rect 67546 109375 67602 109384
rect 67454 97200 67510 97209
rect 67454 97135 67510 97144
rect 67468 92041 67496 97135
rect 67560 95198 67588 109375
rect 67548 95192 67600 95198
rect 67548 95134 67600 95140
rect 67548 93832 67600 93838
rect 67548 93774 67600 93780
rect 67454 92032 67510 92041
rect 67454 91967 67510 91976
rect 67560 89690 67588 93774
rect 67652 92886 67680 238726
rect 68940 231169 68968 241431
rect 69492 239426 69520 241590
rect 69860 241590 70288 241618
rect 71392 241590 71452 241618
rect 71944 241590 72280 241618
rect 72496 241590 72832 241618
rect 69480 239420 69532 239426
rect 69480 239362 69532 239368
rect 69860 238754 69888 241590
rect 71424 240145 71452 241590
rect 71410 240136 71466 240145
rect 70400 240100 70452 240106
rect 71410 240071 71466 240080
rect 71870 240136 71926 240145
rect 71870 240071 71926 240080
rect 70400 240042 70452 240048
rect 70306 239184 70362 239193
rect 70306 239119 70362 239128
rect 69308 238726 69888 238754
rect 68926 231160 68982 231169
rect 68926 231095 68982 231104
rect 67730 165608 67786 165617
rect 67730 165543 67786 165552
rect 67744 164393 67772 165543
rect 67730 164384 67786 164393
rect 67730 164319 67786 164328
rect 67744 132841 67772 164319
rect 69020 142792 69072 142798
rect 69020 142734 69072 142740
rect 67916 138032 67968 138038
rect 67822 138000 67878 138009
rect 67916 137974 67968 137980
rect 67822 137935 67878 137944
rect 67730 132832 67786 132841
rect 67730 132767 67786 132776
rect 67730 129024 67786 129033
rect 67730 128959 67786 128968
rect 67640 92880 67692 92886
rect 67640 92822 67692 92828
rect 67548 89684 67600 89690
rect 67548 89626 67600 89632
rect 67364 86896 67416 86902
rect 67364 86838 67416 86844
rect 67272 60716 67324 60722
rect 67272 60658 67324 60664
rect 67652 59362 67680 92822
rect 67640 59356 67692 59362
rect 67640 59298 67692 59304
rect 65616 46232 65668 46238
rect 65616 46174 65668 46180
rect 67548 46232 67600 46238
rect 67548 46174 67600 46180
rect 66168 24132 66220 24138
rect 66168 24074 66220 24080
rect 65444 6886 65564 6914
rect 64328 3528 64380 3534
rect 61856 3454 62068 3482
rect 64328 3470 64380 3476
rect 64788 3528 64840 3534
rect 64788 3470 64840 3476
rect 62040 480 62068 3454
rect 63224 3460 63276 3466
rect 63224 3402 63276 3408
rect 63236 480 63264 3402
rect 64340 480 64368 3470
rect 65444 2106 65472 6886
rect 66180 3534 66208 24074
rect 67560 3534 67588 46174
rect 67744 36582 67772 128959
rect 67836 112441 67864 137935
rect 67928 128217 67956 137974
rect 69032 134994 69060 142734
rect 69308 140865 69336 238726
rect 70320 215257 70348 239119
rect 70306 215248 70362 215257
rect 70306 215183 70362 215192
rect 70320 214849 70348 215183
rect 69662 214840 69718 214849
rect 69662 214775 69718 214784
rect 70306 214840 70362 214849
rect 70306 214775 70362 214784
rect 69294 140856 69350 140865
rect 69294 140791 69350 140800
rect 69676 135930 69704 214775
rect 70216 138168 70268 138174
rect 70216 138110 70268 138116
rect 69846 137456 69902 137465
rect 69846 137391 69902 137400
rect 69664 135924 69716 135930
rect 69664 135866 69716 135872
rect 68986 134966 69060 134994
rect 68986 134708 69014 134966
rect 69860 134722 69888 137391
rect 70228 134722 70256 138110
rect 70412 138106 70440 240042
rect 70490 153096 70546 153105
rect 70490 153031 70546 153040
rect 70400 138100 70452 138106
rect 70400 138042 70452 138048
rect 70308 135924 70360 135930
rect 70308 135866 70360 135872
rect 70320 135017 70348 135866
rect 70306 135008 70362 135017
rect 70306 134943 70362 134952
rect 69552 134694 69888 134722
rect 70104 134694 70256 134722
rect 70504 134722 70532 153031
rect 71778 146976 71834 146985
rect 71778 146911 71834 146920
rect 70582 143440 70638 143449
rect 70582 143375 70638 143384
rect 70596 142798 70624 143375
rect 70584 142792 70636 142798
rect 70584 142734 70636 142740
rect 71134 140856 71190 140865
rect 71134 140791 71190 140800
rect 71148 134722 71176 140791
rect 71228 138100 71280 138106
rect 71228 138042 71280 138048
rect 70504 134694 70656 134722
rect 71024 134694 71176 134722
rect 71240 134722 71268 138042
rect 71792 134722 71820 146911
rect 71884 138174 71912 240071
rect 72252 240009 72280 241590
rect 72238 240000 72294 240009
rect 72238 239935 72294 239944
rect 72804 239329 72832 241590
rect 72896 241590 73048 241618
rect 73540 241590 73600 241618
rect 73816 241590 74152 241618
rect 74644 241590 74704 241618
rect 74828 241590 75256 241618
rect 75472 241590 75808 241618
rect 75932 241590 76360 241618
rect 76576 241590 76912 241618
rect 72896 239465 72924 241590
rect 73540 241466 73568 241590
rect 73528 241460 73580 241466
rect 73528 241402 73580 241408
rect 72974 240136 73030 240145
rect 72974 240071 73030 240080
rect 72882 239456 72938 239465
rect 72882 239391 72938 239400
rect 72790 239320 72846 239329
rect 72790 239255 72846 239264
rect 72988 236706 73016 240071
rect 73540 239873 73568 241402
rect 73526 239864 73582 239873
rect 73526 239799 73582 239808
rect 73816 238754 73844 241590
rect 74540 240168 74592 240174
rect 74354 240136 74410 240145
rect 74540 240110 74592 240116
rect 74354 240071 74410 240080
rect 73172 238726 73844 238754
rect 72976 236700 73028 236706
rect 72976 236642 73028 236648
rect 73172 232558 73200 238726
rect 74368 238542 74396 240071
rect 74356 238536 74408 238542
rect 74356 238478 74408 238484
rect 73160 232552 73212 232558
rect 73160 232494 73212 232500
rect 73436 231124 73488 231130
rect 73436 231066 73488 231072
rect 73068 149184 73120 149190
rect 73068 149126 73120 149132
rect 72330 138680 72386 138689
rect 72330 138615 72386 138624
rect 71872 138168 71924 138174
rect 71872 138110 71924 138116
rect 72344 134722 72372 138615
rect 73080 137902 73108 149126
rect 73342 147792 73398 147801
rect 73342 147727 73398 147736
rect 73356 138106 73384 147727
rect 73344 138100 73396 138106
rect 73344 138042 73396 138048
rect 73068 137896 73120 137902
rect 73068 137838 73120 137844
rect 73080 136762 73108 137838
rect 73080 136734 73200 136762
rect 73172 134994 73200 136734
rect 73172 134966 73246 134994
rect 71240 134694 71576 134722
rect 71792 134694 72128 134722
rect 72344 134694 72680 134722
rect 73218 134708 73246 134966
rect 73448 134722 73476 231066
rect 74552 199510 74580 240110
rect 74644 238066 74672 241590
rect 74632 238060 74684 238066
rect 74632 238002 74684 238008
rect 74828 220153 74856 241590
rect 75472 240174 75500 241590
rect 75460 240168 75512 240174
rect 75460 240110 75512 240116
rect 75932 238513 75960 241590
rect 76104 240100 76156 240106
rect 76104 240042 76156 240048
rect 75918 238504 75974 238513
rect 75918 238439 75974 238448
rect 76116 237386 76144 240042
rect 76576 239193 76604 241590
rect 77450 241534 77478 241604
rect 77588 241590 78016 241618
rect 78140 241590 78568 241618
rect 78784 241590 79120 241618
rect 79336 241590 79672 241618
rect 80164 241590 80224 241618
rect 80348 241590 80776 241618
rect 80992 241590 81328 241618
rect 81880 241590 82216 241618
rect 77438 241528 77490 241534
rect 77438 241470 77490 241476
rect 77450 241346 77478 241470
rect 77404 241318 77478 241346
rect 76562 239184 76618 239193
rect 76562 239119 76618 239128
rect 76656 238536 76708 238542
rect 76656 238478 76708 238484
rect 76104 237380 76156 237386
rect 76104 237322 76156 237328
rect 76116 236026 76144 237322
rect 76104 236020 76156 236026
rect 76104 235962 76156 235968
rect 76564 233912 76616 233918
rect 76564 233854 76616 233860
rect 76104 228404 76156 228410
rect 76104 228346 76156 228352
rect 74814 220144 74870 220153
rect 74814 220079 74870 220088
rect 74828 219434 74856 220079
rect 74828 219406 75224 219434
rect 74540 199504 74592 199510
rect 74540 199446 74592 199452
rect 74538 162072 74594 162081
rect 74538 162007 74594 162016
rect 73804 138100 73856 138106
rect 73804 138042 73856 138048
rect 73816 134722 73844 138042
rect 74552 134722 74580 162007
rect 75196 153882 75224 219406
rect 75920 169788 75972 169794
rect 75920 169730 75972 169736
rect 75276 158024 75328 158030
rect 75276 157966 75328 157972
rect 75184 153876 75236 153882
rect 75184 153818 75236 153824
rect 74814 145616 74870 145625
rect 74814 145551 74870 145560
rect 74828 134722 74856 145551
rect 75288 138014 75316 157966
rect 75932 151814 75960 169730
rect 75932 151786 76052 151814
rect 75918 140992 75974 141001
rect 75918 140927 75974 140936
rect 75288 137986 75408 138014
rect 75380 136785 75408 137986
rect 75366 136776 75422 136785
rect 75366 136711 75422 136720
rect 75380 134722 75408 136711
rect 75932 134722 75960 140927
rect 76024 134858 76052 151786
rect 76116 138009 76144 228346
rect 76102 138000 76158 138009
rect 76102 137935 76158 137944
rect 76576 136746 76604 233854
rect 76668 170406 76696 238478
rect 76748 236020 76800 236026
rect 76748 235962 76800 235968
rect 76760 224262 76788 235962
rect 77404 233918 77432 241318
rect 77588 240394 77616 241590
rect 78140 240938 78168 241590
rect 77496 240366 77616 240394
rect 77680 240910 78168 240938
rect 77496 240106 77524 240366
rect 77484 240100 77536 240106
rect 77484 240042 77536 240048
rect 77680 238754 77708 240910
rect 77942 240816 77998 240825
rect 77942 240751 77998 240760
rect 77588 238726 77708 238754
rect 77588 238377 77616 238726
rect 77574 238368 77630 238377
rect 77574 238303 77630 238312
rect 77392 233912 77444 233918
rect 77392 233854 77444 233860
rect 77300 232552 77352 232558
rect 77300 232494 77352 232500
rect 77208 228404 77260 228410
rect 77208 228346 77260 228352
rect 77220 227798 77248 228346
rect 77208 227792 77260 227798
rect 77208 227734 77260 227740
rect 76748 224256 76800 224262
rect 76748 224198 76800 224204
rect 76656 170400 76708 170406
rect 76656 170342 76708 170348
rect 76668 169794 76696 170342
rect 76656 169788 76708 169794
rect 76656 169730 76708 169736
rect 77312 141438 77340 232494
rect 77588 229770 77616 238303
rect 77576 229764 77628 229770
rect 77576 229706 77628 229712
rect 77956 151814 77984 240751
rect 78680 240168 78732 240174
rect 78680 240110 78732 240116
rect 78692 232558 78720 240110
rect 78784 237386 78812 241590
rect 79336 240174 79364 241590
rect 79324 240168 79376 240174
rect 79324 240110 79376 240116
rect 80060 240168 80112 240174
rect 80060 240110 80112 240116
rect 79416 237448 79468 237454
rect 79416 237390 79468 237396
rect 78772 237380 78824 237386
rect 78772 237322 78824 237328
rect 79324 236700 79376 236706
rect 79324 236642 79376 236648
rect 78680 232552 78732 232558
rect 78680 232494 78732 232500
rect 79336 175273 79364 236642
rect 79428 199442 79456 237390
rect 80072 226302 80100 240110
rect 80164 238678 80192 241590
rect 80152 238672 80204 238678
rect 80152 238614 80204 238620
rect 80164 237454 80192 238614
rect 80152 237448 80204 237454
rect 80152 237390 80204 237396
rect 80348 230450 80376 241590
rect 80992 240174 81020 241590
rect 80980 240168 81032 240174
rect 80980 240110 81032 240116
rect 82188 240106 82216 241590
rect 82280 241590 82432 241618
rect 82924 241590 82984 241618
rect 83752 241590 84088 241618
rect 84304 241590 84640 241618
rect 84856 241590 85192 241618
rect 85744 241590 85854 241618
rect 82176 240100 82228 240106
rect 82176 240042 82228 240048
rect 82280 240009 82308 241590
rect 82820 240168 82872 240174
rect 82820 240110 82872 240116
rect 82266 240000 82322 240009
rect 82266 239935 82322 239944
rect 82280 238754 82308 239935
rect 82096 238726 82308 238754
rect 80336 230444 80388 230450
rect 80336 230386 80388 230392
rect 80060 226296 80112 226302
rect 80060 226238 80112 226244
rect 80704 222896 80756 222902
rect 80704 222838 80756 222844
rect 79416 199436 79468 199442
rect 79416 199378 79468 199384
rect 78678 175264 78734 175273
rect 78678 175199 78734 175208
rect 79322 175264 79378 175273
rect 79322 175199 79378 175208
rect 77956 151786 78168 151814
rect 77300 141432 77352 141438
rect 77300 141374 77352 141380
rect 78036 140072 78088 140078
rect 78036 140014 78088 140020
rect 76564 136740 76616 136746
rect 76564 136682 76616 136688
rect 77392 136740 77444 136746
rect 77392 136682 77444 136688
rect 76024 134830 76328 134858
rect 76300 134722 76328 134830
rect 73448 134694 73600 134722
rect 73816 134694 74152 134722
rect 74552 134694 74704 134722
rect 74828 134694 75256 134722
rect 75380 134694 75808 134722
rect 75932 134694 76176 134722
rect 76300 134694 76728 134722
rect 77404 134586 77432 136682
rect 78048 134722 78076 140014
rect 78140 138689 78168 151786
rect 78126 138680 78182 138689
rect 78126 138615 78182 138624
rect 78140 134994 78168 138615
rect 78692 134994 78720 175199
rect 78862 167648 78918 167657
rect 78862 167583 78918 167592
rect 78876 151814 78904 167583
rect 79966 157448 80022 157457
rect 79966 157383 80022 157392
rect 78876 151786 79456 151814
rect 79322 137320 79378 137329
rect 79322 137255 79378 137264
rect 78140 134966 78214 134994
rect 78692 134966 78766 134994
rect 77832 134694 78076 134722
rect 78186 134708 78214 134966
rect 78738 134708 78766 134966
rect 79336 134858 79364 137255
rect 79290 134830 79364 134858
rect 79290 134708 79318 134830
rect 79428 134722 79456 151786
rect 79980 136882 80008 157383
rect 80242 151872 80298 151881
rect 80242 151814 80298 151816
rect 80242 151807 80560 151814
rect 80256 151786 80560 151807
rect 80152 144832 80204 144838
rect 80152 144774 80204 144780
rect 79968 136876 80020 136882
rect 79968 136818 80020 136824
rect 80164 134722 80192 144774
rect 80532 134722 80560 151786
rect 80716 137465 80744 222838
rect 81438 153776 81494 153785
rect 81438 153711 81494 153720
rect 80702 137456 80758 137465
rect 80702 137391 80758 137400
rect 80980 136876 81032 136882
rect 80980 136818 81032 136824
rect 80992 134722 81020 136818
rect 81452 134722 81480 153711
rect 82096 152590 82124 238726
rect 82832 221474 82860 240110
rect 82924 235346 82952 241590
rect 83752 240174 83780 241590
rect 83740 240168 83792 240174
rect 83740 240110 83792 240116
rect 84200 240168 84252 240174
rect 84200 240110 84252 240116
rect 84106 238776 84162 238785
rect 84106 238711 84162 238720
rect 82912 235340 82964 235346
rect 82912 235282 82964 235288
rect 84016 227044 84068 227050
rect 84016 226986 84068 226992
rect 82820 221468 82872 221474
rect 82820 221410 82872 221416
rect 84028 204950 84056 226986
rect 84016 204944 84068 204950
rect 84016 204886 84068 204892
rect 84120 181490 84148 238711
rect 84212 227050 84240 240110
rect 84304 234569 84332 241590
rect 84856 240174 84884 241590
rect 85854 241567 85910 241576
rect 85960 241590 86296 241618
rect 87064 241590 87400 241618
rect 87616 241590 87952 241618
rect 88352 241590 88504 241618
rect 89056 241590 89392 241618
rect 89608 241590 89668 241618
rect 84844 240168 84896 240174
rect 84844 240110 84896 240116
rect 85960 238754 85988 241590
rect 86960 240168 87012 240174
rect 86960 240110 87012 240116
rect 86868 240100 86920 240106
rect 86868 240042 86920 240048
rect 86880 239465 86908 240042
rect 86866 239456 86922 239465
rect 86866 239391 86922 239400
rect 85592 238726 85988 238754
rect 85592 237182 85620 238726
rect 85580 237176 85632 237182
rect 85580 237118 85632 237124
rect 84290 234560 84346 234569
rect 84290 234495 84346 234504
rect 84200 227044 84252 227050
rect 84200 226986 84252 226992
rect 86866 226400 86922 226409
rect 86866 226335 86922 226344
rect 84108 181484 84160 181490
rect 84108 181426 84160 181432
rect 86222 171184 86278 171193
rect 86222 171119 86278 171128
rect 83462 169008 83518 169017
rect 83462 168943 83518 168952
rect 82912 166320 82964 166326
rect 82912 166262 82964 166268
rect 82084 152584 82136 152590
rect 82084 152526 82136 152532
rect 81992 151088 82044 151094
rect 81992 151030 82044 151036
rect 82004 134722 82032 151030
rect 82820 143744 82872 143750
rect 82820 143686 82872 143692
rect 82832 134994 82860 143686
rect 82786 134966 82860 134994
rect 79428 134694 79856 134722
rect 80164 134694 80408 134722
rect 80532 134694 80776 134722
rect 80992 134694 81328 134722
rect 81452 134694 81880 134722
rect 82004 134694 82432 134722
rect 82786 134708 82814 134966
rect 82924 134722 82952 166262
rect 83476 144838 83504 168943
rect 83464 144832 83516 144838
rect 83464 144774 83516 144780
rect 85580 144492 85632 144498
rect 85580 144434 85632 144440
rect 83002 143576 83058 143585
rect 83002 143511 83058 143520
rect 83016 138825 83044 143511
rect 83462 142488 83518 142497
rect 83462 142423 83518 142432
rect 83002 138816 83058 138825
rect 83002 138751 83058 138760
rect 83476 134722 83504 142423
rect 84752 139392 84804 139398
rect 84752 139334 84804 139340
rect 84658 138816 84714 138825
rect 84658 138751 84714 138760
rect 84672 134722 84700 138751
rect 84764 138009 84792 139334
rect 84750 138000 84806 138009
rect 84750 137935 84806 137944
rect 82924 134694 83352 134722
rect 83476 134694 83904 134722
rect 84456 134694 84700 134722
rect 84764 134722 84792 137935
rect 85488 136740 85540 136746
rect 85488 136682 85540 136688
rect 85500 134722 85528 136682
rect 84764 134694 85008 134722
rect 85376 134694 85528 134722
rect 85592 134722 85620 144434
rect 86236 136746 86264 171119
rect 86314 168464 86370 168473
rect 86314 168399 86370 168408
rect 86328 143750 86356 168399
rect 86316 143744 86368 143750
rect 86316 143686 86368 143692
rect 86880 139466 86908 226335
rect 86972 214606 87000 240110
rect 87064 227050 87092 241590
rect 87616 240174 87644 241590
rect 87604 240168 87656 240174
rect 87604 240110 87656 240116
rect 87602 239864 87658 239873
rect 87602 239799 87658 239808
rect 87052 227044 87104 227050
rect 87052 226986 87104 226992
rect 86960 214600 87012 214606
rect 86960 214542 87012 214548
rect 87616 178702 87644 239799
rect 87696 233912 87748 233918
rect 87696 233854 87748 233860
rect 87708 193866 87736 233854
rect 88246 220960 88302 220969
rect 88246 220895 88302 220904
rect 87696 193860 87748 193866
rect 87696 193802 87748 193808
rect 87604 178696 87656 178702
rect 87604 178638 87656 178644
rect 88260 177342 88288 220895
rect 88352 220794 88380 241590
rect 89076 239420 89128 239426
rect 89076 239362 89128 239368
rect 88984 237176 89036 237182
rect 88984 237118 89036 237124
rect 88340 220788 88392 220794
rect 88340 220730 88392 220736
rect 88248 177336 88300 177342
rect 88248 177278 88300 177284
rect 88260 176730 88288 177278
rect 87604 176724 87656 176730
rect 87604 176666 87656 176672
rect 88248 176724 88300 176730
rect 88248 176666 88300 176672
rect 86960 164280 87012 164286
rect 86960 164222 87012 164228
rect 86868 139460 86920 139466
rect 86868 139402 86920 139408
rect 86224 136740 86276 136746
rect 86224 136682 86276 136688
rect 86880 134722 86908 139402
rect 86972 134994 87000 164222
rect 87144 162920 87196 162926
rect 87144 162862 87196 162868
rect 86972 134966 87046 134994
rect 85592 134694 85928 134722
rect 86480 134694 86908 134722
rect 87018 134708 87046 134966
rect 87156 134722 87184 162862
rect 87512 146260 87564 146266
rect 87512 146202 87564 146208
rect 87524 138014 87552 146202
rect 87616 140078 87644 176666
rect 88996 175982 89024 237118
rect 89088 231810 89116 239362
rect 89364 238814 89392 241590
rect 89640 240106 89668 241590
rect 90284 241590 90712 241618
rect 91112 241590 91264 241618
rect 89628 240100 89680 240106
rect 89628 240042 89680 240048
rect 89352 238808 89404 238814
rect 89352 238750 89404 238756
rect 90284 238754 90312 241590
rect 90914 240136 90970 240145
rect 90914 240071 90970 240080
rect 89732 238726 90312 238754
rect 89076 231804 89128 231810
rect 89076 231746 89128 231752
rect 89732 229090 89760 238726
rect 89720 229084 89772 229090
rect 89720 229026 89772 229032
rect 90822 227080 90878 227089
rect 90822 227015 90878 227024
rect 88984 175976 89036 175982
rect 88984 175918 89036 175924
rect 89074 175400 89130 175409
rect 89074 175335 89130 175344
rect 88984 158840 89036 158846
rect 88984 158782 89036 158788
rect 88338 154592 88394 154601
rect 88338 154527 88394 154536
rect 88248 147008 88300 147014
rect 88248 146950 88300 146956
rect 88260 146266 88288 146950
rect 88248 146260 88300 146266
rect 88248 146202 88300 146208
rect 87604 140072 87656 140078
rect 87604 140014 87656 140020
rect 88352 138106 88380 154527
rect 88616 142316 88668 142322
rect 88616 142258 88668 142264
rect 88524 141432 88576 141438
rect 88524 141374 88576 141380
rect 88340 138100 88392 138106
rect 88340 138042 88392 138048
rect 87524 137986 87736 138014
rect 87708 134722 87736 137986
rect 88536 134994 88564 141374
rect 88490 134966 88564 134994
rect 87156 134694 87584 134722
rect 87708 134694 87952 134722
rect 88490 134708 88518 134966
rect 88628 134722 88656 142258
rect 88996 140826 89024 158782
rect 89088 144498 89116 175335
rect 90836 173942 90864 227015
rect 90928 184210 90956 240071
rect 91112 236314 91140 241590
rect 92216 238754 92244 241726
rect 95344 241726 95882 241754
rect 94964 241664 95016 241670
rect 92354 241505 92382 241604
rect 92492 241590 92920 241618
rect 92340 241496 92396 241505
rect 92340 241431 92396 241440
rect 92216 238726 92428 238754
rect 91020 236286 91140 236314
rect 91020 233918 91048 236286
rect 91008 233912 91060 233918
rect 91008 233854 91060 233860
rect 91008 232552 91060 232558
rect 91008 232494 91060 232500
rect 90916 184204 90968 184210
rect 90916 184146 90968 184152
rect 89720 173936 89772 173942
rect 89720 173878 89772 173884
rect 90824 173936 90876 173942
rect 90824 173878 90876 173884
rect 89168 172576 89220 172582
rect 89168 172518 89220 172524
rect 89180 158030 89208 172518
rect 89168 158024 89220 158030
rect 89168 157966 89220 157972
rect 89732 151814 89760 173878
rect 91020 167793 91048 232494
rect 92400 198014 92428 238726
rect 92492 232529 92520 241590
rect 93458 241369 93486 241604
rect 93872 241590 94024 241618
rect 94148 241590 94576 241618
rect 95016 241612 95128 241618
rect 94964 241606 95128 241612
rect 94976 241590 95128 241606
rect 93122 241360 93178 241369
rect 93122 241295 93178 241304
rect 93444 241360 93500 241369
rect 93444 241295 93500 241304
rect 92478 232520 92534 232529
rect 92478 232455 92534 232464
rect 93136 207126 93164 241295
rect 93768 238740 93820 238746
rect 93768 238682 93820 238688
rect 93124 207120 93176 207126
rect 93124 207062 93176 207068
rect 92388 198008 92440 198014
rect 92388 197950 92440 197956
rect 91192 176724 91244 176730
rect 91192 176666 91244 176672
rect 91006 167784 91062 167793
rect 91006 167719 91062 167728
rect 91008 160744 91060 160750
rect 91008 160686 91060 160692
rect 91020 151814 91048 160686
rect 89732 151786 89852 151814
rect 89076 144492 89128 144498
rect 89076 144434 89128 144440
rect 88984 140820 89036 140826
rect 88984 140762 89036 140768
rect 88996 137766 89024 140762
rect 89260 138100 89312 138106
rect 89260 138042 89312 138048
rect 88984 137760 89036 137766
rect 88984 137702 89036 137708
rect 89272 134722 89300 138042
rect 89718 136776 89774 136785
rect 89718 136711 89774 136720
rect 89732 134722 89760 136711
rect 89824 134858 89852 151786
rect 90836 151786 91048 151814
rect 91204 151814 91232 176666
rect 92662 166288 92718 166297
rect 92662 166223 92718 166232
rect 91204 151786 91784 151814
rect 89904 142384 89956 142390
rect 89904 142326 89956 142332
rect 89916 139534 89944 142326
rect 89994 139632 90050 139641
rect 89994 139567 90050 139576
rect 89904 139528 89956 139534
rect 89904 139470 89956 139476
rect 90008 136649 90036 139567
rect 89994 136640 90050 136649
rect 89994 136575 90050 136584
rect 90836 135998 90864 151786
rect 90916 142248 90968 142254
rect 90916 142190 90968 142196
rect 90928 139398 90956 142190
rect 91098 140856 91154 140865
rect 91098 140791 91154 140800
rect 90916 139392 90968 139398
rect 90916 139334 90968 139340
rect 91112 137873 91140 140791
rect 91098 137864 91154 137873
rect 91098 137799 91154 137808
rect 91192 137760 91244 137766
rect 91192 137702 91244 137708
rect 90824 135992 90876 135998
rect 90824 135934 90876 135940
rect 89824 134830 90128 134858
rect 90100 134722 90128 134830
rect 88628 134694 89056 134722
rect 89272 134694 89608 134722
rect 89732 134694 89976 134722
rect 90100 134694 90528 134722
rect 91204 134586 91232 137702
rect 91284 135992 91336 135998
rect 91284 135934 91336 135940
rect 91296 134722 91324 135934
rect 91756 134722 91784 151786
rect 92570 136776 92626 136785
rect 92570 136711 92626 136720
rect 92584 134858 92612 136711
rect 92538 134830 92612 134858
rect 91296 134694 91632 134722
rect 91756 134694 92184 134722
rect 92538 134708 92566 134830
rect 92676 134722 92704 166223
rect 93674 140856 93730 140865
rect 93674 140791 93730 140800
rect 93688 134994 93716 140791
rect 93642 134966 93716 134994
rect 92676 134694 93104 134722
rect 93642 134708 93670 134966
rect 93780 134638 93808 238682
rect 93872 205018 93900 241590
rect 93952 241528 94004 241534
rect 93952 241470 94004 241476
rect 93964 237425 93992 241470
rect 93950 237416 94006 237425
rect 93950 237351 94006 237360
rect 94148 236745 94176 241590
rect 95240 240168 95292 240174
rect 95240 240110 95292 240116
rect 95056 237448 95108 237454
rect 95056 237390 95108 237396
rect 94134 236736 94190 236745
rect 94134 236671 94190 236680
rect 94688 233980 94740 233986
rect 94688 233922 94740 233928
rect 93860 205012 93912 205018
rect 93860 204954 93912 204960
rect 93860 153264 93912 153270
rect 93860 153206 93912 153212
rect 93872 151814 93900 153206
rect 93872 151786 94360 151814
rect 94226 140040 94282 140049
rect 94226 139975 94282 139984
rect 94240 134994 94268 139975
rect 94194 134966 94268 134994
rect 94194 134708 94222 134966
rect 94332 134722 94360 151786
rect 94504 136672 94556 136678
rect 94504 136614 94556 136620
rect 94516 135250 94544 136614
rect 94504 135244 94556 135250
rect 94504 135186 94556 135192
rect 94332 134694 94576 134722
rect 77280 134558 77432 134586
rect 91080 134558 91232 134586
rect 93768 134632 93820 134638
rect 93768 134574 93820 134580
rect 67914 128208 67970 128217
rect 67914 128143 67970 128152
rect 67822 112432 67878 112441
rect 67822 112367 67878 112376
rect 94596 102808 94648 102814
rect 94596 102750 94648 102756
rect 67822 101008 67878 101017
rect 67822 100943 67878 100952
rect 67836 84182 67864 100943
rect 68284 95192 68336 95198
rect 68284 95134 68336 95140
rect 67914 93936 67970 93945
rect 67914 93871 67970 93880
rect 67928 93838 67956 93871
rect 67916 93832 67968 93838
rect 67916 93774 67968 93780
rect 67824 84176 67876 84182
rect 67824 84118 67876 84124
rect 68296 81297 68324 95134
rect 68468 92880 68520 92886
rect 68520 92828 68816 92834
rect 68468 92822 68816 92828
rect 68480 92806 68816 92822
rect 69170 92562 69198 92820
rect 69722 92721 69750 92820
rect 69708 92712 69764 92721
rect 70274 92698 70302 92820
rect 70274 92670 70348 92698
rect 69708 92647 69764 92656
rect 69722 92562 69750 92647
rect 69170 92534 69244 92562
rect 69216 85474 69244 92534
rect 69676 92534 69750 92562
rect 69204 85468 69256 85474
rect 69204 85410 69256 85416
rect 69676 84194 69704 92534
rect 70320 90982 70348 92670
rect 70826 92562 70854 92820
rect 71194 92721 71222 92820
rect 71746 92750 71774 92820
rect 71734 92744 71786 92750
rect 71180 92712 71236 92721
rect 71734 92686 71786 92692
rect 71180 92647 71236 92656
rect 70412 92534 70854 92562
rect 71780 92608 71832 92614
rect 72298 92562 72326 92820
rect 72850 92562 72878 92820
rect 73402 92698 73430 92820
rect 73770 92698 73798 92820
rect 71780 92550 71832 92556
rect 70308 90976 70360 90982
rect 70308 90918 70360 90924
rect 70320 90302 70348 90918
rect 70308 90296 70360 90302
rect 70308 90238 70360 90244
rect 69216 84166 69704 84194
rect 68282 81288 68338 81297
rect 68282 81223 68338 81232
rect 69216 69018 69244 84166
rect 70412 84114 70440 92534
rect 71792 91089 71820 92550
rect 71884 92534 72326 92562
rect 72804 92534 72878 92562
rect 73356 92670 73430 92698
rect 73724 92670 73798 92698
rect 71778 91080 71834 91089
rect 71778 91015 71834 91024
rect 71044 90296 71096 90302
rect 71044 90238 71096 90244
rect 70400 84108 70452 84114
rect 70400 84050 70452 84056
rect 70306 82104 70362 82113
rect 70306 82039 70362 82048
rect 69204 69012 69256 69018
rect 69204 68954 69256 68960
rect 68928 37936 68980 37942
rect 68928 37878 68980 37884
rect 67732 36576 67784 36582
rect 67732 36518 67784 36524
rect 68940 3534 68968 37878
rect 70216 13116 70268 13122
rect 70216 13058 70268 13064
rect 70228 3534 70256 13058
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 65432 2100 65484 2106
rect 65432 2042 65484 2048
rect 65536 480 65564 3470
rect 66732 480 66760 3470
rect 67928 480 67956 3470
rect 69124 480 69152 3470
rect 70320 480 70348 82039
rect 71056 62014 71084 90238
rect 71792 86873 71820 91015
rect 71778 86864 71834 86873
rect 71778 86799 71834 86808
rect 71688 69692 71740 69698
rect 71688 69634 71740 69640
rect 71044 62008 71096 62014
rect 71044 61950 71096 61956
rect 71700 6914 71728 69634
rect 71884 67590 71912 92534
rect 72804 92478 72832 92534
rect 72792 92472 72844 92478
rect 73356 92449 73384 92670
rect 72792 92414 72844 92420
rect 73342 92440 73398 92449
rect 73342 92375 73398 92384
rect 73724 91050 73752 92670
rect 74322 92562 74350 92820
rect 74276 92534 74350 92562
rect 74540 92608 74592 92614
rect 74874 92562 74902 92820
rect 74540 92550 74592 92556
rect 73712 91044 73764 91050
rect 73712 90986 73764 90992
rect 73724 88262 73752 90986
rect 74276 90817 74304 92534
rect 74262 90808 74318 90817
rect 74262 90743 74318 90752
rect 73712 88256 73764 88262
rect 73712 88198 73764 88204
rect 74276 84194 74304 90743
rect 73816 84166 74304 84194
rect 71872 67584 71924 67590
rect 71872 67526 71924 67532
rect 73816 57866 73844 84166
rect 73804 57860 73856 57866
rect 73804 57802 73856 57808
rect 74552 56574 74580 92550
rect 74828 92534 74902 92562
rect 75426 92562 75454 92820
rect 75794 92614 75822 92820
rect 76346 92698 76374 92820
rect 76300 92670 76374 92698
rect 75782 92608 75834 92614
rect 75426 92534 75500 92562
rect 75782 92550 75834 92556
rect 74828 89622 74856 92534
rect 75472 92478 75500 92534
rect 75460 92472 75512 92478
rect 75460 92414 75512 92420
rect 76300 90953 76328 92670
rect 76898 92562 76926 92820
rect 77450 92562 77478 92820
rect 76576 92534 76926 92562
rect 77312 92534 77478 92562
rect 78002 92562 78030 92820
rect 78370 92562 78398 92820
rect 78922 92562 78950 92820
rect 79474 92562 79502 92820
rect 78002 92534 78076 92562
rect 78370 92534 78444 92562
rect 78922 92534 78996 92562
rect 76286 90944 76342 90953
rect 76286 90879 76342 90888
rect 74816 89616 74868 89622
rect 74816 89558 74868 89564
rect 76576 84194 76604 92534
rect 75932 84166 76604 84194
rect 75932 82822 75960 84166
rect 75920 82816 75972 82822
rect 75920 82758 75972 82764
rect 77312 81161 77340 92534
rect 78048 89593 78076 92534
rect 78034 89584 78090 89593
rect 78034 89519 78090 89528
rect 78416 85377 78444 92534
rect 78968 90370 78996 92534
rect 79428 92534 79502 92562
rect 80026 92562 80054 92820
rect 80578 92562 80606 92820
rect 80026 92534 80100 92562
rect 78956 90364 79008 90370
rect 78956 90306 79008 90312
rect 79428 88330 79456 92534
rect 79416 88324 79468 88330
rect 79416 88266 79468 88272
rect 80072 86970 80100 92534
rect 80164 92534 80606 92562
rect 80946 92562 80974 92820
rect 81498 92562 81526 92820
rect 80946 92534 81020 92562
rect 80060 86964 80112 86970
rect 80060 86906 80112 86912
rect 78402 85368 78458 85377
rect 78402 85303 78458 85312
rect 80164 81394 80192 92534
rect 80992 87961 81020 92534
rect 81452 92534 81526 92562
rect 81624 92608 81676 92614
rect 82050 92562 82078 92820
rect 82602 92614 82630 92820
rect 82970 92698 82998 92820
rect 82970 92670 83044 92698
rect 81624 92550 81676 92556
rect 81452 92410 81480 92534
rect 81440 92404 81492 92410
rect 81440 92346 81492 92352
rect 80978 87952 81034 87961
rect 80978 87887 81034 87896
rect 80152 81388 80204 81394
rect 80152 81330 80204 81336
rect 77298 81152 77354 81161
rect 77298 81087 77354 81096
rect 81636 74526 81664 92550
rect 81728 92534 82078 92562
rect 82590 92608 82642 92614
rect 82590 92550 82642 92556
rect 81728 80034 81756 92534
rect 83016 89729 83044 92670
rect 83522 92562 83550 92820
rect 83200 92534 83550 92562
rect 84074 92562 84102 92820
rect 84626 92698 84654 92820
rect 84626 92670 84700 92698
rect 84074 92534 84148 92562
rect 83002 89720 83058 89729
rect 83002 89655 83058 89664
rect 83200 84194 83228 92534
rect 84120 86601 84148 92534
rect 84672 92313 84700 92670
rect 85178 92562 85206 92820
rect 84856 92534 85206 92562
rect 85546 92562 85574 92820
rect 86098 92562 86126 92820
rect 85546 92534 85620 92562
rect 84658 92304 84714 92313
rect 84658 92239 84714 92248
rect 84106 86592 84162 86601
rect 84106 86527 84162 86536
rect 84856 84194 84884 92534
rect 82832 84166 83228 84194
rect 84212 84166 84884 84194
rect 81716 80028 81768 80034
rect 81716 79970 81768 79976
rect 82832 78606 82860 84166
rect 84212 82754 84240 84166
rect 84200 82748 84252 82754
rect 84200 82690 84252 82696
rect 82820 78600 82872 78606
rect 82820 78542 82872 78548
rect 81624 74520 81676 74526
rect 81624 74462 81676 74468
rect 75828 65544 75880 65550
rect 75828 65486 75880 65492
rect 74540 56568 74592 56574
rect 74540 56510 74592 56516
rect 73068 54528 73120 54534
rect 73068 54470 73120 54476
rect 71516 6886 71728 6914
rect 71516 480 71544 6886
rect 73080 3534 73108 54470
rect 75184 35216 75236 35222
rect 75184 35158 75236 35164
rect 74448 21412 74500 21418
rect 74448 21354 74500 21360
rect 74460 3534 74488 21354
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 72620 480 72648 3470
rect 73816 480 73844 3470
rect 75012 480 75040 3470
rect 75196 3466 75224 35158
rect 75840 3534 75868 65486
rect 85592 64870 85620 92534
rect 85684 92534 86126 92562
rect 86650 92562 86678 92820
rect 86960 92608 87012 92614
rect 86650 92534 86724 92562
rect 86960 92550 87012 92556
rect 87202 92562 87230 92820
rect 87570 92750 87598 92820
rect 87558 92744 87610 92750
rect 87558 92686 87610 92692
rect 87570 92562 87598 92686
rect 88122 92614 88150 92820
rect 88110 92608 88162 92614
rect 85684 84017 85712 92534
rect 86696 92177 86724 92534
rect 86682 92168 86738 92177
rect 86682 92103 86738 92112
rect 85670 84008 85726 84017
rect 85670 83943 85726 83952
rect 86866 77888 86922 77897
rect 86866 77823 86922 77832
rect 85580 64864 85632 64870
rect 85580 64806 85632 64812
rect 85488 62892 85540 62898
rect 85488 62834 85540 62840
rect 81348 62824 81400 62830
rect 81348 62766 81400 62772
rect 77208 43444 77260 43450
rect 77208 43386 77260 43392
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 75184 3460 75236 3466
rect 75184 3402 75236 3408
rect 77220 3262 77248 43386
rect 79324 42084 79376 42090
rect 79324 42026 79376 42032
rect 78588 22772 78640 22778
rect 78588 22714 78640 22720
rect 77392 3460 77444 3466
rect 77392 3402 77444 3408
rect 76196 3256 76248 3262
rect 76196 3198 76248 3204
rect 77208 3256 77260 3262
rect 77208 3198 77260 3204
rect 76208 480 76236 3198
rect 77404 480 77432 3402
rect 78600 480 78628 22714
rect 79336 2174 79364 42026
rect 79692 10328 79744 10334
rect 79692 10270 79744 10276
rect 79324 2168 79376 2174
rect 79324 2110 79376 2116
rect 79704 480 79732 10270
rect 81360 3534 81388 62766
rect 82728 39364 82780 39370
rect 82728 39306 82780 39312
rect 82740 3534 82768 39306
rect 84108 11756 84160 11762
rect 84108 11698 84160 11704
rect 84120 3534 84148 11698
rect 85500 3534 85528 62834
rect 86776 28280 86828 28286
rect 86776 28222 86828 28228
rect 86788 3534 86816 28222
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 84108 3528 84160 3534
rect 84108 3470 84160 3476
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 85672 3528 85724 3534
rect 85672 3470 85724 3476
rect 86776 3528 86828 3534
rect 86776 3470 86828 3476
rect 80900 480 80928 3470
rect 82096 480 82124 3470
rect 83292 480 83320 3470
rect 84488 480 84516 3470
rect 85684 480 85712 3470
rect 86880 480 86908 77823
rect 86972 73166 87000 92550
rect 87202 92534 87276 92562
rect 87570 92534 87644 92562
rect 88674 92562 88702 92820
rect 88110 92550 88162 92556
rect 87248 88097 87276 92534
rect 87616 88330 87644 92534
rect 88352 92534 88702 92562
rect 89226 92562 89254 92820
rect 89778 92562 89806 92820
rect 89226 92534 89300 92562
rect 87604 88324 87656 88330
rect 87604 88266 87656 88272
rect 88156 88324 88208 88330
rect 88156 88266 88208 88272
rect 87234 88088 87290 88097
rect 87234 88023 87290 88032
rect 86960 73160 87012 73166
rect 86960 73102 87012 73108
rect 88168 62082 88196 88266
rect 88352 77246 88380 92534
rect 89272 89622 89300 92534
rect 89732 92534 89806 92562
rect 89904 92608 89956 92614
rect 90146 92562 90174 92820
rect 90698 92614 90726 92820
rect 89904 92550 89956 92556
rect 89260 89616 89312 89622
rect 89260 89558 89312 89564
rect 89732 81326 89760 92534
rect 89720 81320 89772 81326
rect 89720 81262 89772 81268
rect 89916 80073 89944 92550
rect 90008 92534 90174 92562
rect 90686 92608 90738 92614
rect 90686 92550 90738 92556
rect 91250 92562 91278 92820
rect 91802 92562 91830 92820
rect 92354 92562 92382 92820
rect 92722 92562 92750 92820
rect 93274 92721 93302 92820
rect 93826 92750 93854 92820
rect 94392 92806 94544 92834
rect 93814 92744 93866 92750
rect 93260 92712 93316 92721
rect 93814 92686 93866 92692
rect 93260 92647 93316 92656
rect 93274 92562 93302 92647
rect 93826 92562 93854 92686
rect 91250 92534 91324 92562
rect 91802 92534 91876 92562
rect 92354 92534 92428 92562
rect 92722 92534 92796 92562
rect 93274 92534 93348 92562
rect 93826 92534 93900 92562
rect 94516 92546 94544 92806
rect 90008 82793 90036 92534
rect 91296 85241 91324 92534
rect 91848 92449 91876 92534
rect 91834 92440 91890 92449
rect 92400 92410 92428 92534
rect 91834 92375 91890 92384
rect 92388 92404 92440 92410
rect 92388 92346 92440 92352
rect 92768 86737 92796 92534
rect 92754 86728 92810 86737
rect 92754 86663 92810 86672
rect 91282 85232 91338 85241
rect 91282 85167 91338 85176
rect 93320 84194 93348 92534
rect 93872 84194 93900 92534
rect 94504 92540 94556 92546
rect 94504 92482 94556 92488
rect 93320 84166 93808 84194
rect 93872 84166 94544 84194
rect 94608 84182 94636 102750
rect 94700 92750 94728 233922
rect 95068 153270 95096 237390
rect 95148 226364 95200 226370
rect 95148 226306 95200 226312
rect 95056 153264 95108 153270
rect 95056 153206 95108 153212
rect 95160 103601 95188 226306
rect 95252 206310 95280 240110
rect 95344 233986 95372 241726
rect 95882 241703 95938 241712
rect 95896 241590 96232 241618
rect 96724 241590 96784 241618
rect 97336 241590 97580 241618
rect 95896 240174 95924 241590
rect 95976 241528 96028 241534
rect 95976 241470 96028 241476
rect 95884 240168 95936 240174
rect 95884 240110 95936 240116
rect 95988 238678 96016 241470
rect 96620 240168 96672 240174
rect 96620 240110 96672 240116
rect 96526 238776 96582 238785
rect 96526 238711 96582 238720
rect 95976 238672 96028 238678
rect 95976 238614 96028 238620
rect 95332 233980 95384 233986
rect 95332 233922 95384 233928
rect 96068 207120 96120 207126
rect 96068 207062 96120 207068
rect 95240 206304 95292 206310
rect 95240 206246 95292 206252
rect 95884 199504 95936 199510
rect 95884 199446 95936 199452
rect 95240 134632 95292 134638
rect 95240 134574 95292 134580
rect 95146 103592 95202 103601
rect 95146 103527 95202 103536
rect 95252 92818 95280 134574
rect 95330 120320 95386 120329
rect 95330 120255 95386 120264
rect 95240 92812 95292 92818
rect 95240 92754 95292 92760
rect 94688 92744 94740 92750
rect 94688 92686 94740 92692
rect 93122 83464 93178 83473
rect 93122 83399 93178 83408
rect 89994 82784 90050 82793
rect 89994 82719 90050 82728
rect 89902 80064 89958 80073
rect 89902 79999 89958 80008
rect 90364 79348 90416 79354
rect 90364 79290 90416 79296
rect 88340 77240 88392 77246
rect 88340 77182 88392 77188
rect 88248 71052 88300 71058
rect 88248 70994 88300 71000
rect 88156 62076 88208 62082
rect 88156 62018 88208 62024
rect 88260 6914 88288 70994
rect 89628 68332 89680 68338
rect 89628 68274 89680 68280
rect 87984 6886 88288 6914
rect 87984 480 88012 6886
rect 89640 3534 89668 68274
rect 90376 6914 90404 79290
rect 93136 20670 93164 83399
rect 93780 57934 93808 84166
rect 94516 70378 94544 84166
rect 94596 84176 94648 84182
rect 94596 84118 94648 84124
rect 95344 76566 95372 120255
rect 95516 94512 95568 94518
rect 95516 94454 95568 94460
rect 95528 88262 95556 94454
rect 95896 92993 95924 199446
rect 95976 178084 96028 178090
rect 95976 178026 96028 178032
rect 95988 105097 96016 178026
rect 96080 134065 96108 207062
rect 96540 200802 96568 238711
rect 96632 231878 96660 240110
rect 96724 234025 96752 241590
rect 97552 240145 97580 241590
rect 97644 241590 97888 241618
rect 97644 240174 97672 241590
rect 97632 240168 97684 240174
rect 97538 240136 97594 240145
rect 97632 240110 97684 240116
rect 97538 240071 97594 240080
rect 97908 236020 97960 236026
rect 97908 235962 97960 235968
rect 96710 234016 96766 234025
rect 96710 233951 96766 233960
rect 97814 234016 97870 234025
rect 97814 233951 97870 233960
rect 96620 231872 96672 231878
rect 96620 231814 96672 231820
rect 97264 231872 97316 231878
rect 97264 231814 97316 231820
rect 97276 209098 97304 231814
rect 97264 209092 97316 209098
rect 97264 209034 97316 209040
rect 96528 200796 96580 200802
rect 96528 200738 96580 200744
rect 97828 155174 97856 233951
rect 97264 155168 97316 155174
rect 97264 155110 97316 155116
rect 97816 155168 97868 155174
rect 97816 155110 97868 155116
rect 96710 145752 96766 145761
rect 96710 145687 96766 145696
rect 96160 139528 96212 139534
rect 96160 139470 96212 139476
rect 96066 134056 96122 134065
rect 96066 133991 96122 134000
rect 96172 132462 96200 139470
rect 96620 133884 96672 133890
rect 96620 133826 96672 133832
rect 96632 133113 96660 133826
rect 96618 133104 96674 133113
rect 96618 133039 96674 133048
rect 96160 132456 96212 132462
rect 96160 132398 96212 132404
rect 96620 132388 96672 132394
rect 96620 132330 96672 132336
rect 96632 132297 96660 132330
rect 96618 132288 96674 132297
rect 96618 132223 96674 132232
rect 96618 130928 96674 130937
rect 96618 130863 96674 130872
rect 96632 130422 96660 130863
rect 96620 130416 96672 130422
rect 96540 130364 96620 130370
rect 96540 130358 96672 130364
rect 96540 130342 96660 130358
rect 96540 129962 96568 130342
rect 96620 130212 96672 130218
rect 96620 130154 96672 130160
rect 96632 130121 96660 130154
rect 96618 130112 96674 130121
rect 96618 130047 96674 130056
rect 96540 129934 96660 129962
rect 96068 120352 96120 120358
rect 96066 120320 96068 120329
rect 96120 120320 96122 120329
rect 96066 120255 96122 120264
rect 95974 105088 96030 105097
rect 95974 105023 96030 105032
rect 96528 103556 96580 103562
rect 96528 103498 96580 103504
rect 96540 103465 96568 103498
rect 96526 103456 96582 103465
rect 96526 103391 96582 103400
rect 95882 92984 95938 92993
rect 95882 92919 95938 92928
rect 95896 92478 95924 92919
rect 95884 92472 95936 92478
rect 95884 92414 95936 92420
rect 95516 88256 95568 88262
rect 95516 88198 95568 88204
rect 96632 83473 96660 129934
rect 96724 127673 96752 145687
rect 96804 135176 96856 135182
rect 96804 135118 96856 135124
rect 96816 133929 96844 135118
rect 96802 133920 96858 133929
rect 96802 133855 96858 133864
rect 96710 127664 96766 127673
rect 96710 127599 96766 127608
rect 97080 127628 97132 127634
rect 97080 127570 97132 127576
rect 97092 124681 97120 127570
rect 97078 124672 97134 124681
rect 97078 124607 97134 124616
rect 97172 124092 97224 124098
rect 97172 124034 97224 124040
rect 97184 123321 97212 124034
rect 97170 123312 97226 123321
rect 97170 123247 97226 123256
rect 97276 122505 97304 155110
rect 97356 144084 97408 144090
rect 97356 144026 97408 144032
rect 97368 131481 97396 144026
rect 97354 131472 97410 131481
rect 97354 131407 97410 131416
rect 97540 128308 97592 128314
rect 97540 128250 97592 128256
rect 97552 127129 97580 128250
rect 97538 127120 97594 127129
rect 97538 127055 97594 127064
rect 97816 126948 97868 126954
rect 97816 126890 97868 126896
rect 97828 126313 97856 126890
rect 97814 126304 97870 126313
rect 97814 126239 97870 126248
rect 97816 124160 97868 124166
rect 97814 124128 97816 124137
rect 97868 124128 97870 124137
rect 97814 124063 97870 124072
rect 97540 122800 97592 122806
rect 97540 122742 97592 122748
rect 97262 122496 97318 122505
rect 97262 122431 97318 122440
rect 97552 121689 97580 122742
rect 97538 121680 97594 121689
rect 97538 121615 97594 121624
rect 96988 121440 97040 121446
rect 96988 121382 97040 121388
rect 97000 120873 97028 121382
rect 96986 120864 97042 120873
rect 96986 120799 97042 120808
rect 97920 120170 97948 235962
rect 97736 120142 97948 120170
rect 97356 117224 97408 117230
rect 97356 117166 97408 117172
rect 97368 117065 97396 117166
rect 97354 117056 97410 117065
rect 97354 116991 97410 117000
rect 97736 114050 97764 120142
rect 97908 120080 97960 120086
rect 97908 120022 97960 120028
rect 97920 119513 97948 120022
rect 97906 119504 97962 119513
rect 97906 119439 97962 119448
rect 97906 118688 97962 118697
rect 97906 118623 97908 118632
rect 97960 118623 97962 118632
rect 97908 118594 97960 118600
rect 97908 117292 97960 117298
rect 97908 117234 97960 117240
rect 97920 116521 97948 117234
rect 97906 116512 97962 116521
rect 97906 116447 97962 116456
rect 97816 115932 97868 115938
rect 97816 115874 97868 115880
rect 97828 114889 97856 115874
rect 97906 115696 97962 115705
rect 97906 115631 97962 115640
rect 97814 114880 97870 114889
rect 97814 114815 97870 114824
rect 97920 114578 97948 115631
rect 97908 114572 97960 114578
rect 97908 114514 97960 114520
rect 97814 114064 97870 114073
rect 97736 114022 97814 114050
rect 97814 113999 97816 114008
rect 97868 113999 97870 114008
rect 97816 113970 97868 113976
rect 97906 113520 97962 113529
rect 97906 113455 97962 113464
rect 97920 113218 97948 113455
rect 97908 113212 97960 113218
rect 97908 113154 97960 113160
rect 97080 111920 97132 111926
rect 97078 111888 97080 111897
rect 97132 111888 97134 111897
rect 97078 111823 97134 111832
rect 96712 111716 96764 111722
rect 96712 111658 96764 111664
rect 96724 111081 96752 111658
rect 96710 111072 96766 111081
rect 96710 111007 96766 111016
rect 97908 110424 97960 110430
rect 97908 110366 97960 110372
rect 97920 110265 97948 110366
rect 97906 110256 97962 110265
rect 97906 110191 97962 110200
rect 97814 109712 97870 109721
rect 97814 109647 97870 109656
rect 96710 107264 96766 107273
rect 96710 107199 96766 107208
rect 96724 106418 96752 107199
rect 97828 106962 97856 109647
rect 97908 108384 97960 108390
rect 97908 108326 97960 108332
rect 97920 108089 97948 108326
rect 97906 108080 97962 108089
rect 97906 108015 97962 108024
rect 97816 106956 97868 106962
rect 97816 106898 97868 106904
rect 96712 106412 96764 106418
rect 96712 106354 96764 106360
rect 96802 104272 96858 104281
rect 96802 104207 96858 104216
rect 96816 104174 96844 104207
rect 96804 104168 96856 104174
rect 96804 104110 96856 104116
rect 97906 102912 97962 102921
rect 98012 102898 98040 243510
rect 98104 237454 98132 277366
rect 98748 269822 98776 284815
rect 99380 284436 99432 284442
rect 99380 284378 99432 284384
rect 98920 283076 98972 283082
rect 98920 283018 98972 283024
rect 98828 283008 98880 283014
rect 98828 282950 98880 282956
rect 98840 271182 98868 282950
rect 98932 276690 98960 283018
rect 99392 280838 99420 284378
rect 99380 280832 99432 280838
rect 99380 280774 99432 280780
rect 99378 280256 99434 280265
rect 99378 280191 99434 280200
rect 98920 276684 98972 276690
rect 98920 276626 98972 276632
rect 98828 271176 98880 271182
rect 98828 271118 98880 271124
rect 98736 269816 98788 269822
rect 98736 269758 98788 269764
rect 98182 261352 98238 261361
rect 98182 261287 98238 261296
rect 98092 237448 98144 237454
rect 98092 237390 98144 237396
rect 98196 236026 98224 261287
rect 99286 258088 99342 258097
rect 99286 258023 99342 258032
rect 98274 248840 98330 248849
rect 98274 248775 98330 248784
rect 98288 243574 98316 248775
rect 98276 243568 98328 243574
rect 98276 243510 98328 243516
rect 98276 243432 98328 243438
rect 98276 243374 98328 243380
rect 98288 240009 98316 243374
rect 98734 242584 98790 242593
rect 98734 242519 98790 242528
rect 98748 241777 98776 242519
rect 99102 242448 99158 242457
rect 99102 242383 99158 242392
rect 98734 241768 98790 241777
rect 98734 241703 98790 241712
rect 98440 241590 98776 241618
rect 98748 240009 98776 241590
rect 99116 241534 99144 242383
rect 99104 241528 99156 241534
rect 99104 241470 99156 241476
rect 98274 240000 98330 240009
rect 98274 239935 98330 239944
rect 98734 240000 98790 240009
rect 98734 239935 98790 239944
rect 98184 236020 98236 236026
rect 98184 235962 98236 235968
rect 98644 207052 98696 207058
rect 98644 206994 98696 207000
rect 98460 125588 98512 125594
rect 98460 125530 98512 125536
rect 98472 125497 98500 125530
rect 98458 125488 98514 125497
rect 98458 125423 98514 125432
rect 98092 111852 98144 111858
rect 98092 111794 98144 111800
rect 98104 108905 98132 111794
rect 98090 108896 98146 108905
rect 98090 108831 98146 108840
rect 97962 102882 98040 102898
rect 97962 102876 98052 102882
rect 97962 102870 98000 102876
rect 97906 102847 97962 102856
rect 98000 102818 98052 102824
rect 97908 102128 97960 102134
rect 97906 102096 97908 102105
rect 97960 102096 97962 102105
rect 97906 102031 97962 102040
rect 97538 100464 97594 100473
rect 97538 100399 97594 100408
rect 97552 99414 97580 100399
rect 97908 100020 97960 100026
rect 97908 99962 97960 99968
rect 97920 99657 97948 99962
rect 97906 99648 97962 99657
rect 97906 99583 97962 99592
rect 97540 99408 97592 99414
rect 97540 99350 97592 99356
rect 97814 99104 97870 99113
rect 97814 99039 97870 99048
rect 97828 98122 97856 99039
rect 97906 98288 97962 98297
rect 97906 98223 97962 98232
rect 97816 98116 97868 98122
rect 97816 98058 97868 98064
rect 97920 98054 97948 98223
rect 97908 98048 97960 98054
rect 97908 97990 97960 97996
rect 98656 97782 98684 206994
rect 99300 147694 99328 258023
rect 98736 147688 98788 147694
rect 98736 147630 98788 147636
rect 99288 147688 99340 147694
rect 99288 147630 99340 147636
rect 98748 111722 98776 147630
rect 98826 146432 98882 146441
rect 98826 146367 98882 146376
rect 98840 120358 98868 146367
rect 99392 144090 99420 280191
rect 100036 272542 100064 297463
rect 100114 282976 100170 282985
rect 100114 282911 100170 282920
rect 100024 272536 100076 272542
rect 100024 272478 100076 272484
rect 100128 268462 100156 282911
rect 100116 268456 100168 268462
rect 100116 268398 100168 268404
rect 100022 259040 100078 259049
rect 100022 258975 100078 258984
rect 100036 225010 100064 258975
rect 100588 254969 100616 373254
rect 100850 283384 100906 283393
rect 100850 283319 100906 283328
rect 100758 282704 100814 282713
rect 100758 282639 100814 282648
rect 100772 281586 100800 282639
rect 100760 281580 100812 281586
rect 100760 281522 100812 281528
rect 100864 280158 100892 283319
rect 100852 280152 100904 280158
rect 100852 280094 100904 280100
rect 100760 278656 100812 278662
rect 100758 278624 100760 278633
rect 100812 278624 100814 278633
rect 100758 278559 100814 278568
rect 100760 277364 100812 277370
rect 100760 277306 100812 277312
rect 100772 276185 100800 277306
rect 100758 276176 100814 276185
rect 100758 276111 100814 276120
rect 100944 275324 100996 275330
rect 100944 275266 100996 275272
rect 100760 274644 100812 274650
rect 100760 274586 100812 274592
rect 100772 274553 100800 274586
rect 100852 274576 100904 274582
rect 100758 274544 100814 274553
rect 100852 274518 100904 274524
rect 100758 274479 100814 274488
rect 100864 273737 100892 274518
rect 100850 273728 100906 273737
rect 100850 273663 100906 273672
rect 100760 273216 100812 273222
rect 100760 273158 100812 273164
rect 100772 272921 100800 273158
rect 100758 272912 100814 272921
rect 100758 272847 100814 272856
rect 100760 270496 100812 270502
rect 100758 270464 100760 270473
rect 100812 270464 100814 270473
rect 100758 270399 100814 270408
rect 100956 268841 100984 275266
rect 101416 272105 101444 381482
rect 101678 281072 101734 281081
rect 101678 281007 101734 281016
rect 101692 275398 101720 281007
rect 101968 277394 101996 385630
rect 102152 369170 102180 390102
rect 103164 389230 103192 390374
rect 103578 390130 103606 390388
rect 103532 390102 103606 390130
rect 103716 390374 104144 390402
rect 104880 390374 105216 390402
rect 103152 389224 103204 389230
rect 103152 389166 103204 389172
rect 102140 369164 102192 369170
rect 102140 369106 102192 369112
rect 103532 357406 103560 390102
rect 103716 382129 103744 390374
rect 105188 386374 105216 390374
rect 106738 390416 106794 390425
rect 105322 390374 106044 390402
rect 105266 390351 105322 390360
rect 105542 388920 105598 388929
rect 105542 388855 105598 388864
rect 105176 386368 105228 386374
rect 105176 386310 105228 386316
rect 103702 382120 103758 382129
rect 103702 382055 103758 382064
rect 104254 382120 104310 382129
rect 104254 382055 104310 382064
rect 104164 370592 104216 370598
rect 104164 370534 104216 370540
rect 103520 357400 103572 357406
rect 103520 357342 103572 357348
rect 102140 354000 102192 354006
rect 102140 353942 102192 353948
rect 101876 277366 101996 277394
rect 101680 275392 101732 275398
rect 101680 275334 101732 275340
rect 101402 272096 101458 272105
rect 101402 272031 101458 272040
rect 101128 271856 101180 271862
rect 101128 271798 101180 271804
rect 101140 271289 101168 271798
rect 101126 271280 101182 271289
rect 101126 271215 101182 271224
rect 100942 268832 100998 268841
rect 100942 268767 100998 268776
rect 100760 268048 100812 268054
rect 100758 268016 100760 268025
rect 100812 268016 100814 268025
rect 100758 267951 100814 267960
rect 100760 266416 100812 266422
rect 100758 266384 100760 266393
rect 100812 266384 100814 266393
rect 100758 266319 100814 266328
rect 100758 265568 100814 265577
rect 100758 265503 100814 265512
rect 100772 264994 100800 265503
rect 100760 264988 100812 264994
rect 100760 264930 100812 264936
rect 100850 264752 100906 264761
rect 100850 264687 100906 264696
rect 100864 263634 100892 264687
rect 100944 264240 100996 264246
rect 100944 264182 100996 264188
rect 100852 263628 100904 263634
rect 100852 263570 100904 263576
rect 100760 263560 100812 263566
rect 100760 263502 100812 263508
rect 100772 263129 100800 263502
rect 100758 263120 100814 263129
rect 100758 263055 100814 263064
rect 100956 262313 100984 264182
rect 100666 262304 100722 262313
rect 100666 262239 100722 262248
rect 100942 262304 100998 262313
rect 100942 262239 100998 262248
rect 100574 254960 100630 254969
rect 100574 254895 100630 254904
rect 100114 247616 100170 247625
rect 100114 247551 100170 247560
rect 100024 225004 100076 225010
rect 100024 224946 100076 224952
rect 99472 202836 99524 202842
rect 99472 202778 99524 202784
rect 99484 202162 99512 202778
rect 99472 202156 99524 202162
rect 99472 202098 99524 202104
rect 99380 144084 99432 144090
rect 99380 144026 99432 144032
rect 98828 120352 98880 120358
rect 98828 120294 98880 120300
rect 99380 117360 99432 117366
rect 99380 117302 99432 117308
rect 99392 115938 99420 117302
rect 99380 115932 99432 115938
rect 99380 115874 99432 115880
rect 98736 111716 98788 111722
rect 98736 111658 98788 111664
rect 98736 106412 98788 106418
rect 98736 106354 98788 106360
rect 96712 97776 96764 97782
rect 96712 97718 96764 97724
rect 98644 97776 98696 97782
rect 98644 97718 98696 97724
rect 96724 96665 96752 97718
rect 97816 97300 97868 97306
rect 97816 97242 97868 97248
rect 96710 96656 96766 96665
rect 96710 96591 96766 96600
rect 97080 95328 97132 95334
rect 97078 95296 97080 95305
rect 97132 95296 97134 95305
rect 97078 95231 97134 95240
rect 97828 94489 97856 97242
rect 97906 96112 97962 96121
rect 97906 96047 97962 96056
rect 97920 95266 97948 96047
rect 97908 95260 97960 95266
rect 97908 95202 97960 95208
rect 97814 94480 97870 94489
rect 97814 94415 97870 94424
rect 97908 93832 97960 93838
rect 97908 93774 97960 93780
rect 97920 93673 97948 93774
rect 97906 93664 97962 93673
rect 97906 93599 97962 93608
rect 96710 90400 96766 90409
rect 96710 90335 96712 90344
rect 96764 90335 96766 90344
rect 97264 90364 97316 90370
rect 96712 90306 96764 90312
rect 97264 90306 97316 90312
rect 96618 83464 96674 83473
rect 96618 83399 96674 83408
rect 95332 76560 95384 76566
rect 95332 76502 95384 76508
rect 95146 75168 95202 75177
rect 95146 75103 95202 75112
rect 94504 70372 94556 70378
rect 94504 70314 94556 70320
rect 93768 57928 93820 57934
rect 93768 57870 93820 57876
rect 93768 26920 93820 26926
rect 93768 26862 93820 26868
rect 93124 20664 93176 20670
rect 93124 20606 93176 20612
rect 91008 19984 91060 19990
rect 91008 19926 91060 19932
rect 90284 6886 90404 6914
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89628 3528 89680 3534
rect 89628 3470 89680 3476
rect 89180 480 89208 3470
rect 90284 3466 90312 6886
rect 91020 3534 91048 19926
rect 93780 3534 93808 26862
rect 95056 14476 95108 14482
rect 95056 14418 95108 14424
rect 95068 3534 95096 14418
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 92756 3528 92808 3534
rect 92756 3470 92808 3476
rect 93768 3528 93820 3534
rect 93768 3470 93820 3476
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 95056 3528 95108 3534
rect 95056 3470 95108 3476
rect 90272 3460 90324 3466
rect 90272 3402 90324 3408
rect 90376 480 90404 3470
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 91572 480 91600 3402
rect 92768 480 92796 3470
rect 93964 480 93992 3470
rect 95160 480 95188 75103
rect 97276 60654 97304 90306
rect 98642 85504 98698 85513
rect 98642 85439 98698 85448
rect 98656 85241 98684 85439
rect 98642 85232 98698 85241
rect 98642 85167 98698 85176
rect 98748 74497 98776 106354
rect 98828 101448 98880 101454
rect 98828 101390 98880 101396
rect 98840 86902 98868 101390
rect 99484 101289 99512 202098
rect 100036 111926 100064 224946
rect 100128 213246 100156 247551
rect 100116 213240 100168 213246
rect 100116 213182 100168 213188
rect 100128 202842 100156 213182
rect 100116 202836 100168 202842
rect 100116 202778 100168 202784
rect 100680 117366 100708 262239
rect 100850 260672 100906 260681
rect 100850 260607 100906 260616
rect 100758 259856 100814 259865
rect 100758 259791 100814 259800
rect 100772 259554 100800 259791
rect 100760 259548 100812 259554
rect 100760 259490 100812 259496
rect 100864 259486 100892 260607
rect 100852 259480 100904 259486
rect 100852 259422 100904 259428
rect 101416 259418 101444 272031
rect 101876 271862 101904 277366
rect 101864 271856 101916 271862
rect 101864 271798 101916 271804
rect 101404 259412 101456 259418
rect 101404 259354 101456 259360
rect 100758 258224 100814 258233
rect 100758 258159 100814 258168
rect 100772 258058 100800 258159
rect 100760 258052 100812 258058
rect 100760 257994 100812 258000
rect 102048 257440 102100 257446
rect 102046 257408 102048 257417
rect 102100 257408 102102 257417
rect 102046 257343 102102 257352
rect 100758 256592 100814 256601
rect 100758 256527 100814 256536
rect 100772 255338 100800 256527
rect 100852 256012 100904 256018
rect 100852 255954 100904 255960
rect 100864 255785 100892 255954
rect 100850 255776 100906 255785
rect 100906 255734 100984 255762
rect 100850 255711 100906 255720
rect 100760 255332 100812 255338
rect 100760 255274 100812 255280
rect 100758 254960 100814 254969
rect 100758 254895 100760 254904
rect 100812 254895 100814 254904
rect 100760 254866 100812 254872
rect 100758 254144 100814 254153
rect 100758 254079 100814 254088
rect 100772 253978 100800 254079
rect 100760 253972 100812 253978
rect 100760 253914 100812 253920
rect 100758 253328 100814 253337
rect 100758 253263 100814 253272
rect 100772 252618 100800 253263
rect 100760 252612 100812 252618
rect 100760 252554 100812 252560
rect 100852 252544 100904 252550
rect 100850 252512 100852 252521
rect 100904 252512 100906 252521
rect 100850 252447 100906 252456
rect 100758 251696 100814 251705
rect 100758 251631 100814 251640
rect 100772 251394 100800 251631
rect 100760 251388 100812 251394
rect 100760 251330 100812 251336
rect 100758 250880 100814 250889
rect 100758 250815 100814 250824
rect 100772 250578 100800 250815
rect 100760 250572 100812 250578
rect 100760 250514 100812 250520
rect 100956 250458 100984 255734
rect 100772 250430 100984 250458
rect 100668 117360 100720 117366
rect 100668 117302 100720 117308
rect 100024 111920 100076 111926
rect 100024 111862 100076 111868
rect 100772 111858 100800 250430
rect 100850 250064 100906 250073
rect 100850 249999 100906 250008
rect 100864 226370 100892 249999
rect 100944 249756 100996 249762
rect 100944 249698 100996 249704
rect 100956 248441 100984 249698
rect 100942 248432 100998 248441
rect 100942 248367 100998 248376
rect 100944 247036 100996 247042
rect 100944 246978 100996 246984
rect 100956 246809 100984 246978
rect 100942 246800 100998 246809
rect 100942 246735 100998 246744
rect 101402 246256 101458 246265
rect 101402 246191 101458 246200
rect 100942 245168 100998 245177
rect 100942 245103 100998 245112
rect 100956 245002 100984 245103
rect 100944 244996 100996 245002
rect 100944 244938 100996 244944
rect 101036 244928 101088 244934
rect 101036 244870 101088 244876
rect 101048 244361 101076 244870
rect 101034 244352 101090 244361
rect 101034 244287 101090 244296
rect 100852 226364 100904 226370
rect 100852 226306 100904 226312
rect 100760 111852 100812 111858
rect 100760 111794 100812 111800
rect 100116 109744 100168 109750
rect 100116 109686 100168 109692
rect 99470 101280 99526 101289
rect 99470 101215 99526 101224
rect 100024 95328 100076 95334
rect 100024 95270 100076 95276
rect 99012 94580 99064 94586
rect 99012 94522 99064 94528
rect 99024 89690 99052 94522
rect 99012 89684 99064 89690
rect 99012 89626 99064 89632
rect 98828 86896 98880 86902
rect 98828 86838 98880 86844
rect 98734 74488 98790 74497
rect 98734 74423 98790 74432
rect 100036 66230 100064 95270
rect 100128 92177 100156 109686
rect 100298 100056 100354 100065
rect 101416 100026 101444 246191
rect 101496 218000 101548 218006
rect 101496 217942 101548 217948
rect 101508 178090 101536 217942
rect 101496 178084 101548 178090
rect 101496 178026 101548 178032
rect 101496 114028 101548 114034
rect 101496 113970 101548 113976
rect 100298 99991 100354 100000
rect 101404 100020 101456 100026
rect 100312 92313 100340 99991
rect 101404 99962 101456 99968
rect 100298 92304 100354 92313
rect 100298 92239 100354 92248
rect 100114 92168 100170 92177
rect 100114 92103 100170 92112
rect 100116 87644 100168 87650
rect 100116 87586 100168 87592
rect 100128 81326 100156 87586
rect 100116 81320 100168 81326
rect 100116 81262 100168 81268
rect 101508 77217 101536 113970
rect 101588 111104 101640 111110
rect 101588 111046 101640 111052
rect 101600 86601 101628 111046
rect 102060 110498 102088 257343
rect 102152 232558 102180 353942
rect 103428 318096 103480 318102
rect 103428 318038 103480 318044
rect 102784 281648 102836 281654
rect 102784 281590 102836 281596
rect 102232 267028 102284 267034
rect 102232 266970 102284 266976
rect 102244 261497 102272 266970
rect 102230 261488 102286 261497
rect 102230 261423 102286 261432
rect 102796 250510 102824 281590
rect 103440 281489 103468 318038
rect 103426 281480 103482 281489
rect 103426 281415 103482 281424
rect 103440 280265 103468 281415
rect 103426 280256 103482 280265
rect 103426 280191 103482 280200
rect 103428 261520 103480 261526
rect 103428 261462 103480 261468
rect 102784 250504 102836 250510
rect 102784 250446 102836 250452
rect 102324 246356 102376 246362
rect 102324 246298 102376 246304
rect 102230 242720 102286 242729
rect 102230 242655 102286 242664
rect 102140 232552 102192 232558
rect 102140 232494 102192 232500
rect 102244 208350 102272 242655
rect 102336 241398 102364 246298
rect 102324 241392 102376 241398
rect 102324 241334 102376 241340
rect 103440 240009 103468 261462
rect 104176 258058 104204 370534
rect 104268 363633 104296 382055
rect 105556 380866 105584 388855
rect 105544 380860 105596 380866
rect 105544 380802 105596 380808
rect 104254 363624 104310 363633
rect 104254 363559 104310 363568
rect 104256 322312 104308 322318
rect 104256 322254 104308 322260
rect 104268 268054 104296 322254
rect 104348 320272 104400 320278
rect 104348 320214 104400 320220
rect 104360 297430 104388 320214
rect 104438 304192 104494 304201
rect 104438 304127 104494 304136
rect 104348 297424 104400 297430
rect 104348 297366 104400 297372
rect 104348 287088 104400 287094
rect 104348 287030 104400 287036
rect 104256 268048 104308 268054
rect 104256 267990 104308 267996
rect 104360 261594 104388 287030
rect 104452 278662 104480 304127
rect 104900 291304 104952 291310
rect 104900 291246 104952 291252
rect 104440 278656 104492 278662
rect 104440 278598 104492 278604
rect 104440 263628 104492 263634
rect 104440 263570 104492 263576
rect 104348 261588 104400 261594
rect 104348 261530 104400 261536
rect 104164 258052 104216 258058
rect 104164 257994 104216 258000
rect 104256 254924 104308 254930
rect 104256 254866 104308 254872
rect 103520 251388 103572 251394
rect 103520 251330 103572 251336
rect 103426 240000 103482 240009
rect 103426 239935 103482 239944
rect 103426 238096 103482 238105
rect 103426 238031 103482 238040
rect 102232 208344 102284 208350
rect 102232 208286 102284 208292
rect 102244 207058 102272 208286
rect 102232 207052 102284 207058
rect 102232 206994 102284 207000
rect 102784 193860 102836 193866
rect 102784 193802 102836 193808
rect 102048 110492 102100 110498
rect 102048 110434 102100 110440
rect 101680 108316 101732 108322
rect 101680 108258 101732 108264
rect 101692 88233 101720 108258
rect 102796 90409 102824 193802
rect 102874 162888 102930 162897
rect 102874 162823 102930 162832
rect 102888 133890 102916 162823
rect 102966 144936 103022 144945
rect 102966 144871 103022 144880
rect 102876 133884 102928 133890
rect 102876 133826 102928 133832
rect 102980 130218 103008 144871
rect 103060 133272 103112 133278
rect 103060 133214 103112 133220
rect 102968 130212 103020 130218
rect 102968 130154 103020 130160
rect 103072 121446 103100 133214
rect 103060 121440 103112 121446
rect 103060 121382 103112 121388
rect 102782 90400 102838 90409
rect 102782 90335 102838 90344
rect 101678 88224 101734 88233
rect 101678 88159 101734 88168
rect 101586 86592 101642 86601
rect 101586 86527 101642 86536
rect 102796 82822 102824 90335
rect 102784 82816 102836 82822
rect 102784 82758 102836 82764
rect 101494 77208 101550 77217
rect 101494 77143 101550 77152
rect 100024 66224 100076 66230
rect 100024 66166 100076 66172
rect 101508 64874 101536 77143
rect 101416 64846 101536 64874
rect 97264 60648 97316 60654
rect 97264 60590 97316 60596
rect 97264 53100 97316 53106
rect 97264 53042 97316 53048
rect 96252 4888 96304 4894
rect 96252 4830 96304 4836
rect 96264 480 96292 4830
rect 97276 4826 97304 53042
rect 99288 40724 99340 40730
rect 99288 40666 99340 40672
rect 97264 4820 97316 4826
rect 97264 4762 97316 4768
rect 99300 3534 99328 40666
rect 99840 9036 99892 9042
rect 99840 8978 99892 8984
rect 98644 3528 98696 3534
rect 97446 3496 97502 3505
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 97446 3431 97502 3440
rect 97460 480 97488 3431
rect 98656 480 98684 3470
rect 99852 480 99880 8978
rect 101416 8974 101444 64846
rect 103336 54596 103388 54602
rect 103336 54538 103388 54544
rect 103348 16574 103376 54538
rect 103256 16546 103376 16574
rect 101404 8968 101456 8974
rect 101404 8910 101456 8916
rect 101036 3596 101088 3602
rect 101036 3538 101088 3544
rect 101048 480 101076 3538
rect 103256 3534 103284 16546
rect 103440 6914 103468 238031
rect 103532 218006 103560 251330
rect 104164 227044 104216 227050
rect 104164 226986 104216 226992
rect 103520 218000 103572 218006
rect 103520 217942 103572 217948
rect 103520 205012 103572 205018
rect 103520 204954 103572 204960
rect 103532 92410 103560 204954
rect 103520 92404 103572 92410
rect 103520 92346 103572 92352
rect 104176 84182 104204 226986
rect 104268 225593 104296 254866
rect 104452 244905 104480 263570
rect 104808 258868 104860 258874
rect 104808 258810 104860 258816
rect 104820 247110 104848 258810
rect 104808 247104 104860 247110
rect 104808 247046 104860 247052
rect 104438 244896 104494 244905
rect 104438 244831 104494 244840
rect 104346 241904 104402 241913
rect 104346 241839 104402 241848
rect 104254 225584 104310 225593
rect 104254 225519 104310 225528
rect 104360 217938 104388 241839
rect 104348 217932 104400 217938
rect 104348 217874 104400 217880
rect 104716 205012 104768 205018
rect 104716 204954 104768 204960
rect 104728 204406 104756 204954
rect 104716 204400 104768 204406
rect 104716 204342 104768 204348
rect 104254 182880 104310 182889
rect 104254 182815 104310 182824
rect 104164 84176 104216 84182
rect 104164 84118 104216 84124
rect 104176 84017 104204 84118
rect 104162 84008 104218 84017
rect 104162 83943 104218 83952
rect 104268 75177 104296 182815
rect 104912 151094 104940 291246
rect 104992 289876 105044 289882
rect 104992 289818 105044 289824
rect 105004 222902 105032 289818
rect 105556 229090 105584 380802
rect 106016 379506 106044 390374
rect 106338 390130 106366 390388
rect 107750 390416 107806 390425
rect 106794 390374 107516 390402
rect 107640 390374 107750 390402
rect 106738 390351 106794 390360
rect 106292 390102 106366 390130
rect 106004 379500 106056 379506
rect 106004 379442 106056 379448
rect 106188 290488 106240 290494
rect 106188 290430 106240 290436
rect 106200 289882 106228 290430
rect 106188 289876 106240 289882
rect 106188 289818 106240 289824
rect 106292 261526 106320 390102
rect 106924 377528 106976 377534
rect 106924 377470 106976 377476
rect 106280 261520 106332 261526
rect 106280 261462 106332 261468
rect 106936 250578 106964 377470
rect 107488 375358 107516 390374
rect 107948 390402 107976 390623
rect 111984 390594 112036 390600
rect 107806 390374 107884 390402
rect 107750 390351 107806 390360
rect 107764 390291 107792 390351
rect 107856 389337 107884 390374
rect 107948 390374 108376 390402
rect 109112 390374 109448 390402
rect 107842 389328 107898 389337
rect 107842 389263 107898 389272
rect 107856 389162 107884 389263
rect 107844 389156 107896 389162
rect 107844 389098 107896 389104
rect 107476 375352 107528 375358
rect 107476 375294 107528 375300
rect 107948 373994 107976 390374
rect 109420 389298 109448 390374
rect 109696 390374 109848 390402
rect 109408 389292 109460 389298
rect 109408 389234 109460 389240
rect 109696 384985 109724 390374
rect 110386 390130 110414 390388
rect 110524 390374 111136 390402
rect 111872 390374 112024 390402
rect 110386 390102 110460 390130
rect 110432 387122 110460 390102
rect 110420 387116 110472 387122
rect 110420 387058 110472 387064
rect 109682 384976 109738 384985
rect 109682 384911 109738 384920
rect 107764 373966 107976 373994
rect 107660 370524 107712 370530
rect 107660 370466 107712 370472
rect 107014 260808 107070 260817
rect 107014 260743 107070 260752
rect 106924 250572 106976 250578
rect 106924 250514 106976 250520
rect 106280 244996 106332 245002
rect 106280 244938 106332 244944
rect 105636 229764 105688 229770
rect 105636 229706 105688 229712
rect 105544 229084 105596 229090
rect 105544 229026 105596 229032
rect 105556 227118 105584 229026
rect 105544 227112 105596 227118
rect 105544 227054 105596 227060
rect 104992 222896 105044 222902
rect 104992 222838 105044 222844
rect 105544 175976 105596 175982
rect 105544 175918 105596 175924
rect 104900 151088 104952 151094
rect 104900 151030 104952 151036
rect 104806 150512 104862 150521
rect 104806 150447 104862 150456
rect 104820 145761 104848 150447
rect 104806 145752 104862 145761
rect 104806 145687 104862 145696
rect 104346 139496 104402 139505
rect 104346 139431 104402 139440
rect 104360 129062 104388 139431
rect 104348 129056 104400 129062
rect 104348 128998 104400 129004
rect 104348 91112 104400 91118
rect 104348 91054 104400 91060
rect 104254 75168 104310 75177
rect 104254 75103 104310 75112
rect 103348 6886 103468 6914
rect 102232 3528 102284 3534
rect 102232 3470 102284 3476
rect 103244 3528 103296 3534
rect 103244 3470 103296 3476
rect 102244 480 102272 3470
rect 103348 480 103376 6886
rect 104360 3466 104388 91054
rect 105450 90536 105506 90545
rect 105450 90471 105506 90480
rect 105464 89593 105492 90471
rect 105556 90370 105584 175918
rect 105648 90545 105676 229706
rect 106292 98122 106320 244938
rect 106936 237114 106964 250514
rect 107028 245002 107056 260743
rect 107016 244996 107068 245002
rect 107016 244938 107068 244944
rect 107672 238746 107700 370466
rect 107764 366450 107792 373966
rect 107752 366444 107804 366450
rect 107752 366386 107804 366392
rect 108948 335776 109000 335782
rect 108948 335718 109000 335724
rect 108396 323604 108448 323610
rect 108396 323546 108448 323552
rect 108304 320204 108356 320210
rect 108304 320146 108356 320152
rect 107660 238740 107712 238746
rect 107660 238682 107712 238688
rect 107568 238060 107620 238066
rect 107568 238002 107620 238008
rect 106924 237108 106976 237114
rect 106924 237050 106976 237056
rect 106370 210352 106426 210361
rect 106370 210287 106426 210296
rect 106384 209817 106412 210287
rect 106370 209808 106426 209817
rect 106370 209743 106426 209752
rect 106280 98116 106332 98122
rect 106280 98058 106332 98064
rect 106292 97866 106320 98058
rect 106200 97838 106320 97866
rect 105634 90536 105690 90545
rect 105634 90471 105690 90480
rect 105544 90364 105596 90370
rect 105544 90306 105596 90312
rect 105450 89584 105506 89593
rect 105450 89519 105506 89528
rect 105556 82754 105584 90306
rect 105544 82748 105596 82754
rect 105544 82690 105596 82696
rect 106200 81433 106228 97838
rect 106384 93838 106412 209743
rect 106464 181484 106516 181490
rect 106464 181426 106516 181432
rect 106372 93832 106424 93838
rect 106372 93774 106424 93780
rect 106186 81424 106242 81433
rect 106186 81359 106242 81368
rect 106476 74526 106504 181426
rect 107474 109032 107530 109041
rect 107474 108967 107530 108976
rect 107488 108390 107516 108967
rect 107476 108384 107528 108390
rect 107476 108326 107528 108332
rect 107476 93152 107528 93158
rect 107476 93094 107528 93100
rect 107488 85474 107516 93094
rect 107476 85468 107528 85474
rect 107476 85410 107528 85416
rect 106464 74520 106516 74526
rect 106464 74462 106516 74468
rect 106188 64184 106240 64190
rect 106188 64126 106240 64132
rect 106200 3466 106228 64126
rect 107580 3466 107608 238002
rect 107660 236496 107712 236502
rect 107660 236438 107712 236444
rect 107672 85377 107700 236438
rect 108316 233238 108344 320146
rect 108408 304366 108436 323546
rect 108396 304360 108448 304366
rect 108396 304302 108448 304308
rect 108396 253224 108448 253230
rect 108396 253166 108448 253172
rect 108408 237386 108436 253166
rect 108960 249762 108988 335718
rect 109040 288448 109092 288454
rect 109040 288390 109092 288396
rect 108488 249756 108540 249762
rect 108488 249698 108540 249704
rect 108948 249756 109000 249762
rect 108948 249698 109000 249704
rect 108500 249150 108528 249698
rect 108488 249144 108540 249150
rect 108488 249086 108540 249092
rect 108396 237380 108448 237386
rect 108396 237322 108448 237328
rect 108408 236502 108436 237322
rect 108396 236496 108448 236502
rect 108396 236438 108448 236444
rect 108304 233232 108356 233238
rect 108304 233174 108356 233180
rect 108948 233232 109000 233238
rect 108948 233174 109000 233180
rect 108304 224256 108356 224262
rect 108304 224198 108356 224204
rect 108316 90681 108344 224198
rect 108960 147014 108988 233174
rect 109052 160750 109080 288390
rect 109696 260817 109724 384911
rect 110524 352918 110552 390374
rect 110602 389464 110658 389473
rect 110602 389399 110658 389408
rect 110512 352912 110564 352918
rect 110512 352854 110564 352860
rect 110512 316056 110564 316062
rect 110512 315998 110564 316004
rect 109682 260808 109738 260817
rect 109682 260743 109738 260752
rect 110524 227050 110552 315998
rect 110616 238513 110644 389399
rect 111996 389094 112024 390374
rect 112088 390374 112608 390402
rect 111984 389088 112036 389094
rect 111984 389030 112036 389036
rect 112088 373994 112116 390374
rect 112732 385694 112760 418066
rect 113192 413817 113220 561682
rect 117320 560312 117372 560318
rect 117320 560254 117372 560260
rect 115202 537432 115258 537441
rect 115202 537367 115258 537376
rect 115216 463758 115244 537367
rect 115940 527876 115992 527882
rect 115940 527818 115992 527824
rect 115204 463752 115256 463758
rect 115204 463694 115256 463700
rect 113272 463004 113324 463010
rect 113272 462946 113324 462952
rect 113284 436937 113312 462946
rect 114742 442232 114798 442241
rect 114742 442167 114798 442176
rect 113270 436928 113326 436937
rect 113270 436863 113326 436872
rect 114008 433696 114060 433702
rect 114008 433638 114060 433644
rect 114020 429894 114048 433638
rect 114558 430128 114614 430137
rect 114558 430063 114614 430072
rect 114008 429888 114060 429894
rect 114008 429830 114060 429836
rect 113362 426048 113418 426057
rect 113362 425983 113418 425992
rect 113270 416800 113326 416809
rect 113270 416735 113326 416744
rect 113178 413808 113234 413817
rect 113178 413743 113234 413752
rect 113192 413030 113220 413743
rect 113180 413024 113232 413030
rect 113180 412966 113232 412972
rect 112720 385688 112772 385694
rect 112720 385630 112772 385636
rect 113180 382288 113232 382294
rect 113180 382230 113232 382236
rect 111812 373966 112116 373994
rect 111812 372570 111840 373966
rect 111800 372564 111852 372570
rect 111800 372506 111852 372512
rect 112536 372564 112588 372570
rect 112536 372506 112588 372512
rect 111064 353252 111116 353258
rect 111064 353194 111116 353200
rect 111076 352918 111104 353194
rect 111064 352912 111116 352918
rect 111064 352854 111116 352860
rect 111076 258874 111104 352854
rect 112444 338156 112496 338162
rect 112444 338098 112496 338104
rect 111064 258868 111116 258874
rect 111064 258810 111116 258816
rect 111064 253292 111116 253298
rect 111064 253234 111116 253240
rect 110602 238504 110658 238513
rect 110602 238439 110658 238448
rect 110512 227044 110564 227050
rect 110512 226986 110564 226992
rect 109684 200796 109736 200802
rect 109684 200738 109736 200744
rect 109040 160744 109092 160750
rect 109040 160686 109092 160692
rect 108488 147008 108540 147014
rect 108486 146976 108488 146985
rect 108948 147008 109000 147014
rect 108540 146976 108542 146985
rect 108948 146950 109000 146956
rect 108486 146911 108542 146920
rect 108394 143712 108450 143721
rect 108394 143647 108450 143656
rect 108408 126274 108436 143647
rect 108396 126268 108448 126274
rect 108396 126210 108448 126216
rect 108396 120760 108448 120766
rect 108396 120702 108448 120708
rect 108302 90672 108358 90681
rect 108302 90607 108358 90616
rect 108120 85468 108172 85474
rect 108120 85410 108172 85416
rect 108132 85377 108160 85410
rect 107658 85368 107714 85377
rect 107658 85303 107714 85312
rect 108118 85368 108174 85377
rect 108118 85303 108174 85312
rect 108316 81161 108344 90607
rect 108302 81152 108358 81161
rect 108302 81087 108358 81096
rect 108408 21418 108436 120702
rect 109696 118726 109724 200738
rect 109776 144968 109828 144974
rect 109776 144910 109828 144916
rect 109684 118720 109736 118726
rect 109684 118662 109736 118668
rect 108488 117360 108540 117366
rect 108488 117302 108540 117308
rect 108500 108390 108528 117302
rect 108488 108384 108540 108390
rect 108488 108326 108540 108332
rect 109696 87961 109724 118662
rect 109788 106282 109816 144910
rect 110880 133204 110932 133210
rect 110880 133146 110932 133152
rect 110892 126954 110920 133146
rect 110880 126948 110932 126954
rect 110880 126890 110932 126896
rect 110328 120828 110380 120834
rect 110328 120770 110380 120776
rect 109776 106276 109828 106282
rect 109776 106218 109828 106224
rect 109682 87952 109738 87961
rect 109682 87887 109738 87896
rect 108396 21412 108448 21418
rect 108396 21354 108448 21360
rect 110340 3466 110368 120770
rect 111076 91118 111104 253234
rect 111156 252612 111208 252618
rect 111156 252554 111208 252560
rect 111168 219337 111196 252554
rect 112456 242593 112484 338098
rect 112548 335782 112576 372506
rect 113192 370598 113220 382230
rect 113180 370592 113232 370598
rect 113180 370534 113232 370540
rect 112536 335776 112588 335782
rect 112536 335718 112588 335724
rect 112536 310480 112588 310486
rect 112536 310422 112588 310428
rect 112548 270502 112576 310422
rect 112810 278216 112866 278225
rect 112810 278151 112866 278160
rect 112824 278118 112852 278151
rect 112812 278112 112864 278118
rect 112812 278054 112864 278060
rect 112628 278044 112680 278050
rect 112628 277986 112680 277992
rect 112536 270496 112588 270502
rect 112536 270438 112588 270444
rect 112442 242584 112498 242593
rect 112442 242519 112498 242528
rect 112536 242276 112588 242282
rect 112536 242218 112588 242224
rect 111246 232520 111302 232529
rect 111246 232455 111302 232464
rect 111154 219328 111210 219337
rect 111154 219263 111210 219272
rect 111260 202842 111288 232455
rect 112548 231742 112576 242218
rect 112640 241466 112668 277986
rect 113284 269385 113312 416735
rect 113376 384305 113404 425983
rect 113546 420064 113602 420073
rect 113546 419999 113602 420008
rect 113468 402422 113496 402453
rect 113456 402416 113508 402422
rect 113454 402384 113456 402393
rect 113508 402384 113510 402393
rect 113454 402319 113510 402328
rect 113362 384296 113418 384305
rect 113362 384231 113418 384240
rect 113468 382294 113496 402319
rect 113456 382288 113508 382294
rect 113456 382230 113508 382236
rect 113560 381546 113588 419999
rect 113916 417104 113968 417110
rect 113916 417046 113968 417052
rect 113928 416809 113956 417046
rect 113914 416800 113970 416809
rect 113914 416735 113970 416744
rect 113548 381540 113600 381546
rect 113548 381482 113600 381488
rect 114468 371204 114520 371210
rect 114468 371146 114520 371152
rect 114480 370598 114508 371146
rect 114468 370592 114520 370598
rect 114468 370534 114520 370540
rect 114572 318102 114600 430063
rect 114650 417888 114706 417897
rect 114650 417823 114706 417832
rect 114560 318096 114612 318102
rect 114560 318038 114612 318044
rect 114664 310486 114692 417823
rect 114756 412634 114784 442167
rect 115020 425060 115072 425066
rect 115020 425002 115072 425008
rect 115032 424153 115060 425002
rect 115018 424144 115074 424153
rect 115018 424079 115074 424088
rect 115020 423564 115072 423570
rect 115020 423506 115072 423512
rect 115032 423065 115060 423506
rect 115018 423056 115074 423065
rect 115018 422991 115074 423000
rect 115216 421977 115244 463694
rect 115756 434716 115808 434722
rect 115756 434658 115808 434664
rect 115296 434036 115348 434042
rect 115296 433978 115348 433984
rect 115202 421968 115258 421977
rect 115202 421903 115258 421912
rect 115308 420986 115336 433978
rect 115768 433401 115796 434658
rect 115754 433392 115810 433401
rect 115754 433327 115810 433336
rect 115848 433220 115900 433226
rect 115848 433162 115900 433168
rect 115860 432313 115888 433162
rect 115846 432304 115902 432313
rect 115846 432239 115902 432248
rect 115848 431248 115900 431254
rect 115846 431216 115848 431225
rect 115900 431216 115902 431225
rect 115846 431151 115902 431160
rect 115848 428460 115900 428466
rect 115848 428402 115900 428408
rect 115860 428233 115888 428402
rect 115846 428224 115902 428233
rect 115846 428159 115902 428168
rect 115388 426284 115440 426290
rect 115388 426226 115440 426232
rect 115400 426057 115428 426226
rect 115386 426048 115442 426057
rect 115386 425983 115442 425992
rect 115388 424992 115440 424998
rect 115386 424960 115388 424969
rect 115440 424960 115442 424969
rect 115386 424895 115442 424904
rect 115296 420980 115348 420986
rect 115296 420922 115348 420928
rect 115308 412729 115336 420922
rect 115754 420880 115810 420889
rect 115754 420815 115810 420824
rect 115768 419558 115796 420815
rect 115756 419552 115808 419558
rect 115756 419494 115808 419500
rect 115952 415834 115980 527818
rect 116582 456920 116638 456929
rect 116582 456855 116638 456864
rect 116596 437073 116624 456855
rect 117332 442950 117360 560254
rect 118792 494760 118844 494766
rect 118792 494702 118844 494708
rect 117780 468512 117832 468518
rect 117780 468454 117832 468460
rect 117792 467906 117820 468454
rect 117412 467900 117464 467906
rect 117412 467842 117464 467848
rect 117780 467900 117832 467906
rect 117780 467842 117832 467848
rect 117320 442944 117372 442950
rect 117320 442886 117372 442892
rect 116582 437064 116638 437073
rect 116582 436999 116638 437008
rect 116582 434752 116638 434761
rect 116582 434687 116638 434696
rect 116596 427106 116624 434687
rect 116584 427100 116636 427106
rect 116584 427042 116636 427048
rect 117424 424998 117452 467842
rect 118698 461544 118754 461553
rect 118698 461479 118754 461488
rect 118712 461009 118740 461479
rect 118698 461000 118754 461009
rect 118698 460935 118754 460944
rect 117964 450560 118016 450566
rect 117964 450502 118016 450508
rect 117976 448497 118004 450502
rect 117962 448488 118018 448497
rect 117962 448423 118018 448432
rect 117780 442944 117832 442950
rect 117780 442886 117832 442892
rect 117502 442368 117558 442377
rect 117502 442303 117558 442312
rect 117516 425066 117544 442303
rect 117792 442270 117820 442886
rect 117780 442264 117832 442270
rect 117780 442206 117832 442212
rect 117504 425060 117556 425066
rect 117504 425002 117556 425008
rect 117412 424992 117464 424998
rect 117412 424934 117464 424940
rect 117976 417110 118004 448423
rect 118712 431254 118740 460935
rect 118700 431248 118752 431254
rect 118700 431190 118752 431196
rect 117964 417104 118016 417110
rect 117964 417046 118016 417052
rect 116124 416152 116176 416158
rect 116124 416094 116176 416100
rect 115768 415806 115980 415834
rect 115768 414882 115796 415806
rect 115846 415712 115902 415721
rect 116136 415698 116164 416094
rect 116584 416084 116636 416090
rect 116584 416026 116636 416032
rect 115902 415670 116164 415698
rect 115846 415647 115902 415656
rect 115846 414896 115902 414905
rect 115768 414854 115846 414882
rect 115846 414831 115902 414840
rect 115860 414730 115888 414831
rect 115848 414724 115900 414730
rect 115848 414666 115900 414672
rect 115294 412720 115350 412729
rect 115294 412655 115350 412664
rect 114756 412606 115244 412634
rect 114744 410644 114796 410650
rect 114744 410586 114796 410592
rect 114756 410553 114784 410586
rect 114742 410544 114798 410553
rect 114742 410479 114798 410488
rect 115216 406473 115244 412606
rect 115848 412616 115900 412622
rect 115848 412558 115900 412564
rect 115860 411641 115888 412558
rect 115846 411632 115902 411641
rect 115846 411567 115902 411576
rect 115846 408640 115902 408649
rect 115846 408575 115902 408584
rect 115860 408542 115888 408575
rect 115848 408536 115900 408542
rect 115848 408478 115900 408484
rect 115388 408400 115440 408406
rect 115388 408342 115440 408348
rect 115400 407561 115428 408342
rect 115386 407552 115442 407561
rect 115386 407487 115442 407496
rect 115202 406464 115258 406473
rect 115202 406399 115258 406408
rect 114926 405512 114982 405521
rect 114926 405447 114982 405456
rect 114940 404433 114968 405447
rect 114926 404424 114982 404433
rect 114926 404359 114982 404368
rect 114744 401124 114796 401130
rect 114744 401066 114796 401072
rect 114756 400489 114784 401066
rect 114742 400480 114798 400489
rect 114742 400415 114798 400424
rect 114940 396409 114968 404359
rect 115216 397361 115244 406399
rect 115848 405680 115900 405686
rect 115754 405648 115810 405657
rect 115848 405622 115900 405628
rect 115754 405583 115756 405592
rect 115808 405583 115810 405592
rect 115756 405554 115808 405560
rect 115860 404569 115888 405622
rect 115846 404560 115902 404569
rect 115846 404495 115902 404504
rect 115846 403472 115902 403481
rect 115846 403407 115902 403416
rect 115860 403034 115888 403407
rect 115848 403028 115900 403034
rect 115848 402970 115900 402976
rect 115570 401296 115626 401305
rect 115570 401231 115626 401240
rect 115584 400246 115612 401231
rect 115572 400240 115624 400246
rect 115572 400182 115624 400188
rect 115846 399392 115902 399401
rect 115846 399327 115902 399336
rect 115860 398886 115888 399327
rect 115848 398880 115900 398886
rect 115848 398822 115900 398828
rect 115386 398304 115442 398313
rect 115386 398239 115442 398248
rect 115400 397526 115428 398239
rect 115388 397520 115440 397526
rect 115388 397462 115440 397468
rect 115202 397352 115258 397361
rect 115202 397287 115258 397296
rect 115754 397352 115810 397361
rect 115754 397287 115810 397296
rect 115294 397216 115350 397225
rect 115294 397151 115296 397160
rect 115348 397151 115350 397160
rect 115296 397122 115348 397128
rect 114926 396400 114982 396409
rect 114926 396335 114982 396344
rect 115768 396273 115796 397287
rect 115754 396264 115810 396273
rect 115754 396199 115810 396208
rect 115768 394618 115796 396199
rect 115846 395312 115902 395321
rect 115846 395247 115902 395256
rect 115860 394738 115888 395247
rect 115848 394732 115900 394738
rect 115848 394674 115900 394680
rect 115768 394590 115888 394618
rect 115754 394224 115810 394233
rect 115754 394159 115810 394168
rect 115768 393378 115796 394159
rect 115756 393372 115808 393378
rect 115756 393314 115808 393320
rect 115570 393136 115626 393145
rect 115570 393071 115626 393080
rect 115584 392086 115612 393071
rect 115572 392080 115624 392086
rect 115572 392022 115624 392028
rect 115754 392048 115810 392057
rect 115754 391983 115756 391992
rect 115808 391983 115810 391992
rect 115756 391954 115808 391960
rect 114834 391232 114890 391241
rect 114834 391167 114890 391176
rect 114848 390794 114876 391167
rect 114836 390788 114888 390794
rect 114836 390730 114888 390736
rect 115860 329186 115888 394590
rect 116032 392080 116084 392086
rect 116032 392022 116084 392028
rect 116044 377534 116072 392022
rect 116032 377528 116084 377534
rect 116032 377470 116084 377476
rect 116136 376718 116164 415670
rect 116596 410650 116624 416026
rect 117320 413024 117372 413030
rect 117320 412966 117372 412972
rect 116584 410644 116636 410650
rect 116584 410586 116636 410592
rect 117228 403096 117280 403102
rect 117228 403038 117280 403044
rect 117240 401130 117268 403038
rect 117228 401124 117280 401130
rect 117228 401066 117280 401072
rect 117226 391096 117282 391105
rect 117226 391031 117282 391040
rect 116584 390788 116636 390794
rect 116584 390730 116636 390736
rect 116124 376712 116176 376718
rect 116124 376654 116176 376660
rect 116596 362914 116624 390730
rect 117240 390658 117268 391031
rect 117228 390652 117280 390658
rect 117228 390594 117280 390600
rect 116674 388104 116730 388113
rect 116674 388039 116730 388048
rect 116688 387433 116716 388039
rect 116674 387424 116730 387433
rect 116674 387359 116730 387368
rect 116688 364993 116716 387359
rect 116674 364984 116730 364993
rect 116674 364919 116730 364928
rect 116584 362908 116636 362914
rect 116584 362850 116636 362856
rect 115204 329180 115256 329186
rect 115204 329122 115256 329128
rect 115848 329180 115900 329186
rect 115848 329122 115900 329128
rect 114652 310480 114704 310486
rect 114652 310422 114704 310428
rect 113914 285016 113970 285025
rect 113914 284951 113970 284960
rect 113270 269376 113326 269385
rect 113270 269311 113326 269320
rect 113824 268388 113876 268394
rect 113824 268330 113876 268336
rect 113088 261520 113140 261526
rect 113088 261462 113140 261468
rect 112628 241460 112680 241466
rect 112628 241402 112680 241408
rect 112996 235340 113048 235346
rect 112996 235282 113048 235288
rect 112536 231736 112588 231742
rect 112536 231678 112588 231684
rect 111708 222896 111760 222902
rect 111708 222838 111760 222844
rect 111248 202836 111300 202842
rect 111248 202778 111300 202784
rect 111156 193860 111208 193866
rect 111156 193802 111208 193808
rect 111064 91112 111116 91118
rect 111064 91054 111116 91060
rect 111168 71058 111196 193802
rect 111156 71052 111208 71058
rect 111156 70994 111208 71000
rect 111616 21412 111668 21418
rect 111616 21354 111668 21360
rect 104348 3460 104400 3466
rect 104348 3402 104400 3408
rect 105728 3460 105780 3466
rect 105728 3402 105780 3408
rect 106188 3460 106240 3466
rect 106188 3402 106240 3408
rect 106924 3460 106976 3466
rect 106924 3402 106976 3408
rect 107568 3460 107620 3466
rect 107568 3402 107620 3408
rect 109316 3460 109368 3466
rect 109316 3402 109368 3408
rect 110328 3460 110380 3466
rect 110328 3402 110380 3408
rect 110512 3460 110564 3466
rect 110512 3402 110564 3408
rect 104530 3360 104586 3369
rect 104530 3295 104586 3304
rect 104544 480 104572 3295
rect 105740 480 105768 3402
rect 106936 480 106964 3402
rect 108120 3392 108172 3398
rect 108120 3334 108172 3340
rect 108132 480 108160 3334
rect 109328 480 109356 3402
rect 110524 480 110552 3402
rect 111628 480 111656 21354
rect 111720 3466 111748 222838
rect 111800 214600 111852 214606
rect 111800 214542 111852 214548
rect 111812 213994 111840 214542
rect 111800 213988 111852 213994
rect 111800 213930 111852 213936
rect 111812 109750 111840 213930
rect 111800 109744 111852 109750
rect 111800 109686 111852 109692
rect 112444 105392 112496 105398
rect 112444 105334 112496 105340
rect 112456 104174 112484 105334
rect 112444 104168 112496 104174
rect 112444 104110 112496 104116
rect 112456 91798 112484 104110
rect 112444 91792 112496 91798
rect 112444 91734 112496 91740
rect 112444 91044 112496 91050
rect 112444 90986 112496 90992
rect 112456 81394 112484 90986
rect 113008 87961 113036 235282
rect 112534 87952 112590 87961
rect 112534 87887 112590 87896
rect 112994 87952 113050 87961
rect 112994 87887 113050 87896
rect 112444 81388 112496 81394
rect 112444 81330 112496 81336
rect 112456 59294 112484 81330
rect 112548 80034 112576 87887
rect 112536 80028 112588 80034
rect 112536 79970 112588 79976
rect 112444 59288 112496 59294
rect 112444 59230 112496 59236
rect 113100 6914 113128 261462
rect 113836 238241 113864 268330
rect 113928 257378 113956 284951
rect 115216 267034 115244 329122
rect 115860 328574 115888 329122
rect 115848 328568 115900 328574
rect 115848 328510 115900 328516
rect 115848 310548 115900 310554
rect 115848 310490 115900 310496
rect 115204 267028 115256 267034
rect 115204 266970 115256 266976
rect 113916 257372 113968 257378
rect 113916 257314 113968 257320
rect 115296 254584 115348 254590
rect 115296 254526 115348 254532
rect 115204 253972 115256 253978
rect 115204 253914 115256 253920
rect 113916 243636 113968 243642
rect 113916 243578 113968 243584
rect 113822 238232 113878 238241
rect 113822 238167 113878 238176
rect 113272 237108 113324 237114
rect 113272 237050 113324 237056
rect 113180 226296 113232 226302
rect 113180 226238 113232 226244
rect 113192 91050 113220 226238
rect 113284 105398 113312 237050
rect 113928 226302 113956 243578
rect 113916 226296 113968 226302
rect 115216 226273 115244 253914
rect 115308 241670 115336 254526
rect 115296 241664 115348 241670
rect 115296 241606 115348 241612
rect 113916 226238 113968 226244
rect 115202 226264 115258 226273
rect 115202 226199 115258 226208
rect 114558 225584 114614 225593
rect 114558 225519 114614 225528
rect 114466 167784 114522 167793
rect 114466 167719 114522 167728
rect 113272 105392 113324 105398
rect 113272 105334 113324 105340
rect 113180 91044 113232 91050
rect 113180 90986 113232 90992
rect 112824 6886 113128 6914
rect 111708 3460 111760 3466
rect 111708 3402 111760 3408
rect 112824 480 112852 6886
rect 114480 3602 114508 167719
rect 114572 109041 114600 225519
rect 115204 204944 115256 204950
rect 115204 204886 115256 204892
rect 115216 204338 115244 204886
rect 114652 204332 114704 204338
rect 114652 204274 114704 204280
rect 115204 204332 115256 204338
rect 115204 204274 115256 204280
rect 114664 111110 114692 204274
rect 115204 124908 115256 124914
rect 115204 124850 115256 124856
rect 114652 111104 114704 111110
rect 114652 111046 114704 111052
rect 114558 109032 114614 109041
rect 114558 108967 114614 108976
rect 115216 62898 115244 124850
rect 115294 109032 115350 109041
rect 115294 108967 115350 108976
rect 115308 82822 115336 108967
rect 115296 82816 115348 82822
rect 115296 82758 115348 82764
rect 115204 62892 115256 62898
rect 115204 62834 115256 62840
rect 115860 3602 115888 310490
rect 116582 291272 116638 291281
rect 116582 291207 116638 291216
rect 116492 287768 116544 287774
rect 116492 287710 116544 287716
rect 116504 281489 116532 287710
rect 116490 281480 116546 281489
rect 116490 281415 116546 281424
rect 116596 278118 116624 291207
rect 116584 278112 116636 278118
rect 116584 278054 116636 278060
rect 115940 272536 115992 272542
rect 115940 272478 115992 272484
rect 115952 138009 115980 272478
rect 116582 236736 116638 236745
rect 116582 236671 116638 236680
rect 115938 138000 115994 138009
rect 115938 137935 115994 137944
rect 116490 138000 116546 138009
rect 116490 137935 116546 137944
rect 116504 137329 116532 137935
rect 116490 137320 116546 137329
rect 116490 137255 116546 137264
rect 116596 86737 116624 236671
rect 116688 235346 116716 364919
rect 117228 297424 117280 297430
rect 117228 297366 117280 297372
rect 117240 293962 117268 297366
rect 117228 293956 117280 293962
rect 117228 293898 117280 293904
rect 117332 266665 117360 412966
rect 118700 410576 118752 410582
rect 118700 410518 118752 410524
rect 118712 405618 118740 410518
rect 118700 405612 118752 405618
rect 118700 405554 118752 405560
rect 118804 402422 118832 494702
rect 119356 463826 119384 583743
rect 120724 497480 120776 497486
rect 120724 497422 120776 497428
rect 120736 465225 120764 497422
rect 120722 465216 120778 465225
rect 120722 465151 120778 465160
rect 119344 463820 119396 463826
rect 119344 463762 119396 463768
rect 118882 433800 118938 433809
rect 118882 433735 118938 433744
rect 118792 402416 118844 402422
rect 118792 402358 118844 402364
rect 118608 397520 118660 397526
rect 118608 397462 118660 397468
rect 118620 376038 118648 397462
rect 118608 376032 118660 376038
rect 118608 375974 118660 375980
rect 118620 373318 118648 375974
rect 118608 373312 118660 373318
rect 118608 373254 118660 373260
rect 118896 306374 118924 433735
rect 119356 426290 119384 463762
rect 120736 460934 120764 465151
rect 120736 460906 120856 460934
rect 120724 436552 120776 436558
rect 120724 436494 120776 436500
rect 120736 436150 120764 436494
rect 120724 436144 120776 436150
rect 120724 436086 120776 436092
rect 119344 426284 119396 426290
rect 119344 426226 119396 426232
rect 119344 400240 119396 400246
rect 119344 400182 119396 400188
rect 119356 316742 119384 400182
rect 119436 397180 119488 397186
rect 119436 397122 119488 397128
rect 119448 377369 119476 397122
rect 119434 377360 119490 377369
rect 119434 377295 119490 377304
rect 120736 323610 120764 436086
rect 120828 423570 120856 460906
rect 120816 423564 120868 423570
rect 120816 423506 120868 423512
rect 121472 388113 121500 585142
rect 122840 558204 122892 558210
rect 122840 558146 122892 558152
rect 121552 480956 121604 480962
rect 121552 480898 121604 480904
rect 121458 388104 121514 388113
rect 121458 388039 121514 388048
rect 121564 387802 121592 480898
rect 122748 480276 122800 480282
rect 122748 480218 122800 480224
rect 122760 476066 122788 480218
rect 122748 476060 122800 476066
rect 122748 476002 122800 476008
rect 122852 451994 122880 558146
rect 123024 476060 123076 476066
rect 123024 476002 123076 476008
rect 122840 451988 122892 451994
rect 122840 451930 122892 451936
rect 122102 451344 122158 451353
rect 122102 451279 122158 451288
rect 122116 436558 122144 451279
rect 122932 447908 122984 447914
rect 122932 447850 122984 447856
rect 122838 441688 122894 441697
rect 122838 441623 122894 441632
rect 122852 440910 122880 441623
rect 122840 440904 122892 440910
rect 122840 440846 122892 440852
rect 122104 436552 122156 436558
rect 122104 436494 122156 436500
rect 122840 428460 122892 428466
rect 122840 428402 122892 428408
rect 121644 412684 121696 412690
rect 121644 412626 121696 412632
rect 121656 408406 121684 412626
rect 121644 408400 121696 408406
rect 121644 408342 121696 408348
rect 121644 400920 121696 400926
rect 121644 400862 121696 400868
rect 121656 397526 121684 400862
rect 121644 397520 121696 397526
rect 121644 397462 121696 397468
rect 122102 388512 122158 388521
rect 122102 388447 122158 388456
rect 121552 387796 121604 387802
rect 121552 387738 121604 387744
rect 122116 382226 122144 388447
rect 122196 387796 122248 387802
rect 122196 387738 122248 387744
rect 122104 382220 122156 382226
rect 122104 382162 122156 382168
rect 122116 356697 122144 382162
rect 122208 373998 122236 387738
rect 122196 373992 122248 373998
rect 122196 373934 122248 373940
rect 122102 356688 122158 356697
rect 122102 356623 122158 356632
rect 120724 323604 120776 323610
rect 120724 323546 120776 323552
rect 119344 316736 119396 316742
rect 119344 316678 119396 316684
rect 119986 309224 120042 309233
rect 119986 309159 120042 309168
rect 118896 306346 119384 306374
rect 119356 292641 119384 306346
rect 119342 292632 119398 292641
rect 119342 292567 119398 292576
rect 119356 282878 119384 292567
rect 119344 282872 119396 282878
rect 119344 282814 119396 282820
rect 119344 280900 119396 280906
rect 119344 280842 119396 280848
rect 117318 266656 117374 266665
rect 117318 266591 117374 266600
rect 117332 266082 117360 266591
rect 117320 266076 117372 266082
rect 117320 266018 117372 266024
rect 117964 261588 118016 261594
rect 117964 261530 118016 261536
rect 116768 251932 116820 251938
rect 116768 251874 116820 251880
rect 116780 235929 116808 251874
rect 116766 235920 116822 235929
rect 116766 235855 116822 235864
rect 116676 235340 116728 235346
rect 116676 235282 116728 235288
rect 117228 199436 117280 199442
rect 117228 199378 117280 199384
rect 116674 149696 116730 149705
rect 116674 149631 116730 149640
rect 116688 117337 116716 149631
rect 116674 117328 116730 117337
rect 116674 117263 116730 117272
rect 116582 86728 116638 86737
rect 116582 86663 116638 86672
rect 117240 3602 117268 199378
rect 117976 175302 118004 261530
rect 119356 252550 119384 280842
rect 119344 252544 119396 252550
rect 119344 252486 119396 252492
rect 118700 227112 118752 227118
rect 118700 227054 118752 227060
rect 118608 220108 118660 220114
rect 118608 220050 118660 220056
rect 117964 175296 118016 175302
rect 117964 175238 118016 175244
rect 117976 138825 118004 175238
rect 117962 138816 118018 138825
rect 117962 138751 118018 138760
rect 118620 3602 118648 220050
rect 118712 89622 118740 227054
rect 118790 191040 118846 191049
rect 118790 190975 118846 190984
rect 118700 89616 118752 89622
rect 118700 89558 118752 89564
rect 118804 64870 118832 190975
rect 118792 64864 118844 64870
rect 118792 64806 118844 64812
rect 119896 46300 119948 46306
rect 119896 46242 119948 46248
rect 119908 16574 119936 46242
rect 119816 16546 119936 16574
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 114468 3596 114520 3602
rect 114468 3538 114520 3544
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 115848 3596 115900 3602
rect 115848 3538 115900 3544
rect 116400 3596 116452 3602
rect 116400 3538 116452 3544
rect 117228 3596 117280 3602
rect 117228 3538 117280 3544
rect 117596 3596 117648 3602
rect 117596 3538 117648 3544
rect 118608 3596 118660 3602
rect 118608 3538 118660 3544
rect 114020 480 114048 3538
rect 115216 480 115244 3538
rect 116412 480 116440 3538
rect 117608 480 117636 3538
rect 119816 3058 119844 16546
rect 120000 6914 120028 309159
rect 120814 291816 120870 291825
rect 120814 291751 120870 291760
rect 120722 287192 120778 287201
rect 120722 287127 120778 287136
rect 120736 229770 120764 287127
rect 120828 249082 120856 291751
rect 120816 249076 120868 249082
rect 120816 249018 120868 249024
rect 122116 236745 122144 356623
rect 122194 331392 122250 331401
rect 122194 331327 122250 331336
rect 122208 253298 122236 331327
rect 122746 309360 122802 309369
rect 122746 309295 122802 309304
rect 122196 253292 122248 253298
rect 122196 253234 122248 253240
rect 122102 236736 122158 236745
rect 122102 236671 122158 236680
rect 122196 236700 122248 236706
rect 122196 236642 122248 236648
rect 120724 229764 120776 229770
rect 120724 229706 120776 229712
rect 121368 224256 121420 224262
rect 121368 224198 121420 224204
rect 120080 178696 120132 178702
rect 120080 178638 120132 178644
rect 120092 100065 120120 178638
rect 120078 100056 120134 100065
rect 120078 99991 120134 100000
rect 121380 6914 121408 224198
rect 122208 220794 122236 236642
rect 121460 220788 121512 220794
rect 121460 220730 121512 220736
rect 122196 220788 122248 220794
rect 122196 220730 122248 220736
rect 121472 88330 121500 220730
rect 121552 184204 121604 184210
rect 121552 184146 121604 184152
rect 121460 88324 121512 88330
rect 121460 88266 121512 88272
rect 121472 88097 121500 88266
rect 121458 88088 121514 88097
rect 121458 88023 121514 88032
rect 121564 77246 121592 184146
rect 121552 77240 121604 77246
rect 121552 77182 121604 77188
rect 121564 76498 121592 77182
rect 121552 76492 121604 76498
rect 121552 76434 121604 76440
rect 122104 76492 122156 76498
rect 122104 76434 122156 76440
rect 122116 63442 122144 76434
rect 122104 63436 122156 63442
rect 122104 63378 122156 63384
rect 119908 6886 120028 6914
rect 121104 6886 121408 6914
rect 118792 3052 118844 3058
rect 118792 2994 118844 3000
rect 119804 3052 119856 3058
rect 119804 2994 119856 3000
rect 118804 480 118832 2994
rect 119908 480 119936 6886
rect 121104 480 121132 6886
rect 122760 3602 122788 309295
rect 122852 304201 122880 428402
rect 122944 376650 122972 447850
rect 123036 428466 123064 476002
rect 123496 469266 123524 586502
rect 123484 469260 123536 469266
rect 123484 469202 123536 469208
rect 123496 433226 123524 469202
rect 124128 451988 124180 451994
rect 124128 451930 124180 451936
rect 124140 451897 124168 451930
rect 124126 451888 124182 451897
rect 124126 451823 124182 451832
rect 123484 433220 123536 433226
rect 123484 433162 123536 433168
rect 123024 428460 123076 428466
rect 123024 428402 123076 428408
rect 123484 418804 123536 418810
rect 123484 418746 123536 418752
rect 123496 412622 123524 418746
rect 123484 412616 123536 412622
rect 123484 412558 123536 412564
rect 124232 384985 124260 589290
rect 128360 588600 128412 588606
rect 128360 588542 128412 588548
rect 125600 576156 125652 576162
rect 125600 576098 125652 576104
rect 124312 478168 124364 478174
rect 124312 478110 124364 478116
rect 124324 386374 124352 478110
rect 125508 409148 125560 409154
rect 125508 409090 125560 409096
rect 125520 405686 125548 409090
rect 125508 405680 125560 405686
rect 125508 405622 125560 405628
rect 125612 388521 125640 576098
rect 126980 573368 127032 573374
rect 126980 573310 127032 573316
rect 125692 542428 125744 542434
rect 125692 542370 125744 542376
rect 125704 442134 125732 542370
rect 125692 442128 125744 442134
rect 125692 442070 125744 442076
rect 126244 442128 126296 442134
rect 126244 442070 126296 442076
rect 125704 441658 125732 442070
rect 125692 441652 125744 441658
rect 125692 441594 125744 441600
rect 126256 422958 126284 442070
rect 126336 425740 126388 425746
rect 126336 425682 126388 425688
rect 126244 422952 126296 422958
rect 126244 422894 126296 422900
rect 126348 416158 126376 425682
rect 126336 416152 126388 416158
rect 126336 416094 126388 416100
rect 125692 414724 125744 414730
rect 125692 414666 125744 414672
rect 125598 388512 125654 388521
rect 125598 388447 125654 388456
rect 124312 386368 124364 386374
rect 124312 386310 124364 386316
rect 124864 386368 124916 386374
rect 124864 386310 124916 386316
rect 124218 384976 124274 384985
rect 124218 384911 124274 384920
rect 122932 376644 122984 376650
rect 122932 376586 122984 376592
rect 123484 376644 123536 376650
rect 123484 376586 123536 376592
rect 123496 361486 123524 376586
rect 123484 361480 123536 361486
rect 123484 361422 123536 361428
rect 124220 359576 124272 359582
rect 124220 359518 124272 359524
rect 123576 346520 123628 346526
rect 123576 346462 123628 346468
rect 123484 304360 123536 304366
rect 123484 304302 123536 304308
rect 122838 304192 122894 304201
rect 122838 304127 122894 304136
rect 123496 277370 123524 304302
rect 123484 277364 123536 277370
rect 123484 277306 123536 277312
rect 123484 266076 123536 266082
rect 123484 266018 123536 266024
rect 122840 206304 122892 206310
rect 122840 206246 122892 206252
rect 122852 92546 122880 206246
rect 123496 164354 123524 266018
rect 123588 253230 123616 346462
rect 124126 306912 124182 306921
rect 124126 306847 124182 306856
rect 123576 253224 123628 253230
rect 123576 253166 123628 253172
rect 123760 206304 123812 206310
rect 123760 206246 123812 206252
rect 123772 205698 123800 206246
rect 123760 205692 123812 205698
rect 123760 205634 123812 205640
rect 123484 164348 123536 164354
rect 123484 164290 123536 164296
rect 123496 120086 123524 164290
rect 123484 120080 123536 120086
rect 123484 120022 123536 120028
rect 123484 109064 123536 109070
rect 123484 109006 123536 109012
rect 122840 92540 122892 92546
rect 122840 92482 122892 92488
rect 123496 77081 123524 109006
rect 123482 77072 123538 77081
rect 123482 77007 123538 77016
rect 122288 3596 122340 3602
rect 122288 3538 122340 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 122300 480 122328 3538
rect 124140 3534 124168 306847
rect 124232 236706 124260 359518
rect 124876 358737 124904 386310
rect 125048 359576 125100 359582
rect 125048 359518 125100 359524
rect 125060 358834 125088 359518
rect 125048 358828 125100 358834
rect 125048 358770 125100 358776
rect 124862 358728 124918 358737
rect 124862 358663 124918 358672
rect 124864 338224 124916 338230
rect 124864 338166 124916 338172
rect 124220 236700 124272 236706
rect 124220 236642 124272 236648
rect 124876 120766 124904 338166
rect 125704 322930 125732 414666
rect 126992 387818 127020 573310
rect 128372 400926 128400 588542
rect 129738 581088 129794 581097
rect 129738 581023 129794 581032
rect 129004 554804 129056 554810
rect 129004 554746 129056 554752
rect 128360 400920 128412 400926
rect 128360 400862 128412 400868
rect 129016 387841 129044 554746
rect 126900 387790 127020 387818
rect 128358 387832 128414 387841
rect 126900 384946 126928 387790
rect 128358 387767 128414 387776
rect 129002 387832 129058 387841
rect 129002 387767 129058 387776
rect 128372 386345 128400 387767
rect 129752 387705 129780 581023
rect 134524 578264 134576 578270
rect 134524 578206 134576 578212
rect 132592 576904 132644 576910
rect 132592 576846 132644 576852
rect 130384 541000 130436 541006
rect 130384 540942 130436 540948
rect 129832 419552 129884 419558
rect 129832 419494 129884 419500
rect 129738 387696 129794 387705
rect 129738 387631 129794 387640
rect 128358 386336 128414 386345
rect 128358 386271 128414 386280
rect 126888 384940 126940 384946
rect 126888 384882 126940 384888
rect 126900 382226 126928 384882
rect 128360 382968 128412 382974
rect 128360 382910 128412 382916
rect 128372 382294 128400 382910
rect 128360 382288 128412 382294
rect 128360 382230 128412 382236
rect 126888 382220 126940 382226
rect 126888 382162 126940 382168
rect 127622 330032 127678 330041
rect 127622 329967 127678 329976
rect 126334 327176 126390 327185
rect 126334 327111 126390 327120
rect 125692 322924 125744 322930
rect 125692 322866 125744 322872
rect 125704 322318 125732 322866
rect 125692 322312 125744 322318
rect 125692 322254 125744 322260
rect 126242 305008 126298 305017
rect 126242 304943 126298 304952
rect 124956 300144 125008 300150
rect 124956 300086 125008 300092
rect 124968 289241 124996 300086
rect 124954 289232 125010 289241
rect 124954 289167 125010 289176
rect 124956 282872 125008 282878
rect 124956 282814 125008 282820
rect 124968 261594 124996 282814
rect 124956 261588 125008 261594
rect 124956 261530 125008 261536
rect 125508 236700 125560 236706
rect 125508 236642 125560 236648
rect 125416 233912 125468 233918
rect 125416 233854 125468 233860
rect 124864 120760 124916 120766
rect 124864 120702 124916 120708
rect 124864 89752 124916 89758
rect 124864 89694 124916 89700
rect 124876 82793 124904 89694
rect 125428 89622 125456 233854
rect 125416 89616 125468 89622
rect 125416 89558 125468 89564
rect 125428 87650 125456 89558
rect 125416 87644 125468 87650
rect 125416 87586 125468 87592
rect 124862 82784 124918 82793
rect 124862 82719 124918 82728
rect 124876 71670 124904 82719
rect 124864 71664 124916 71670
rect 124864 71606 124916 71612
rect 125520 3534 125548 236642
rect 125600 198008 125652 198014
rect 125600 197950 125652 197956
rect 125612 89758 125640 197950
rect 125600 89752 125652 89758
rect 125600 89694 125652 89700
rect 125600 36576 125652 36582
rect 125600 36518 125652 36524
rect 125612 16574 125640 36518
rect 125612 16546 125916 16574
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125888 480 125916 16546
rect 126256 3602 126284 304943
rect 126348 199442 126376 327111
rect 126888 320884 126940 320890
rect 126888 320826 126940 320832
rect 126900 320278 126928 320826
rect 126888 320272 126940 320278
rect 126888 320214 126940 320220
rect 126336 199436 126388 199442
rect 126336 199378 126388 199384
rect 126900 150482 126928 320214
rect 126888 150476 126940 150482
rect 126888 150418 126940 150424
rect 126900 146266 126928 150418
rect 126888 146260 126940 146266
rect 126888 146202 126940 146208
rect 126336 126336 126388 126342
rect 126336 126278 126388 126284
rect 126348 64190 126376 126278
rect 127636 124914 127664 329967
rect 127716 291236 127768 291242
rect 127716 291178 127768 291184
rect 127728 287026 127756 291178
rect 127716 287020 127768 287026
rect 127716 286962 127768 286968
rect 127728 158846 127756 286962
rect 128372 233918 128400 382230
rect 129004 367872 129056 367878
rect 129004 367814 129056 367820
rect 129016 356046 129044 367814
rect 129004 356040 129056 356046
rect 129004 355982 129056 355988
rect 129002 336832 129058 336841
rect 129002 336767 129058 336776
rect 128728 271856 128780 271862
rect 128728 271798 128780 271804
rect 128740 271250 128768 271798
rect 128728 271244 128780 271250
rect 128728 271186 128780 271192
rect 128360 233912 128412 233918
rect 128360 233854 128412 233860
rect 128358 231160 128414 231169
rect 128358 231095 128414 231104
rect 127716 158840 127768 158846
rect 127716 158782 127768 158788
rect 127806 158808 127862 158817
rect 127728 158030 127756 158782
rect 127806 158743 127862 158752
rect 127716 158024 127768 158030
rect 127716 157966 127768 157972
rect 127716 129940 127768 129946
rect 127716 129882 127768 129888
rect 127624 124908 127676 124914
rect 127624 124850 127676 124856
rect 126336 64184 126388 64190
rect 126336 64126 126388 64132
rect 127728 21418 127756 129882
rect 127820 128314 127848 158743
rect 127808 128308 127860 128314
rect 127808 128250 127860 128256
rect 127716 21412 127768 21418
rect 127716 21354 127768 21360
rect 128372 6914 128400 231095
rect 129016 46238 129044 336767
rect 129646 297528 129702 297537
rect 129646 297463 129702 297472
rect 129660 271250 129688 297463
rect 129844 277394 129872 419494
rect 130396 408474 130424 540942
rect 131120 483676 131172 483682
rect 131120 483618 131172 483624
rect 131132 410582 131160 483618
rect 132498 435296 132554 435305
rect 132498 435231 132554 435240
rect 131120 410576 131172 410582
rect 131120 410518 131172 410524
rect 130384 408468 130436 408474
rect 130384 408410 130436 408416
rect 130396 378049 130424 408410
rect 131764 393440 131816 393446
rect 131764 393382 131816 393388
rect 131776 392086 131804 393382
rect 131764 392080 131816 392086
rect 131764 392022 131816 392028
rect 130474 387696 130530 387705
rect 130474 387631 130530 387640
rect 130382 378040 130438 378049
rect 130382 377975 130438 377984
rect 130488 368490 130516 387631
rect 131776 386374 131804 392022
rect 131764 386368 131816 386374
rect 131764 386310 131816 386316
rect 130476 368484 130528 368490
rect 130476 368426 130528 368432
rect 130476 340944 130528 340950
rect 130476 340886 130528 340892
rect 130382 305144 130438 305153
rect 130382 305079 130438 305088
rect 129752 277366 129872 277394
rect 129752 273222 129780 277366
rect 129740 273216 129792 273222
rect 129740 273158 129792 273164
rect 129752 272542 129780 273158
rect 129740 272536 129792 272542
rect 129740 272478 129792 272484
rect 129648 271244 129700 271250
rect 129648 271186 129700 271192
rect 129188 251864 129240 251870
rect 129188 251806 129240 251812
rect 129096 249144 129148 249150
rect 129096 249086 129148 249092
rect 129108 102134 129136 249086
rect 129200 242457 129228 251806
rect 129186 242448 129242 242457
rect 129186 242383 129242 242392
rect 129740 209092 129792 209098
rect 129740 209034 129792 209040
rect 129752 208418 129780 209034
rect 129740 208412 129792 208418
rect 129740 208354 129792 208360
rect 129096 102128 129148 102134
rect 129096 102070 129148 102076
rect 129108 101522 129136 102070
rect 129096 101516 129148 101522
rect 129096 101458 129148 101464
rect 129752 97306 129780 208354
rect 129740 97300 129792 97306
rect 129740 97242 129792 97248
rect 129004 46232 129056 46238
rect 129004 46174 129056 46180
rect 128280 6886 128400 6914
rect 126244 3596 126296 3602
rect 126244 3538 126296 3544
rect 128280 3534 128308 6886
rect 128268 3528 128320 3534
rect 128268 3470 128320 3476
rect 129372 3528 129424 3534
rect 130396 3505 130424 305079
rect 130488 298790 130516 340886
rect 131854 305280 131910 305289
rect 131854 305215 131910 305224
rect 130476 298784 130528 298790
rect 130476 298726 130528 298732
rect 130568 296064 130620 296070
rect 130568 296006 130620 296012
rect 130476 265668 130528 265674
rect 130476 265610 130528 265616
rect 130488 195294 130516 265610
rect 130580 257446 130608 296006
rect 131764 264308 131816 264314
rect 131764 264250 131816 264256
rect 130658 263664 130714 263673
rect 130658 263599 130714 263608
rect 130568 257440 130620 257446
rect 130568 257382 130620 257388
rect 130672 254561 130700 263599
rect 130658 254552 130714 254561
rect 130658 254487 130714 254496
rect 130476 195288 130528 195294
rect 130476 195230 130528 195236
rect 130476 104168 130528 104174
rect 130476 104110 130528 104116
rect 130488 62830 130516 104110
rect 130476 62824 130528 62830
rect 130476 62766 130528 62772
rect 131776 11762 131804 264250
rect 131868 226953 131896 305215
rect 131854 226944 131910 226953
rect 131854 226879 131910 226888
rect 131856 150544 131908 150550
rect 131856 150486 131908 150492
rect 131868 120766 131896 150486
rect 131856 120760 131908 120766
rect 131856 120702 131908 120708
rect 132512 16574 132540 435231
rect 132604 393446 132632 576846
rect 133880 493332 133932 493338
rect 133880 493274 133932 493280
rect 133142 450120 133198 450129
rect 133142 450055 133198 450064
rect 133156 437481 133184 450055
rect 133142 437472 133198 437481
rect 133142 437407 133198 437416
rect 132592 393440 132644 393446
rect 132592 393382 132644 393388
rect 133892 389094 133920 493274
rect 133880 389088 133932 389094
rect 133880 389030 133932 389036
rect 133142 325952 133198 325961
rect 133142 325887 133198 325896
rect 133156 129946 133184 325887
rect 133326 281616 133382 281625
rect 133326 281551 133382 281560
rect 133236 221536 133288 221542
rect 133236 221478 133288 221484
rect 133144 129940 133196 129946
rect 133144 129882 133196 129888
rect 133248 54602 133276 221478
rect 133340 220833 133368 281551
rect 133880 247104 133932 247110
rect 133880 247046 133932 247052
rect 133326 220824 133382 220833
rect 133326 220759 133382 220768
rect 133892 99498 133920 247046
rect 133800 99470 133920 99498
rect 133800 99414 133828 99470
rect 133788 99408 133840 99414
rect 133788 99350 133840 99356
rect 133800 77246 133828 99350
rect 133788 77240 133840 77246
rect 133788 77182 133840 77188
rect 133236 54596 133288 54602
rect 133236 54538 133288 54544
rect 132512 16546 133000 16574
rect 131764 11756 131816 11762
rect 131764 11698 131816 11704
rect 129372 3470 129424 3476
rect 130382 3496 130438 3505
rect 129384 480 129412 3470
rect 130382 3431 130438 3440
rect 132972 480 133000 16546
rect 134536 4214 134564 578206
rect 136652 536761 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702778 154160 703520
rect 154120 702772 154172 702778
rect 154120 702714 154172 702720
rect 170324 702574 170352 703520
rect 191748 703452 191800 703458
rect 191748 703394 191800 703400
rect 177304 702840 177356 702846
rect 177304 702782 177356 702788
rect 170312 702568 170364 702574
rect 170312 702510 170364 702516
rect 143540 592680 143592 592686
rect 143540 592622 143592 592628
rect 141424 579692 141476 579698
rect 141424 579634 141476 579640
rect 136638 536752 136694 536761
rect 136638 536687 136694 536696
rect 136732 525088 136784 525094
rect 136732 525030 136784 525036
rect 136640 436756 136692 436762
rect 136640 436698 136692 436704
rect 136652 435470 136680 436698
rect 136640 435464 136692 435470
rect 136640 435406 136692 435412
rect 135994 347848 136050 347857
rect 135994 347783 136050 347792
rect 134614 317656 134670 317665
rect 134614 317591 134670 317600
rect 134628 79354 134656 317591
rect 135904 282192 135956 282198
rect 135904 282134 135956 282140
rect 134708 268456 134760 268462
rect 134708 268398 134760 268404
rect 134720 242214 134748 268398
rect 135168 247716 135220 247722
rect 135168 247658 135220 247664
rect 135180 247110 135208 247658
rect 135168 247104 135220 247110
rect 135168 247046 135220 247052
rect 134708 242208 134760 242214
rect 134708 242150 134760 242156
rect 134616 79348 134668 79354
rect 134616 79290 134668 79296
rect 135916 25566 135944 282134
rect 136008 274582 136036 347783
rect 136652 320890 136680 435406
rect 136744 418810 136772 525030
rect 141436 459678 141464 579634
rect 142158 538792 142214 538801
rect 142158 538727 142214 538736
rect 142068 466472 142120 466478
rect 142068 466414 142120 466420
rect 141424 459672 141476 459678
rect 141424 459614 141476 459620
rect 141436 425746 141464 459614
rect 141424 425740 141476 425746
rect 141424 425682 141476 425688
rect 136732 418804 136784 418810
rect 136732 418746 136784 418752
rect 137468 369164 137520 369170
rect 137468 369106 137520 369112
rect 136640 320884 136692 320890
rect 136640 320826 136692 320832
rect 137284 305040 137336 305046
rect 137284 304982 137336 304988
rect 136088 275392 136140 275398
rect 136088 275334 136140 275340
rect 135996 274576 136048 274582
rect 135996 274518 136048 274524
rect 135996 271244 136048 271250
rect 135996 271186 136048 271192
rect 136008 167074 136036 271186
rect 136100 240854 136128 275334
rect 136088 240848 136140 240854
rect 136088 240790 136140 240796
rect 135996 167068 136048 167074
rect 135996 167010 136048 167016
rect 136008 124098 136036 167010
rect 135996 124092 136048 124098
rect 135996 124034 136048 124040
rect 135904 25560 135956 25566
rect 135904 25502 135956 25508
rect 134524 4208 134576 4214
rect 134524 4150 134576 4156
rect 136456 4208 136508 4214
rect 136456 4150 136508 4156
rect 136468 480 136496 4150
rect 137296 3466 137324 304982
rect 137376 271244 137428 271250
rect 137376 271186 137428 271192
rect 137388 42090 137416 271186
rect 137480 255270 137508 369106
rect 141608 345160 141660 345166
rect 141608 345102 141660 345108
rect 141424 343732 141476 343738
rect 141424 343674 141476 343680
rect 140134 324456 140190 324465
rect 140134 324391 140190 324400
rect 138754 299024 138810 299033
rect 138754 298959 138810 298968
rect 138020 293956 138072 293962
rect 138020 293898 138072 293904
rect 138032 290562 138060 293898
rect 138020 290556 138072 290562
rect 138020 290498 138072 290504
rect 137468 255264 137520 255270
rect 137468 255206 137520 255212
rect 137480 254590 137508 255206
rect 137468 254584 137520 254590
rect 137468 254526 137520 254532
rect 138664 253224 138716 253230
rect 138664 253166 138716 253172
rect 137376 42084 137428 42090
rect 137376 42026 137428 42032
rect 138676 24138 138704 253166
rect 138768 192506 138796 298959
rect 140044 285048 140096 285054
rect 140044 284990 140096 284996
rect 138848 264988 138900 264994
rect 138848 264930 138900 264936
rect 138860 231130 138888 264930
rect 138848 231124 138900 231130
rect 138848 231066 138900 231072
rect 138756 192500 138808 192506
rect 138756 192442 138808 192448
rect 140056 33794 140084 284990
rect 140148 243642 140176 324391
rect 141436 319462 141464 343674
rect 141424 319456 141476 319462
rect 141424 319398 141476 319404
rect 141422 308000 141478 308009
rect 141422 307935 141478 307944
rect 140136 243636 140188 243642
rect 140136 243578 140188 243584
rect 140044 33788 140096 33794
rect 140044 33730 140096 33736
rect 138664 24132 138716 24138
rect 138664 24074 138716 24080
rect 141436 19990 141464 307935
rect 141514 293176 141570 293185
rect 141514 293111 141570 293120
rect 141528 53106 141556 293111
rect 141620 126342 141648 345102
rect 142080 343738 142108 466414
rect 142172 416090 142200 538727
rect 142804 465112 142856 465118
rect 142804 465054 142856 465060
rect 142816 443698 142844 465054
rect 142804 443692 142856 443698
rect 142804 443634 142856 443640
rect 142160 416084 142212 416090
rect 142160 416026 142212 416032
rect 142160 414044 142212 414050
rect 142160 413986 142212 413992
rect 142172 408474 142200 413986
rect 142160 408468 142212 408474
rect 142160 408410 142212 408416
rect 142068 343732 142120 343738
rect 142068 343674 142120 343680
rect 141700 327140 141752 327146
rect 141700 327082 141752 327088
rect 141712 293282 141740 327082
rect 142816 317490 142844 443634
rect 143552 409154 143580 592622
rect 147680 530664 147732 530670
rect 147680 530606 147732 530612
rect 147586 454200 147642 454209
rect 147586 454135 147642 454144
rect 143632 429888 143684 429894
rect 143632 429830 143684 429836
rect 143540 409148 143592 409154
rect 143540 409090 143592 409096
rect 142988 346452 143040 346458
rect 142988 346394 143040 346400
rect 142804 317484 142856 317490
rect 142804 317426 142856 317432
rect 142816 316034 142844 317426
rect 142816 316006 142936 316034
rect 142802 314936 142858 314945
rect 142802 314871 142858 314880
rect 141700 293276 141752 293282
rect 141700 293218 141752 293224
rect 141608 126336 141660 126342
rect 141608 126278 141660 126284
rect 141516 53100 141568 53106
rect 141516 53042 141568 53048
rect 141424 19984 141476 19990
rect 141424 19926 141476 19932
rect 142816 13122 142844 314871
rect 142908 287026 142936 316006
rect 142896 287020 142948 287026
rect 142896 286962 142948 286968
rect 142894 282160 142950 282169
rect 142894 282095 142950 282104
rect 142908 50386 142936 282095
rect 143000 120834 143028 346394
rect 143644 293962 143672 429830
rect 145656 334008 145708 334014
rect 145656 333950 145708 333956
rect 144276 323672 144328 323678
rect 144276 323614 144328 323620
rect 143632 293956 143684 293962
rect 143632 293898 143684 293904
rect 144184 278112 144236 278118
rect 144184 278054 144236 278060
rect 142988 120828 143040 120834
rect 142988 120770 143040 120776
rect 144196 51746 144224 278054
rect 144288 227633 144316 323614
rect 144828 317552 144880 317558
rect 144828 317494 144880 317500
rect 144274 227624 144330 227633
rect 144274 227559 144330 227568
rect 144184 51740 144236 51746
rect 144184 51682 144236 51688
rect 142896 50380 142948 50386
rect 142896 50322 142948 50328
rect 142804 13116 142856 13122
rect 142804 13058 142856 13064
rect 144840 3534 144868 317494
rect 145564 268456 145616 268462
rect 145564 268398 145616 268404
rect 145576 54534 145604 268398
rect 145668 263566 145696 333950
rect 147034 328536 147090 328545
rect 147034 328471 147090 328480
rect 145748 273964 145800 273970
rect 145748 273906 145800 273912
rect 145656 263560 145708 263566
rect 145656 263502 145708 263508
rect 145760 242282 145788 273906
rect 146944 272604 146996 272610
rect 146944 272546 146996 272552
rect 145748 242276 145800 242282
rect 145748 242218 145800 242224
rect 145656 172644 145708 172650
rect 145656 172586 145708 172592
rect 145668 140049 145696 172586
rect 145654 140040 145710 140049
rect 145654 139975 145710 139984
rect 145564 54528 145616 54534
rect 145564 54470 145616 54476
rect 146956 43450 146984 272546
rect 147048 265674 147076 328471
rect 147128 266416 147180 266422
rect 147128 266358 147180 266364
rect 147036 265668 147088 265674
rect 147036 265610 147088 265616
rect 147140 218754 147168 266358
rect 147128 218748 147180 218754
rect 147128 218690 147180 218696
rect 147036 161492 147088 161498
rect 147036 161434 147088 161440
rect 147048 124166 147076 161434
rect 147036 124160 147088 124166
rect 147036 124102 147088 124108
rect 146944 43444 146996 43450
rect 146944 43386 146996 43392
rect 147600 3534 147628 454135
rect 147692 403782 147720 530606
rect 155776 470620 155828 470626
rect 155776 470562 155828 470568
rect 151084 449948 151136 449954
rect 151084 449890 151136 449896
rect 151096 426426 151124 449890
rect 152464 445868 152516 445874
rect 152464 445810 152516 445816
rect 152476 431254 152504 445810
rect 152464 431248 152516 431254
rect 152464 431190 152516 431196
rect 151084 426420 151136 426426
rect 151084 426362 151136 426368
rect 148324 412684 148376 412690
rect 148324 412626 148376 412632
rect 147680 403776 147732 403782
rect 147680 403718 147732 403724
rect 147692 403102 147720 403718
rect 147680 403096 147732 403102
rect 147680 403038 147732 403044
rect 148336 384946 148364 412626
rect 151082 410136 151138 410145
rect 151082 410071 151138 410080
rect 148416 403776 148468 403782
rect 148416 403718 148468 403724
rect 148324 384940 148376 384946
rect 148324 384882 148376 384888
rect 148428 376009 148456 403718
rect 148968 384940 149020 384946
rect 148968 384882 149020 384888
rect 148414 376000 148470 376009
rect 148414 375935 148470 375944
rect 148414 342272 148470 342281
rect 148414 342207 148470 342216
rect 148324 307828 148376 307834
rect 148324 307770 148376 307776
rect 147680 264920 147732 264926
rect 147680 264862 147732 264868
rect 147692 264246 147720 264862
rect 147680 264240 147732 264246
rect 147680 264182 147732 264188
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147588 3528 147640 3534
rect 147588 3470 147640 3476
rect 137284 3460 137336 3466
rect 137284 3402 137336 3408
rect 140044 2100 140096 2106
rect 140044 2042 140096 2048
rect 140056 480 140084 2042
rect 143552 480 143580 3470
rect 147140 480 147168 3470
rect 148336 3369 148364 307770
rect 148428 221542 148456 342207
rect 148508 276072 148560 276078
rect 148508 276014 148560 276020
rect 148520 249150 148548 276014
rect 148980 264926 149008 384882
rect 151096 378049 151124 410071
rect 152464 408536 152516 408542
rect 152464 408478 152516 408484
rect 151176 393372 151228 393378
rect 151176 393314 151228 393320
rect 151082 378040 151138 378049
rect 151082 377975 151138 377984
rect 151188 363730 151216 393314
rect 152476 376718 152504 408478
rect 155224 403028 155276 403034
rect 155224 402970 155276 402976
rect 152464 376712 152516 376718
rect 152464 376654 152516 376660
rect 155236 370530 155264 402970
rect 155224 370524 155276 370530
rect 155224 370466 155276 370472
rect 152556 367804 152608 367810
rect 152556 367746 152608 367752
rect 151176 363724 151228 363730
rect 151176 363666 151228 363672
rect 149794 321736 149850 321745
rect 149794 321671 149850 321680
rect 149702 314800 149758 314809
rect 149702 314735 149758 314744
rect 149716 294642 149744 314735
rect 149704 294636 149756 294642
rect 149704 294578 149756 294584
rect 149058 285696 149114 285705
rect 149058 285631 149114 285640
rect 149072 284306 149100 285631
rect 149808 285054 149836 321671
rect 151082 320240 151138 320249
rect 151082 320175 151138 320184
rect 151096 304366 151124 320175
rect 151174 319424 151230 319433
rect 151174 319359 151230 319368
rect 151188 308446 151216 319359
rect 151268 311908 151320 311914
rect 151268 311850 151320 311856
rect 151176 308440 151228 308446
rect 151176 308382 151228 308388
rect 151084 304360 151136 304366
rect 151084 304302 151136 304308
rect 151174 294536 151230 294545
rect 151174 294471 151230 294480
rect 149796 285048 149848 285054
rect 149796 284990 149848 284996
rect 149704 284980 149756 284986
rect 149704 284922 149756 284928
rect 149060 284300 149112 284306
rect 149060 284242 149112 284248
rect 148968 264920 149020 264926
rect 148968 264862 149020 264868
rect 148508 249144 148560 249150
rect 148508 249086 148560 249092
rect 148416 221536 148468 221542
rect 148416 221478 148468 221484
rect 148416 201544 148468 201550
rect 148416 201486 148468 201492
rect 148428 10334 148456 201486
rect 148506 156088 148562 156097
rect 148506 156023 148562 156032
rect 148520 132394 148548 156023
rect 148508 132388 148560 132394
rect 148508 132330 148560 132336
rect 149716 47598 149744 284922
rect 151082 266384 151138 266393
rect 151082 266319 151138 266328
rect 149794 250472 149850 250481
rect 149794 250407 149850 250416
rect 149808 223553 149836 250407
rect 149794 223544 149850 223553
rect 149794 223479 149850 223488
rect 149704 47592 149756 47598
rect 149704 47534 149756 47540
rect 148416 10328 148468 10334
rect 148416 10270 148468 10276
rect 151096 4894 151124 266319
rect 151188 49026 151216 294471
rect 151280 193866 151308 311850
rect 152464 306468 152516 306474
rect 152464 306410 152516 306416
rect 151360 304360 151412 304366
rect 151360 304302 151412 304308
rect 151372 264314 151400 304302
rect 151360 264308 151412 264314
rect 151360 264250 151412 264256
rect 151268 193860 151320 193866
rect 151268 193802 151320 193808
rect 151176 49020 151228 49026
rect 151176 48962 151228 48968
rect 152476 14482 152504 306410
rect 152568 278050 152596 367746
rect 154488 349852 154540 349858
rect 154488 349794 154540 349800
rect 152648 332648 152700 332654
rect 152648 332590 152700 332596
rect 152660 294710 152688 332590
rect 153934 302560 153990 302569
rect 153934 302495 153990 302504
rect 152648 294704 152700 294710
rect 152648 294646 152700 294652
rect 152740 294636 152792 294642
rect 152740 294578 152792 294584
rect 152752 282169 152780 294578
rect 152738 282160 152794 282169
rect 152738 282095 152794 282104
rect 152556 278044 152608 278050
rect 152556 277986 152608 277992
rect 152648 269884 152700 269890
rect 152648 269826 152700 269832
rect 152554 244896 152610 244905
rect 152554 244831 152610 244840
rect 152568 229809 152596 244831
rect 152554 229800 152610 229809
rect 152554 229735 152610 229744
rect 152554 228304 152610 228313
rect 152554 228239 152610 228248
rect 152568 104174 152596 228239
rect 152660 201550 152688 269826
rect 153844 250504 153896 250510
rect 153844 250446 153896 250452
rect 153856 222154 153884 250446
rect 153844 222148 153896 222154
rect 153844 222090 153896 222096
rect 152648 201544 152700 201550
rect 152648 201486 152700 201492
rect 153844 199436 153896 199442
rect 153844 199378 153896 199384
rect 152648 156052 152700 156058
rect 152648 155994 152700 156000
rect 152660 125594 152688 155994
rect 152648 125588 152700 125594
rect 152648 125530 152700 125536
rect 152556 104168 152608 104174
rect 152556 104110 152608 104116
rect 152556 98048 152608 98054
rect 152556 97990 152608 97996
rect 152568 64802 152596 97990
rect 152556 64796 152608 64802
rect 152556 64738 152608 64744
rect 153856 46306 153884 199378
rect 153948 180130 153976 302495
rect 154500 259418 154528 349794
rect 155316 335368 155368 335374
rect 155316 335310 155368 335316
rect 155222 304056 155278 304065
rect 155222 303991 155278 304000
rect 154488 259412 154540 259418
rect 154488 259354 154540 259360
rect 154500 258777 154528 259354
rect 154486 258768 154542 258777
rect 154486 258703 154542 258712
rect 153936 180124 153988 180130
rect 153936 180066 153988 180072
rect 153936 158840 153988 158846
rect 153936 158782 153988 158788
rect 153948 122806 153976 158782
rect 153936 122800 153988 122806
rect 153936 122742 153988 122748
rect 153844 46300 153896 46306
rect 153844 46242 153896 46248
rect 152464 14476 152516 14482
rect 152464 14418 152516 14424
rect 155236 7614 155264 303991
rect 155328 280906 155356 335310
rect 155788 293962 155816 470562
rect 164148 466540 164200 466546
rect 164148 466482 164200 466488
rect 160100 455524 160152 455530
rect 160100 455466 160152 455472
rect 159456 454096 159508 454102
rect 159456 454038 159508 454044
rect 159364 405748 159416 405754
rect 159364 405690 159416 405696
rect 156604 403028 156656 403034
rect 156604 402970 156656 402976
rect 156616 379438 156644 402970
rect 157984 394800 158036 394806
rect 157984 394742 158036 394748
rect 155960 379432 156012 379438
rect 155960 379374 156012 379380
rect 156604 379432 156656 379438
rect 156604 379374 156656 379380
rect 155868 352572 155920 352578
rect 155868 352514 155920 352520
rect 155776 293956 155828 293962
rect 155776 293898 155828 293904
rect 155316 280900 155368 280906
rect 155316 280842 155368 280848
rect 155316 271176 155368 271182
rect 155316 271118 155368 271124
rect 155328 244905 155356 271118
rect 155408 259548 155460 259554
rect 155408 259490 155460 259496
rect 155314 244896 155370 244905
rect 155314 244831 155370 244840
rect 155316 241936 155368 241942
rect 155316 241878 155368 241884
rect 155328 35222 155356 241878
rect 155420 227730 155448 259490
rect 155408 227724 155460 227730
rect 155408 227666 155460 227672
rect 155406 153232 155462 153241
rect 155406 153167 155462 153176
rect 155420 117230 155448 153167
rect 155880 143449 155908 352514
rect 155972 246362 156000 379374
rect 157996 375329 158024 394742
rect 157982 375320 158038 375329
rect 157982 375255 158038 375264
rect 157996 373994 158024 375255
rect 157996 373966 158208 373994
rect 156604 366376 156656 366382
rect 156604 366318 156656 366324
rect 155960 246356 156012 246362
rect 155960 246298 156012 246304
rect 156616 230450 156644 366318
rect 158074 327720 158130 327729
rect 158074 327655 158130 327664
rect 157984 264988 158036 264994
rect 157984 264930 158036 264936
rect 156696 258732 156748 258738
rect 156696 258674 156748 258680
rect 156708 233209 156736 258674
rect 156788 235272 156840 235278
rect 156788 235214 156840 235220
rect 156694 233200 156750 233209
rect 156694 233135 156750 233144
rect 156604 230444 156656 230450
rect 156604 230386 156656 230392
rect 156708 219434 156736 233135
rect 156800 229090 156828 235214
rect 156788 229084 156840 229090
rect 156788 229026 156840 229032
rect 156800 227866 156828 229026
rect 156788 227860 156840 227866
rect 156788 227802 156840 227808
rect 157248 227860 157300 227866
rect 157248 227802 157300 227808
rect 156616 219406 156736 219434
rect 156616 216617 156644 219406
rect 156602 216608 156658 216617
rect 156602 216543 156658 216552
rect 155866 143440 155922 143449
rect 155866 143375 155922 143384
rect 155408 117224 155460 117230
rect 155408 117166 155460 117172
rect 156616 109002 156644 216543
rect 157260 112470 157288 227802
rect 157248 112464 157300 112470
rect 157248 112406 157300 112412
rect 157260 111858 157288 112406
rect 156696 111852 156748 111858
rect 156696 111794 156748 111800
rect 157248 111852 157300 111858
rect 157248 111794 157300 111800
rect 156604 108996 156656 109002
rect 156604 108938 156656 108944
rect 155408 108384 155460 108390
rect 155408 108326 155460 108332
rect 155420 82754 155448 108326
rect 155408 82748 155460 82754
rect 155408 82690 155460 82696
rect 156708 81297 156736 111794
rect 156694 81288 156750 81297
rect 156694 81223 156750 81232
rect 155316 35216 155368 35222
rect 155316 35158 155368 35164
rect 157996 26926 158024 264930
rect 158088 136649 158116 327655
rect 158180 252822 158208 373966
rect 159376 369753 159404 405690
rect 159362 369744 159418 369753
rect 159362 369679 159418 369688
rect 159376 324358 159404 369679
rect 159364 324352 159416 324358
rect 159364 324294 159416 324300
rect 159376 323678 159404 324294
rect 159364 323672 159416 323678
rect 159364 323614 159416 323620
rect 159362 323096 159418 323105
rect 159362 323031 159418 323040
rect 158168 252816 158220 252822
rect 158168 252758 158220 252764
rect 158180 251938 158208 252758
rect 158168 251932 158220 251938
rect 158168 251874 158220 251880
rect 158074 136640 158130 136649
rect 158074 136575 158130 136584
rect 158088 105602 158116 136575
rect 158076 105596 158128 105602
rect 158076 105538 158128 105544
rect 157984 26920 158036 26926
rect 157984 26862 158036 26868
rect 155224 7608 155276 7614
rect 155224 7550 155276 7556
rect 159376 6186 159404 323031
rect 159468 300150 159496 454038
rect 159548 397520 159600 397526
rect 159548 397462 159600 397468
rect 159560 371249 159588 397462
rect 159546 371240 159602 371249
rect 159546 371175 159602 371184
rect 159560 339522 159588 371175
rect 159548 339516 159600 339522
rect 159548 339458 159600 339464
rect 159456 300144 159508 300150
rect 159456 300086 159508 300092
rect 159456 280084 159508 280090
rect 159456 280026 159508 280032
rect 159468 138038 159496 280026
rect 159560 273970 159588 339458
rect 160112 284374 160140 455466
rect 162124 427100 162176 427106
rect 162124 427042 162176 427048
rect 162136 417450 162164 427042
rect 162124 417444 162176 417450
rect 162124 417386 162176 417392
rect 162768 417444 162820 417450
rect 162768 417386 162820 417392
rect 162124 404388 162176 404394
rect 162124 404330 162176 404336
rect 160744 396772 160796 396778
rect 160744 396714 160796 396720
rect 160756 372609 160784 396714
rect 160742 372600 160798 372609
rect 160742 372535 160798 372544
rect 160756 371385 160784 372535
rect 160190 371376 160246 371385
rect 160190 371311 160246 371320
rect 160742 371376 160798 371385
rect 160742 371311 160798 371320
rect 160100 284368 160152 284374
rect 160100 284310 160152 284316
rect 160112 280090 160140 284310
rect 160100 280084 160152 280090
rect 160100 280026 160152 280032
rect 159548 273964 159600 273970
rect 159548 273906 159600 273912
rect 159548 272536 159600 272542
rect 159548 272478 159600 272484
rect 159560 245614 159588 272478
rect 160204 267734 160232 371311
rect 160742 301608 160798 301617
rect 160742 301543 160798 301552
rect 160112 267706 160232 267734
rect 160112 260794 160140 267706
rect 160020 260766 160140 260794
rect 159548 245608 159600 245614
rect 159548 245550 159600 245556
rect 160020 235929 160048 260766
rect 160756 241942 160784 301543
rect 162136 280158 162164 404330
rect 162780 325009 162808 417386
rect 163596 325712 163648 325718
rect 163596 325654 163648 325660
rect 162766 325000 162822 325009
rect 162766 324935 162822 324944
rect 162400 323672 162452 323678
rect 162400 323614 162452 323620
rect 162306 300112 162362 300121
rect 162306 300047 162362 300056
rect 162124 280152 162176 280158
rect 162124 280094 162176 280100
rect 162214 280120 162270 280129
rect 160928 269816 160980 269822
rect 160928 269758 160980 269764
rect 160836 249076 160888 249082
rect 160836 249018 160888 249024
rect 160744 241936 160796 241942
rect 160744 241878 160796 241884
rect 160742 237416 160798 237425
rect 160742 237351 160798 237360
rect 159546 235920 159602 235929
rect 159546 235855 159602 235864
rect 160006 235920 160062 235929
rect 160006 235855 160062 235864
rect 159560 211818 159588 235855
rect 159548 211812 159600 211818
rect 159548 211754 159600 211760
rect 159456 138032 159508 138038
rect 159456 137974 159508 137980
rect 159468 129742 159496 137974
rect 159456 129736 159508 129742
rect 159456 129678 159508 129684
rect 159560 97986 159588 211754
rect 160756 180849 160784 237351
rect 160848 209574 160876 249018
rect 160940 238649 160968 269758
rect 161020 252816 161072 252822
rect 161020 252758 161072 252764
rect 160926 238640 160982 238649
rect 160926 238575 160982 238584
rect 160940 237425 160968 238575
rect 160926 237416 160982 237425
rect 160926 237351 160982 237360
rect 161032 229770 161060 252758
rect 162136 249762 162164 280094
rect 162214 280055 162270 280064
rect 162124 249756 162176 249762
rect 162124 249698 162176 249704
rect 160928 229764 160980 229770
rect 160928 229706 160980 229712
rect 161020 229764 161072 229770
rect 161020 229706 161072 229712
rect 160940 216646 160968 229706
rect 162228 228313 162256 280055
rect 162320 253230 162348 300047
rect 162412 278905 162440 323614
rect 162676 280832 162728 280838
rect 162676 280774 162728 280780
rect 162398 278896 162454 278905
rect 162398 278831 162454 278840
rect 162308 253224 162360 253230
rect 162308 253166 162360 253172
rect 162214 228304 162270 228313
rect 162214 228239 162270 228248
rect 160928 216640 160980 216646
rect 160928 216582 160980 216588
rect 161388 216640 161440 216646
rect 161388 216582 161440 216588
rect 161296 209772 161348 209778
rect 161296 209714 161348 209720
rect 161308 209574 161336 209714
rect 160836 209568 160888 209574
rect 160836 209510 160888 209516
rect 161296 209568 161348 209574
rect 161296 209510 161348 209516
rect 160742 180840 160798 180849
rect 160742 180775 160798 180784
rect 160756 155281 160784 180775
rect 161308 167657 161336 209510
rect 161294 167648 161350 167657
rect 161294 167583 161350 167592
rect 160742 155272 160798 155281
rect 160742 155207 160798 155216
rect 160834 150648 160890 150657
rect 160834 150583 160890 150592
rect 160744 135312 160796 135318
rect 160744 135254 160796 135260
rect 159548 97980 159600 97986
rect 159548 97922 159600 97928
rect 159364 6180 159416 6186
rect 159364 6122 159416 6128
rect 151084 4888 151136 4894
rect 151084 4830 151136 4836
rect 148322 3360 148378 3369
rect 148322 3295 148378 3304
rect 160756 2106 160784 135254
rect 160848 133278 160876 150583
rect 160926 140040 160982 140049
rect 160926 139975 160982 139984
rect 160836 133272 160888 133278
rect 160836 133214 160888 133220
rect 160940 128489 160968 139975
rect 161400 135969 161428 216582
rect 162124 215960 162176 215966
rect 162124 215902 162176 215908
rect 162136 198286 162164 215902
rect 162584 198688 162636 198694
rect 162584 198630 162636 198636
rect 162596 198286 162624 198630
rect 162124 198280 162176 198286
rect 162124 198222 162176 198228
rect 162584 198280 162636 198286
rect 162584 198222 162636 198228
rect 162596 151842 162624 198222
rect 161480 151836 161532 151842
rect 161480 151778 161532 151784
rect 162584 151836 162636 151842
rect 162584 151778 162636 151784
rect 161492 151065 161520 151778
rect 161478 151056 161534 151065
rect 161478 150991 161534 151000
rect 162688 143682 162716 280774
rect 163504 265056 163556 265062
rect 163504 264998 163556 265004
rect 162768 246356 162820 246362
rect 162768 246298 162820 246304
rect 162780 242962 162808 246298
rect 162768 242956 162820 242962
rect 162768 242898 162820 242904
rect 161480 143676 161532 143682
rect 161480 143618 161532 143624
rect 162676 143676 162728 143682
rect 162676 143618 162728 143624
rect 161386 135960 161442 135969
rect 161492 135930 161520 143618
rect 161386 135895 161442 135904
rect 161480 135924 161532 135930
rect 161480 135866 161532 135872
rect 160926 128480 160982 128489
rect 160926 128415 160982 128424
rect 162124 123480 162176 123486
rect 162124 123422 162176 123428
rect 160836 109744 160888 109750
rect 160836 109686 160888 109692
rect 160848 85542 160876 109686
rect 160836 85536 160888 85542
rect 160836 85478 160888 85484
rect 162136 40730 162164 123422
rect 162216 101516 162268 101522
rect 162216 101458 162268 101464
rect 162228 73098 162256 101458
rect 162780 101454 162808 242898
rect 162768 101448 162820 101454
rect 162768 101390 162820 101396
rect 162216 73092 162268 73098
rect 162216 73034 162268 73040
rect 163516 68338 163544 264998
rect 163608 156670 163636 325654
rect 164160 298110 164188 466482
rect 170496 465180 170548 465186
rect 170496 465122 170548 465128
rect 170404 452668 170456 452674
rect 170404 452610 170456 452616
rect 169024 447908 169076 447914
rect 169024 447850 169076 447856
rect 166356 440292 166408 440298
rect 166356 440234 166408 440240
rect 166264 422952 166316 422958
rect 166264 422894 166316 422900
rect 166276 422346 166304 422894
rect 166264 422340 166316 422346
rect 166264 422282 166316 422288
rect 165526 393408 165582 393417
rect 165526 393343 165582 393352
rect 164884 313336 164936 313342
rect 164884 313278 164936 313284
rect 164896 304366 164924 313278
rect 164884 304360 164936 304366
rect 164884 304302 164936 304308
rect 164240 300144 164292 300150
rect 164240 300086 164292 300092
rect 164252 299538 164280 300086
rect 164240 299532 164292 299538
rect 164240 299474 164292 299480
rect 164148 298104 164200 298110
rect 164148 298046 164200 298052
rect 164160 297430 164188 298046
rect 164148 297424 164200 297430
rect 164148 297366 164200 297372
rect 163688 291848 163740 291854
rect 163688 291790 163740 291796
rect 163700 265577 163728 291790
rect 163686 265568 163742 265577
rect 163686 265503 163742 265512
rect 163688 249756 163740 249762
rect 163688 249698 163740 249704
rect 163700 220794 163728 249698
rect 163688 220788 163740 220794
rect 163688 220730 163740 220736
rect 164148 220788 164200 220794
rect 164148 220730 164200 220736
rect 163596 156664 163648 156670
rect 163596 156606 163648 156612
rect 163608 128314 163636 156606
rect 163596 128308 163648 128314
rect 163596 128250 163648 128256
rect 164160 103494 164188 220730
rect 164252 154562 164280 299474
rect 165540 280158 165568 393343
rect 165620 389292 165672 389298
rect 165620 389234 165672 389240
rect 165528 280152 165580 280158
rect 165528 280094 165580 280100
rect 164884 263628 164936 263634
rect 164884 263570 164936 263576
rect 164240 154556 164292 154562
rect 164240 154498 164292 154504
rect 164148 103488 164200 103494
rect 164148 103430 164200 103436
rect 164160 102814 164188 103430
rect 164148 102808 164200 102814
rect 164148 102750 164200 102756
rect 163504 68332 163556 68338
rect 163504 68274 163556 68280
rect 162124 40724 162176 40730
rect 162124 40666 162176 40672
rect 164896 28286 164924 263570
rect 164976 255332 165028 255338
rect 164976 255274 165028 255280
rect 164988 240786 165016 255274
rect 165632 244934 165660 389234
rect 166276 322250 166304 422282
rect 166368 411942 166396 440234
rect 166356 411936 166408 411942
rect 166356 411878 166408 411884
rect 166908 411936 166960 411942
rect 166908 411878 166960 411884
rect 166920 329390 166948 411878
rect 167734 388784 167790 388793
rect 167734 388719 167790 388728
rect 166356 329384 166408 329390
rect 166356 329326 166408 329332
rect 166908 329384 166960 329390
rect 166908 329326 166960 329332
rect 166368 328506 166396 329326
rect 166356 328500 166408 328506
rect 166356 328442 166408 328448
rect 166264 322244 166316 322250
rect 166264 322186 166316 322192
rect 166262 316296 166318 316305
rect 166262 316231 166318 316240
rect 166276 261526 166304 316231
rect 166368 268394 166396 328442
rect 167644 313404 167696 313410
rect 167644 313346 167696 313352
rect 166908 293276 166960 293282
rect 166908 293218 166960 293224
rect 166816 268660 166868 268666
rect 166816 268602 166868 268608
rect 166356 268388 166408 268394
rect 166356 268330 166408 268336
rect 166264 261520 166316 261526
rect 166264 261462 166316 261468
rect 166264 251252 166316 251258
rect 166264 251194 166316 251200
rect 165620 244928 165672 244934
rect 165620 244870 165672 244876
rect 165632 244322 165660 244870
rect 165620 244316 165672 244322
rect 165620 244258 165672 244264
rect 164976 240780 165028 240786
rect 164976 240722 165028 240728
rect 164976 235272 165028 235278
rect 164976 235214 165028 235220
rect 164988 230450 165016 235214
rect 164976 230444 165028 230450
rect 164976 230386 165028 230392
rect 164988 87650 165016 230386
rect 165068 154556 165120 154562
rect 165068 154498 165120 154504
rect 165080 153338 165108 154498
rect 165068 153332 165120 153338
rect 165068 153274 165120 153280
rect 165080 131102 165108 153274
rect 165068 131096 165120 131102
rect 165068 131038 165120 131044
rect 164976 87644 165028 87650
rect 164976 87586 165028 87592
rect 165528 87644 165580 87650
rect 165528 87586 165580 87592
rect 165540 86970 165568 87586
rect 165528 86964 165580 86970
rect 165528 86906 165580 86912
rect 166276 29646 166304 251194
rect 166448 244316 166500 244322
rect 166448 244258 166500 244264
rect 166356 234184 166408 234190
rect 166356 234126 166408 234132
rect 166368 137873 166396 234126
rect 166460 232558 166488 244258
rect 166828 234598 166856 268602
rect 166816 234592 166868 234598
rect 166816 234534 166868 234540
rect 166828 234190 166856 234534
rect 166816 234184 166868 234190
rect 166816 234126 166868 234132
rect 166448 232552 166500 232558
rect 166448 232494 166500 232500
rect 166354 137864 166410 137873
rect 166354 137799 166410 137808
rect 166368 125594 166396 137799
rect 166356 125588 166408 125594
rect 166356 125530 166408 125536
rect 166356 102876 166408 102882
rect 166356 102818 166408 102824
rect 166368 67522 166396 102818
rect 166448 94580 166500 94586
rect 166448 94522 166500 94528
rect 166460 94489 166488 94522
rect 166920 94489 166948 293218
rect 167656 278118 167684 313346
rect 167644 278112 167696 278118
rect 167644 278054 167696 278060
rect 167644 262268 167696 262274
rect 167644 262210 167696 262216
rect 166446 94480 166502 94489
rect 166446 94415 166502 94424
rect 166906 94480 166962 94489
rect 166906 94415 166962 94424
rect 166356 67516 166408 67522
rect 166356 67458 166408 67464
rect 167656 39370 167684 262210
rect 167748 211138 167776 388719
rect 168378 380216 168434 380225
rect 168378 380151 168380 380160
rect 168432 380151 168434 380160
rect 168380 380122 168432 380128
rect 169036 310486 169064 447850
rect 170416 430574 170444 452610
rect 170404 430568 170456 430574
rect 170404 430510 170456 430516
rect 170404 426420 170456 426426
rect 170404 426362 170456 426368
rect 169206 404424 169262 404433
rect 169206 404359 169262 404368
rect 169114 380216 169170 380225
rect 169114 380151 169170 380160
rect 168380 310480 168432 310486
rect 168380 310422 168432 310428
rect 169024 310480 169076 310486
rect 169024 310422 169076 310428
rect 168392 309806 168420 310422
rect 168380 309800 168432 309806
rect 168380 309742 168432 309748
rect 167828 284368 167880 284374
rect 167828 284310 167880 284316
rect 167840 247722 167868 284310
rect 168392 268666 168420 309742
rect 168380 268660 168432 268666
rect 168380 268602 168432 268608
rect 169024 249824 169076 249830
rect 169024 249766 169076 249772
rect 167828 247716 167880 247722
rect 167828 247658 167880 247664
rect 168288 246356 168340 246362
rect 168288 246298 168340 246304
rect 167736 211132 167788 211138
rect 167736 211074 167788 211080
rect 168300 93226 168328 246298
rect 168378 240136 168434 240145
rect 168378 240071 168434 240080
rect 168392 239329 168420 240071
rect 168378 239320 168434 239329
rect 168378 239255 168434 239264
rect 168288 93220 168340 93226
rect 168288 93162 168340 93168
rect 167644 39364 167696 39370
rect 167644 39306 167696 39312
rect 169036 31074 169064 249766
rect 169128 240145 169156 380151
rect 169220 369753 169248 404359
rect 169206 369744 169262 369753
rect 169206 369679 169262 369688
rect 170416 326398 170444 426362
rect 170508 418130 170536 465122
rect 173806 457056 173862 457065
rect 173806 456991 173862 457000
rect 173820 456822 173848 456991
rect 173624 456816 173676 456822
rect 173624 456758 173676 456764
rect 173808 456816 173860 456822
rect 173808 456758 173860 456764
rect 171876 419552 171928 419558
rect 171876 419494 171928 419500
rect 170496 418124 170548 418130
rect 170496 418066 170548 418072
rect 170494 387832 170550 387841
rect 170494 387767 170550 387776
rect 170508 372065 170536 387767
rect 170494 372056 170550 372065
rect 170494 371991 170550 372000
rect 171046 372056 171102 372065
rect 171046 371991 171102 372000
rect 170956 340196 171008 340202
rect 170956 340138 171008 340144
rect 170404 326392 170456 326398
rect 170404 326334 170456 326340
rect 170494 320376 170550 320385
rect 170494 320311 170550 320320
rect 169206 312216 169262 312225
rect 169206 312151 169262 312160
rect 169220 275330 169248 312151
rect 170404 309188 170456 309194
rect 170404 309130 170456 309136
rect 169666 280936 169722 280945
rect 169666 280871 169722 280880
rect 169208 275324 169260 275330
rect 169208 275266 169260 275272
rect 169576 261588 169628 261594
rect 169576 261530 169628 261536
rect 169114 240136 169170 240145
rect 169114 240071 169170 240080
rect 169588 228993 169616 261530
rect 169574 228984 169630 228993
rect 169574 228919 169630 228928
rect 169588 162081 169616 228919
rect 169574 162072 169630 162081
rect 169574 162007 169630 162016
rect 169116 114572 169168 114578
rect 169116 114514 169168 114520
rect 169128 80034 169156 114514
rect 169680 84114 169708 280871
rect 170416 274650 170444 309130
rect 170508 304298 170536 320311
rect 170496 304292 170548 304298
rect 170496 304234 170548 304240
rect 170496 298784 170548 298790
rect 170496 298726 170548 298732
rect 170404 274644 170456 274650
rect 170404 274586 170456 274592
rect 170404 252612 170456 252618
rect 170404 252554 170456 252560
rect 169760 198620 169812 198626
rect 169760 198562 169812 198568
rect 169772 197946 169800 198562
rect 169760 197940 169812 197946
rect 169760 197882 169812 197888
rect 169668 84108 169720 84114
rect 169668 84050 169720 84056
rect 169116 80028 169168 80034
rect 169116 79970 169168 79976
rect 169024 31068 169076 31074
rect 169024 31010 169076 31016
rect 166264 29640 166316 29646
rect 166264 29582 166316 29588
rect 164884 28280 164936 28286
rect 164884 28222 164936 28228
rect 170416 18630 170444 252554
rect 170508 246265 170536 298726
rect 170588 269136 170640 269142
rect 170588 269078 170640 269084
rect 170494 246256 170550 246265
rect 170494 246191 170550 246200
rect 170496 238128 170548 238134
rect 170496 238070 170548 238076
rect 170508 231810 170536 238070
rect 170600 238066 170628 269078
rect 170968 240009 170996 340138
rect 171060 254590 171088 371991
rect 171782 310720 171838 310729
rect 171782 310655 171838 310664
rect 171796 269890 171824 310655
rect 171784 269884 171836 269890
rect 171784 269826 171836 269832
rect 171782 259584 171838 259593
rect 171782 259519 171838 259528
rect 171048 254584 171100 254590
rect 171048 254526 171100 254532
rect 171140 240848 171192 240854
rect 171140 240790 171192 240796
rect 170954 240000 171010 240009
rect 170954 239935 171010 239944
rect 170588 238060 170640 238066
rect 170588 238002 170640 238008
rect 171152 234025 171180 240790
rect 171138 234016 171194 234025
rect 171138 233951 171194 233960
rect 170496 231804 170548 231810
rect 170496 231746 170548 231752
rect 170508 93906 170536 231746
rect 171046 202192 171102 202201
rect 171046 202127 171102 202136
rect 171060 197946 171088 202127
rect 171048 197940 171100 197946
rect 171048 197882 171100 197888
rect 170586 146568 170642 146577
rect 170586 146503 170642 146512
rect 170600 130422 170628 146503
rect 170588 130416 170640 130422
rect 170588 130358 170640 130364
rect 170496 93900 170548 93906
rect 170496 93842 170548 93848
rect 170508 93158 170536 93842
rect 170496 93152 170548 93158
rect 170496 93094 170548 93100
rect 171796 69698 171824 259519
rect 171888 258738 171916 419494
rect 173164 416084 173216 416090
rect 173164 416026 173216 416032
rect 173070 388376 173126 388385
rect 173070 388311 173126 388320
rect 173084 382265 173112 388311
rect 173176 387569 173204 416026
rect 173162 387560 173218 387569
rect 173162 387495 173218 387504
rect 173070 382256 173126 382265
rect 173070 382191 173126 382200
rect 173084 379438 173112 382191
rect 173072 379432 173124 379438
rect 173072 379374 173124 379380
rect 172428 342916 172480 342922
rect 172428 342858 172480 342864
rect 171968 274712 172020 274718
rect 171968 274654 172020 274660
rect 171876 258732 171928 258738
rect 171876 258674 171928 258680
rect 171980 236706 172008 274654
rect 171968 236700 172020 236706
rect 171968 236642 172020 236648
rect 171876 197940 171928 197946
rect 171876 197882 171928 197888
rect 171888 107642 171916 197882
rect 172440 175273 172468 342858
rect 173636 331294 173664 456758
rect 176658 454336 176714 454345
rect 176658 454271 176714 454280
rect 176672 454073 176700 454271
rect 176658 454064 176714 454073
rect 176658 453999 176714 454008
rect 173808 449200 173860 449206
rect 173808 449142 173860 449148
rect 173716 379432 173768 379438
rect 173716 379374 173768 379380
rect 173624 331288 173676 331294
rect 173624 331230 173676 331236
rect 173254 309496 173310 309505
rect 173254 309431 173310 309440
rect 173164 290556 173216 290562
rect 173164 290498 173216 290504
rect 173176 272610 173204 290498
rect 173164 272604 173216 272610
rect 173164 272546 173216 272552
rect 173268 268462 173296 309431
rect 173636 301510 173664 331230
rect 173624 301504 173676 301510
rect 173624 301446 173676 301452
rect 173256 268456 173308 268462
rect 173256 268398 173308 268404
rect 173164 267776 173216 267782
rect 173164 267718 173216 267724
rect 172426 175264 172482 175273
rect 172426 175199 172482 175208
rect 172440 174593 172468 175199
rect 172426 174584 172482 174593
rect 172426 174519 172482 174528
rect 171876 107636 171928 107642
rect 171876 107578 171928 107584
rect 171784 69692 171836 69698
rect 171784 69634 171836 69640
rect 170404 18624 170456 18630
rect 170404 18566 170456 18572
rect 173176 9042 173204 267718
rect 173346 247616 173402 247625
rect 173346 247551 173402 247560
rect 173360 199442 173388 247551
rect 173728 240825 173756 379374
rect 173820 289814 173848 449142
rect 176568 446412 176620 446418
rect 176568 446354 176620 446360
rect 174544 425740 174596 425746
rect 174544 425682 174596 425688
rect 174556 290465 174584 425682
rect 176476 377460 176528 377466
rect 176476 377402 176528 377408
rect 174636 331356 174688 331362
rect 174636 331298 174688 331304
rect 174542 290456 174598 290465
rect 174542 290391 174598 290400
rect 173808 289808 173860 289814
rect 173808 289750 173860 289756
rect 173808 282940 173860 282946
rect 173808 282882 173860 282888
rect 173714 240816 173770 240825
rect 173714 240751 173770 240760
rect 173348 199436 173400 199442
rect 173348 199378 173400 199384
rect 173254 199336 173310 199345
rect 173254 199271 173310 199280
rect 173268 123486 173296 199271
rect 173348 137284 173400 137290
rect 173348 137226 173400 137232
rect 173256 123480 173308 123486
rect 173256 123422 173308 123428
rect 173360 118658 173388 137226
rect 173820 136610 173848 282882
rect 174556 267170 174584 290391
rect 174544 267164 174596 267170
rect 174544 267106 174596 267112
rect 174544 258120 174596 258126
rect 174544 258062 174596 258068
rect 173808 136604 173860 136610
rect 173808 136546 173860 136552
rect 173808 118720 173860 118726
rect 173808 118662 173860 118668
rect 173348 118652 173400 118658
rect 173348 118594 173400 118600
rect 173256 113212 173308 113218
rect 173256 113154 173308 113160
rect 173268 75857 173296 113154
rect 173820 81326 173848 118662
rect 173808 81320 173860 81326
rect 173808 81262 173860 81268
rect 173254 75848 173310 75857
rect 173254 75783 173310 75792
rect 174556 37942 174584 258062
rect 174648 118726 174676 331298
rect 175924 319524 175976 319530
rect 175924 319466 175976 319472
rect 175936 318850 175964 319466
rect 175924 318844 175976 318850
rect 175924 318786 175976 318792
rect 175936 282946 175964 318786
rect 176108 301504 176160 301510
rect 176108 301446 176160 301452
rect 175924 282940 175976 282946
rect 175924 282882 175976 282888
rect 175278 280800 175334 280809
rect 175278 280735 175334 280744
rect 175292 280158 175320 280735
rect 175280 280152 175332 280158
rect 175280 280094 175332 280100
rect 175188 267028 175240 267034
rect 175188 266970 175240 266976
rect 175200 237289 175228 266970
rect 175292 246362 175320 280094
rect 175924 256760 175976 256766
rect 175924 256702 175976 256708
rect 175280 246356 175332 246362
rect 175280 246298 175332 246304
rect 175186 237280 175242 237289
rect 175186 237215 175242 237224
rect 175200 145625 175228 237215
rect 175186 145616 175242 145625
rect 175186 145551 175242 145560
rect 174636 118720 174688 118726
rect 174636 118662 174688 118668
rect 174544 37936 174596 37942
rect 174544 37878 174596 37884
rect 175936 32434 175964 256702
rect 176016 254584 176068 254590
rect 176016 254526 176068 254532
rect 176028 224942 176056 254526
rect 176016 224936 176068 224942
rect 176016 224878 176068 224884
rect 176028 220153 176056 224878
rect 176014 220144 176070 220153
rect 176014 220079 176070 220088
rect 176028 92177 176056 220079
rect 176120 198014 176148 301446
rect 176488 280906 176516 377402
rect 176580 319530 176608 446354
rect 176660 440292 176712 440298
rect 176660 440234 176712 440240
rect 176672 435402 176700 440234
rect 176660 435396 176712 435402
rect 176660 435338 176712 435344
rect 177316 388385 177344 702782
rect 184848 702568 184900 702574
rect 184848 702510 184900 702516
rect 184204 462460 184256 462466
rect 184204 462402 184256 462408
rect 182824 461032 182876 461038
rect 182824 460974 182876 460980
rect 179234 458416 179290 458425
rect 179234 458351 179290 458360
rect 177946 454336 178002 454345
rect 177946 454271 178002 454280
rect 177302 388376 177358 388385
rect 177302 388311 177358 388320
rect 177960 329934 177988 454271
rect 178684 449948 178736 449954
rect 178684 449890 178736 449896
rect 178696 437442 178724 449890
rect 179248 449857 179276 458351
rect 179328 456816 179380 456822
rect 179328 456758 179380 456764
rect 179234 449848 179290 449857
rect 179234 449783 179290 449792
rect 179248 448633 179276 449783
rect 179234 448624 179290 448633
rect 179234 448559 179290 448568
rect 178684 437436 178736 437442
rect 178684 437378 178736 437384
rect 178684 418192 178736 418198
rect 178684 418134 178736 418140
rect 178040 390584 178092 390590
rect 178040 390526 178092 390532
rect 178052 389065 178080 390526
rect 178038 389056 178094 389065
rect 178038 388991 178094 389000
rect 178696 379409 178724 418134
rect 178774 389056 178830 389065
rect 178774 388991 178830 389000
rect 178682 379400 178738 379409
rect 178682 379335 178738 379344
rect 177488 329928 177540 329934
rect 177488 329870 177540 329876
rect 177948 329928 178000 329934
rect 177948 329870 178000 329876
rect 177304 329860 177356 329866
rect 177304 329802 177356 329808
rect 176568 319524 176620 319530
rect 176568 319466 176620 319472
rect 176660 302932 176712 302938
rect 176660 302874 176712 302880
rect 176672 302326 176700 302874
rect 176660 302320 176712 302326
rect 176660 302262 176712 302268
rect 177316 280945 177344 329802
rect 177396 302932 177448 302938
rect 177396 302874 177448 302880
rect 177302 280936 177358 280945
rect 176476 280900 176528 280906
rect 177302 280871 177358 280880
rect 176476 280842 176528 280848
rect 176660 276684 176712 276690
rect 176660 276626 176712 276632
rect 176672 276010 176700 276626
rect 176660 276004 176712 276010
rect 176660 275946 176712 275952
rect 177304 259548 177356 259554
rect 177304 259490 177356 259496
rect 176108 198008 176160 198014
rect 176108 197950 176160 197956
rect 176014 92168 176070 92177
rect 176014 92103 176070 92112
rect 177316 65550 177344 259490
rect 177408 153785 177436 302874
rect 177500 290494 177528 329870
rect 178684 314696 178736 314702
rect 178684 314638 178736 314644
rect 177488 290488 177540 290494
rect 177488 290430 177540 290436
rect 177580 289876 177632 289882
rect 177580 289818 177632 289824
rect 177592 255270 177620 289818
rect 178696 280838 178724 314638
rect 178684 280832 178736 280838
rect 178684 280774 178736 280780
rect 177856 276004 177908 276010
rect 177856 275946 177908 275952
rect 177580 255264 177632 255270
rect 177580 255206 177632 255212
rect 177868 166326 177896 275946
rect 178684 260908 178736 260914
rect 178684 260850 178736 260856
rect 177948 239692 178000 239698
rect 177948 239634 178000 239640
rect 177960 238678 177988 239634
rect 177948 238672 178000 238678
rect 177948 238614 178000 238620
rect 177960 238134 177988 238614
rect 177948 238128 178000 238134
rect 177948 238070 178000 238076
rect 177948 167680 178000 167686
rect 177948 167622 178000 167628
rect 177856 166320 177908 166326
rect 177856 166262 177908 166268
rect 177394 153776 177450 153785
rect 177394 153711 177450 153720
rect 177394 149152 177450 149161
rect 177394 149087 177450 149096
rect 177408 117298 177436 149087
rect 177396 117292 177448 117298
rect 177396 117234 177448 117240
rect 177394 106312 177450 106321
rect 177394 106247 177450 106256
rect 177408 75721 177436 106247
rect 177960 94518 177988 167622
rect 177948 94512 178000 94518
rect 177948 94454 178000 94460
rect 177394 75712 177450 75721
rect 177394 75647 177450 75656
rect 177304 65544 177356 65550
rect 177304 65486 177356 65492
rect 175924 32428 175976 32434
rect 175924 32370 175976 32376
rect 178696 22778 178724 260850
rect 178788 239698 178816 388991
rect 178958 318880 179014 318889
rect 178958 318815 179014 318824
rect 178868 300960 178920 300966
rect 178868 300902 178920 300908
rect 178880 256018 178908 300902
rect 178972 291854 179000 318815
rect 179340 314702 179368 456758
rect 180154 454472 180210 454481
rect 180154 454407 180210 454416
rect 180062 448624 180118 448633
rect 180062 448559 180118 448568
rect 179328 314696 179380 314702
rect 179328 314638 179380 314644
rect 178960 291848 179012 291854
rect 178960 291790 179012 291796
rect 179328 279472 179380 279478
rect 179328 279414 179380 279420
rect 178868 256012 178920 256018
rect 178868 255954 178920 255960
rect 178958 255368 179014 255377
rect 178958 255303 179014 255312
rect 178776 239692 178828 239698
rect 178776 239634 178828 239640
rect 178972 230489 179000 255303
rect 178958 230480 179014 230489
rect 178958 230415 179014 230424
rect 178972 229094 179000 230415
rect 178972 229066 179276 229094
rect 178774 112160 178830 112169
rect 178774 112095 178830 112104
rect 178788 77081 178816 112095
rect 179248 107681 179276 229066
rect 179234 107672 179290 107681
rect 179234 107607 179290 107616
rect 178868 100088 178920 100094
rect 178868 100030 178920 100036
rect 178774 77072 178830 77081
rect 178774 77007 178830 77016
rect 178880 71738 178908 100030
rect 179340 91050 179368 279414
rect 180076 237969 180104 448559
rect 180168 434722 180196 454407
rect 182086 447944 182142 447953
rect 182086 447879 182142 447888
rect 181444 447840 181496 447846
rect 181444 447782 181496 447788
rect 180156 434716 180208 434722
rect 180156 434658 180208 434664
rect 180708 434036 180760 434042
rect 180708 433978 180760 433984
rect 180156 410576 180208 410582
rect 180156 410518 180208 410524
rect 180168 382265 180196 410518
rect 180246 388240 180302 388249
rect 180246 388175 180302 388184
rect 180154 382256 180210 382265
rect 180154 382191 180210 382200
rect 180154 302424 180210 302433
rect 180154 302359 180210 302368
rect 180168 284986 180196 302359
rect 180156 284980 180208 284986
rect 180156 284922 180208 284928
rect 180156 255332 180208 255338
rect 180156 255274 180208 255280
rect 180062 237960 180118 237969
rect 180062 237895 180118 237904
rect 180062 229800 180118 229809
rect 180062 229735 180118 229744
rect 180076 220153 180104 229735
rect 180062 220144 180118 220153
rect 180062 220079 180118 220088
rect 180062 135960 180118 135969
rect 180062 135895 180118 135904
rect 180076 124166 180104 135895
rect 180064 124160 180116 124166
rect 180064 124102 180116 124108
rect 180064 106956 180116 106962
rect 180064 106898 180116 106904
rect 179328 91044 179380 91050
rect 179328 90986 179380 90992
rect 180076 71738 180104 106898
rect 180168 72457 180196 255274
rect 180260 251870 180288 388175
rect 180720 289134 180748 433978
rect 181456 429146 181484 447782
rect 181444 429140 181496 429146
rect 181444 429082 181496 429088
rect 180800 366444 180852 366450
rect 180800 366386 180852 366392
rect 181352 366444 181404 366450
rect 181352 366386 181404 366392
rect 180708 289128 180760 289134
rect 180708 289070 180760 289076
rect 180812 288561 180840 366386
rect 181364 365809 181392 366386
rect 181350 365800 181406 365809
rect 181350 365735 181406 365744
rect 181996 327752 182048 327758
rect 181996 327694 182048 327700
rect 181444 310616 181496 310622
rect 181444 310558 181496 310564
rect 180798 288552 180854 288561
rect 180798 288487 180854 288496
rect 180340 281580 180392 281586
rect 180340 281522 180392 281528
rect 180248 251864 180300 251870
rect 180248 251806 180300 251812
rect 180352 240009 180380 281522
rect 181456 276010 181484 310558
rect 181536 281580 181588 281586
rect 181536 281522 181588 281528
rect 181444 276004 181496 276010
rect 181444 275946 181496 275952
rect 181444 271924 181496 271930
rect 181444 271866 181496 271872
rect 180800 267164 180852 267170
rect 180800 267106 180852 267112
rect 180812 246378 180840 267106
rect 180720 246350 180840 246378
rect 180338 240000 180394 240009
rect 180338 239935 180394 239944
rect 180720 233209 180748 246350
rect 180706 233200 180762 233209
rect 180706 233135 180762 233144
rect 180720 115938 180748 233135
rect 181456 167793 181484 271866
rect 181548 264926 181576 281522
rect 181536 264920 181588 264926
rect 181536 264862 181588 264868
rect 181626 244896 181682 244905
rect 181626 244831 181682 244840
rect 181536 240372 181588 240378
rect 181536 240314 181588 240320
rect 181548 234569 181576 240314
rect 181640 235385 181668 244831
rect 182008 241534 182036 327694
rect 182100 320113 182128 447879
rect 182180 351892 182232 351898
rect 182180 351834 182232 351840
rect 182086 320104 182142 320113
rect 182086 320039 182142 320048
rect 182100 319462 182128 320039
rect 182088 319456 182140 319462
rect 182088 319398 182140 319404
rect 181996 241528 182048 241534
rect 181996 241470 182048 241476
rect 182192 240106 182220 351834
rect 182836 261526 182864 460974
rect 183466 452976 183522 452985
rect 183466 452911 183522 452920
rect 182916 365016 182968 365022
rect 182916 364958 182968 364964
rect 182928 351898 182956 364958
rect 182916 351892 182968 351898
rect 182916 351834 182968 351840
rect 183480 342922 183508 452911
rect 184216 439521 184244 462402
rect 184202 439512 184258 439521
rect 184202 439447 184258 439456
rect 183468 342916 183520 342922
rect 183468 342858 183520 342864
rect 184216 338745 184244 439447
rect 184296 398880 184348 398886
rect 184296 398822 184348 398828
rect 184308 365702 184336 398822
rect 184860 396778 184888 702510
rect 188988 484424 189040 484430
rect 188988 484366 189040 484372
rect 186964 462392 187016 462398
rect 186964 462334 187016 462340
rect 187056 462392 187108 462398
rect 187056 462334 187108 462340
rect 185584 460964 185636 460970
rect 185584 460906 185636 460912
rect 185596 433226 185624 460906
rect 186320 445732 186372 445738
rect 186320 445674 186372 445680
rect 186332 445058 186360 445674
rect 186320 445052 186372 445058
rect 186320 444994 186372 445000
rect 185768 439544 185820 439550
rect 185768 439486 185820 439492
rect 185780 439006 185808 439486
rect 185768 439000 185820 439006
rect 185768 438942 185820 438948
rect 186136 439000 186188 439006
rect 186136 438942 186188 438948
rect 185584 433220 185636 433226
rect 185584 433162 185636 433168
rect 184848 396772 184900 396778
rect 184848 396714 184900 396720
rect 184388 392080 184440 392086
rect 184388 392022 184440 392028
rect 184296 365696 184348 365702
rect 184296 365638 184348 365644
rect 184202 338736 184258 338745
rect 184202 338671 184258 338680
rect 184308 334626 184336 365638
rect 184400 359514 184428 392022
rect 186044 387184 186096 387190
rect 186044 387126 186096 387132
rect 186056 382226 186084 387126
rect 186044 382220 186096 382226
rect 186044 382162 186096 382168
rect 186056 380934 186084 382162
rect 186044 380928 186096 380934
rect 186044 380870 186096 380876
rect 184388 359508 184440 359514
rect 184388 359450 184440 359456
rect 184296 334620 184348 334626
rect 184296 334562 184348 334568
rect 183468 333260 183520 333266
rect 183468 333202 183520 333208
rect 182916 273284 182968 273290
rect 182916 273226 182968 273232
rect 182824 261520 182876 261526
rect 182824 261462 182876 261468
rect 182824 253972 182876 253978
rect 182824 253914 182876 253920
rect 182270 240816 182326 240825
rect 182270 240751 182326 240760
rect 182180 240100 182232 240106
rect 182180 240042 182232 240048
rect 181626 235376 181682 235385
rect 181626 235311 181682 235320
rect 181534 234560 181590 234569
rect 181534 234495 181590 234504
rect 181548 212498 181576 234495
rect 182284 214713 182312 240751
rect 182270 214704 182326 214713
rect 182270 214639 182326 214648
rect 181536 212492 181588 212498
rect 181536 212434 181588 212440
rect 182088 212492 182140 212498
rect 182088 212434 182140 212440
rect 181536 181552 181588 181558
rect 181536 181494 181588 181500
rect 181442 167784 181498 167793
rect 181442 167719 181498 167728
rect 181444 149116 181496 149122
rect 181444 149058 181496 149064
rect 181456 120086 181484 149058
rect 181548 146946 181576 181494
rect 181536 146940 181588 146946
rect 181536 146882 181588 146888
rect 181548 122126 181576 146882
rect 181536 122120 181588 122126
rect 181536 122062 181588 122068
rect 181996 122120 182048 122126
rect 181996 122062 182048 122068
rect 181444 120080 181496 120086
rect 181444 120022 181496 120028
rect 182008 118658 182036 122062
rect 181996 118652 182048 118658
rect 181996 118594 182048 118600
rect 181996 117972 182048 117978
rect 181996 117914 182048 117920
rect 180708 115932 180760 115938
rect 180708 115874 180760 115880
rect 181258 79928 181314 79937
rect 181258 79863 181314 79872
rect 181272 78606 181300 79863
rect 181260 78600 181312 78606
rect 181260 78542 181312 78548
rect 180154 72448 180210 72457
rect 180154 72383 180210 72392
rect 178868 71732 178920 71738
rect 178868 71674 178920 71680
rect 180064 71732 180116 71738
rect 180064 71674 180116 71680
rect 182008 47598 182036 117914
rect 182100 79937 182128 212434
rect 182836 148374 182864 253914
rect 182928 220114 182956 273226
rect 183480 245682 183508 333202
rect 184400 328681 184428 359450
rect 184756 341556 184808 341562
rect 184756 341498 184808 341504
rect 184386 328672 184442 328681
rect 184386 328607 184442 328616
rect 184204 326392 184256 326398
rect 184204 326334 184256 326340
rect 184216 317422 184244 326334
rect 184400 325694 184428 328607
rect 184400 325666 184612 325694
rect 184204 317416 184256 317422
rect 184204 317358 184256 317364
rect 184584 309126 184612 325666
rect 184664 317416 184716 317422
rect 184664 317358 184716 317364
rect 184676 316062 184704 317358
rect 184664 316056 184716 316062
rect 184664 315998 184716 316004
rect 184572 309120 184624 309126
rect 184572 309062 184624 309068
rect 184202 305280 184258 305289
rect 184202 305215 184258 305224
rect 184216 290562 184244 305215
rect 184204 290556 184256 290562
rect 184204 290498 184256 290504
rect 184204 289128 184256 289134
rect 184204 289070 184256 289076
rect 184216 256222 184244 289070
rect 184676 283286 184704 315998
rect 184664 283280 184716 283286
rect 184664 283222 184716 283228
rect 184296 257372 184348 257378
rect 184296 257314 184348 257320
rect 184204 256216 184256 256222
rect 184204 256158 184256 256164
rect 184202 254552 184258 254561
rect 184202 254487 184258 254496
rect 183468 245676 183520 245682
rect 183468 245618 183520 245624
rect 184216 240825 184244 254487
rect 184202 240816 184258 240825
rect 184202 240751 184258 240760
rect 184308 233918 184336 257314
rect 184768 237386 184796 341498
rect 184848 337476 184900 337482
rect 184848 337418 184900 337424
rect 184860 287774 184888 337418
rect 186148 311982 186176 438942
rect 186976 436082 187004 462334
rect 187068 448497 187096 462334
rect 187606 455560 187662 455569
rect 187606 455495 187662 455504
rect 187514 452840 187570 452849
rect 187514 452775 187570 452784
rect 187146 450256 187202 450265
rect 187146 450191 187202 450200
rect 187054 448488 187110 448497
rect 187054 448423 187110 448432
rect 187160 436801 187188 450191
rect 187146 436792 187202 436801
rect 187146 436727 187202 436736
rect 186964 436076 187016 436082
rect 186964 436018 187016 436024
rect 187056 418804 187108 418810
rect 187056 418746 187108 418752
rect 186228 408536 186280 408542
rect 186228 408478 186280 408484
rect 185584 311976 185636 311982
rect 185584 311918 185636 311924
rect 186136 311976 186188 311982
rect 186136 311918 186188 311924
rect 184848 287768 184900 287774
rect 184848 287710 184900 287716
rect 185596 286346 185624 311918
rect 186044 303748 186096 303754
rect 186044 303690 186096 303696
rect 185584 286340 185636 286346
rect 185584 286282 185636 286288
rect 184848 274780 184900 274786
rect 184848 274722 184900 274728
rect 184756 237380 184808 237386
rect 184756 237322 184808 237328
rect 184296 233912 184348 233918
rect 184296 233854 184348 233860
rect 182916 220108 182968 220114
rect 182916 220050 182968 220056
rect 184756 191140 184808 191146
rect 184756 191082 184808 191088
rect 183468 182844 183520 182850
rect 183468 182786 183520 182792
rect 183008 161560 183060 161566
rect 183008 161502 183060 161508
rect 182824 148368 182876 148374
rect 182824 148310 182876 148316
rect 182916 143608 182968 143614
rect 182916 143550 182968 143556
rect 182824 136672 182876 136678
rect 182824 136614 182876 136620
rect 182836 131102 182864 136614
rect 182824 131096 182876 131102
rect 182824 131038 182876 131044
rect 182086 79928 182142 79937
rect 182086 79863 182142 79872
rect 182836 50386 182864 131038
rect 182928 117298 182956 143550
rect 183020 137290 183048 161502
rect 183480 160857 183508 182786
rect 183466 160848 183522 160857
rect 183466 160783 183522 160792
rect 183480 160138 183508 160783
rect 183468 160132 183520 160138
rect 183468 160074 183520 160080
rect 184204 160132 184256 160138
rect 184204 160074 184256 160080
rect 183098 143712 183154 143721
rect 183098 143647 183154 143656
rect 183008 137284 183060 137290
rect 183008 137226 183060 137232
rect 183112 127634 183140 143647
rect 184216 131209 184244 160074
rect 184664 148368 184716 148374
rect 184664 148310 184716 148316
rect 184296 146260 184348 146266
rect 184296 146202 184348 146208
rect 184308 144974 184336 146202
rect 184296 144968 184348 144974
rect 184296 144910 184348 144916
rect 184308 141438 184336 144910
rect 184296 141432 184348 141438
rect 184296 141374 184348 141380
rect 184202 131200 184258 131209
rect 184202 131135 184258 131144
rect 183100 127628 183152 127634
rect 183100 127570 183152 127576
rect 184204 118652 184256 118658
rect 184204 118594 184256 118600
rect 182916 117292 182968 117298
rect 182916 117234 182968 117240
rect 183008 103556 183060 103562
rect 183008 103498 183060 103504
rect 182916 102264 182968 102270
rect 182916 102206 182968 102212
rect 182928 75818 182956 102206
rect 183020 81394 183048 103498
rect 183560 93220 183612 93226
rect 183560 93162 183612 93168
rect 183008 81388 183060 81394
rect 183008 81330 183060 81336
rect 182916 75812 182968 75818
rect 182916 75754 182968 75760
rect 183572 60722 183600 93162
rect 183560 60716 183612 60722
rect 183560 60658 183612 60664
rect 182824 50380 182876 50386
rect 182824 50322 182876 50328
rect 181996 47592 182048 47598
rect 181996 47534 182048 47540
rect 184216 37942 184244 118594
rect 184296 100020 184348 100026
rect 184296 99962 184348 99968
rect 184308 92478 184336 99962
rect 184296 92472 184348 92478
rect 184296 92414 184348 92420
rect 184676 86970 184704 148310
rect 184768 108225 184796 191082
rect 184860 146266 184888 274722
rect 185676 259480 185728 259486
rect 185676 259422 185728 259428
rect 185584 254040 185636 254046
rect 185584 253982 185636 253988
rect 184848 146260 184900 146266
rect 184848 146202 184900 146208
rect 185490 129840 185546 129849
rect 185490 129775 185546 129784
rect 185504 129742 185532 129775
rect 185492 129736 185544 129742
rect 185492 129678 185544 129684
rect 184754 108216 184810 108225
rect 184754 108151 184810 108160
rect 184664 86964 184716 86970
rect 184664 86906 184716 86912
rect 185596 73846 185624 253982
rect 185688 230450 185716 259422
rect 186056 254017 186084 303690
rect 186134 292360 186190 292369
rect 186134 292295 186190 292304
rect 186148 291281 186176 292295
rect 186134 291272 186190 291281
rect 186134 291207 186190 291216
rect 186042 254008 186098 254017
rect 186042 253943 186098 253952
rect 185676 230444 185728 230450
rect 185676 230386 185728 230392
rect 186148 222873 186176 291207
rect 186240 246362 186268 408478
rect 187068 387705 187096 418746
rect 187148 409148 187200 409154
rect 187148 409090 187200 409096
rect 187054 387696 187110 387705
rect 187054 387631 187110 387640
rect 186964 387116 187016 387122
rect 186964 387058 187016 387064
rect 186320 380928 186372 380934
rect 186320 380870 186372 380876
rect 186228 246356 186280 246362
rect 186228 246298 186280 246304
rect 186332 240378 186360 380870
rect 186976 351898 187004 387058
rect 187160 383489 187188 409090
rect 187146 383480 187202 383489
rect 187146 383415 187202 383424
rect 187528 381614 187556 452775
rect 187620 451926 187648 455495
rect 187608 451920 187660 451926
rect 187608 451862 187660 451868
rect 188344 451920 188396 451926
rect 188344 451862 188396 451868
rect 187608 445732 187660 445738
rect 187608 445674 187660 445680
rect 187516 381608 187568 381614
rect 187516 381550 187568 381556
rect 186964 351892 187016 351898
rect 186964 351834 187016 351840
rect 187516 351892 187568 351898
rect 187516 351834 187568 351840
rect 186962 321600 187018 321609
rect 186962 321535 187018 321544
rect 186976 287706 187004 321535
rect 187056 309256 187108 309262
rect 187056 309198 187108 309204
rect 186964 287700 187016 287706
rect 186964 287642 187016 287648
rect 187068 282985 187096 309198
rect 187528 298790 187556 351834
rect 187620 321609 187648 445674
rect 187698 415984 187754 415993
rect 187698 415919 187700 415928
rect 187752 415919 187754 415928
rect 187700 415890 187752 415896
rect 188356 326398 188384 451862
rect 188436 447160 188488 447166
rect 188436 447102 188488 447108
rect 188448 433294 188476 447102
rect 188436 433288 188488 433294
rect 188436 433230 188488 433236
rect 188436 420980 188488 420986
rect 188436 420922 188488 420928
rect 188448 385801 188476 420922
rect 189000 415954 189028 484366
rect 189722 459640 189778 459649
rect 189722 459575 189778 459584
rect 188988 415948 189040 415954
rect 188988 415890 189040 415896
rect 188896 409896 188948 409902
rect 188896 409838 188948 409844
rect 188528 393372 188580 393378
rect 188528 393314 188580 393320
rect 188540 387297 188568 393314
rect 188526 387288 188582 387297
rect 188526 387223 188582 387232
rect 188434 385792 188490 385801
rect 188434 385727 188490 385736
rect 188540 375329 188568 387223
rect 188526 375320 188582 375329
rect 188526 375255 188582 375264
rect 188908 327729 188936 409838
rect 188988 380316 189040 380322
rect 188988 380258 189040 380264
rect 188894 327720 188950 327729
rect 188894 327655 188950 327664
rect 188344 326392 188396 326398
rect 188344 326334 188396 326340
rect 187606 321600 187662 321609
rect 187606 321535 187662 321544
rect 188342 317520 188398 317529
rect 188342 317455 188398 317464
rect 187700 309120 187752 309126
rect 187700 309062 187752 309068
rect 187516 298784 187568 298790
rect 187516 298726 187568 298732
rect 187712 293282 187740 309062
rect 187700 293276 187752 293282
rect 187700 293218 187752 293224
rect 188356 286385 188384 317455
rect 188528 301028 188580 301034
rect 188528 300970 188580 300976
rect 188342 286376 188398 286385
rect 188342 286311 188398 286320
rect 187700 283280 187752 283286
rect 187700 283222 187752 283228
rect 186410 282976 186466 282985
rect 186410 282911 186466 282920
rect 187054 282976 187110 282985
rect 187054 282911 187110 282920
rect 186424 274786 186452 282911
rect 186412 274780 186464 274786
rect 186412 274722 186464 274728
rect 187056 274780 187108 274786
rect 187056 274722 187108 274728
rect 186962 241632 187018 241641
rect 186962 241567 187018 241576
rect 186320 240372 186372 240378
rect 186320 240314 186372 240320
rect 186134 222864 186190 222873
rect 186134 222799 186190 222808
rect 186228 187672 186280 187678
rect 186228 187614 186280 187620
rect 185768 151836 185820 151842
rect 185768 151778 185820 151784
rect 185676 129736 185728 129742
rect 185676 129678 185728 129684
rect 185584 73840 185636 73846
rect 185584 73782 185636 73788
rect 184296 60716 184348 60722
rect 184296 60658 184348 60664
rect 184308 54534 184336 60658
rect 184296 54528 184348 54534
rect 184296 54470 184348 54476
rect 184204 37936 184256 37942
rect 184204 37878 184256 37884
rect 178684 22772 178736 22778
rect 178684 22714 178736 22720
rect 185688 19990 185716 129678
rect 185780 121446 185808 151778
rect 185768 121440 185820 121446
rect 185768 121382 185820 121388
rect 186240 100706 186268 187614
rect 186320 166388 186372 166394
rect 186320 166330 186372 166336
rect 186332 165646 186360 166330
rect 186320 165640 186372 165646
rect 186320 165582 186372 165588
rect 186976 156641 187004 241567
rect 187068 224262 187096 274722
rect 187148 269204 187200 269210
rect 187148 269146 187200 269152
rect 187160 238105 187188 269146
rect 187146 238096 187202 238105
rect 187146 238031 187202 238040
rect 187712 227798 187740 283222
rect 188540 271250 188568 300970
rect 188528 271244 188580 271250
rect 188528 271186 188580 271192
rect 188436 270632 188488 270638
rect 188436 270574 188488 270580
rect 188344 248464 188396 248470
rect 188344 248406 188396 248412
rect 188356 233889 188384 248406
rect 188342 233880 188398 233889
rect 188342 233815 188398 233824
rect 187700 227792 187752 227798
rect 187700 227734 187752 227740
rect 188344 227792 188396 227798
rect 188344 227734 188396 227740
rect 187056 224256 187108 224262
rect 187056 224198 187108 224204
rect 187608 166388 187660 166394
rect 187608 166330 187660 166336
rect 187054 162072 187110 162081
rect 187054 162007 187110 162016
rect 186962 156632 187018 156641
rect 186962 156567 187018 156576
rect 186964 154624 187016 154630
rect 186964 154566 187016 154572
rect 186976 133929 187004 154566
rect 187068 144129 187096 162007
rect 187054 144120 187110 144129
rect 187054 144055 187110 144064
rect 187148 143608 187200 143614
rect 187148 143550 187200 143556
rect 186962 133920 187018 133929
rect 186962 133855 187018 133864
rect 187160 133210 187188 143550
rect 187148 133204 187200 133210
rect 187148 133146 187200 133152
rect 187620 131510 187648 166330
rect 187608 131504 187660 131510
rect 187608 131446 187660 131452
rect 186320 129804 186372 129810
rect 186320 129746 186372 129752
rect 186332 125594 186360 129746
rect 187608 128444 187660 128450
rect 187608 128386 187660 128392
rect 186320 125588 186372 125594
rect 186320 125530 186372 125536
rect 186964 110492 187016 110498
rect 186964 110434 187016 110440
rect 186318 108216 186374 108225
rect 186318 108151 186374 108160
rect 186332 107817 186360 108151
rect 186318 107808 186374 107817
rect 186318 107743 186374 107752
rect 186228 100700 186280 100706
rect 186228 100642 186280 100648
rect 186332 84153 186360 107743
rect 186976 93838 187004 110434
rect 187516 98048 187568 98054
rect 187516 97990 187568 97996
rect 186964 93832 187016 93838
rect 186964 93774 187016 93780
rect 187528 92041 187556 97990
rect 187514 92032 187570 92041
rect 187514 91967 187570 91976
rect 186318 84144 186374 84153
rect 186318 84079 186374 84088
rect 186332 82929 186360 84079
rect 186318 82920 186374 82929
rect 186318 82855 186374 82864
rect 186962 82920 187018 82929
rect 186962 82855 187018 82864
rect 186976 51746 187004 82855
rect 187620 65550 187648 128386
rect 187700 120760 187752 120766
rect 187700 120702 187752 120708
rect 187712 120222 187740 120702
rect 187700 120216 187752 120222
rect 187700 120158 187752 120164
rect 188356 117230 188384 227734
rect 188448 222902 188476 270574
rect 189000 238746 189028 380258
rect 189078 327312 189134 327321
rect 189078 327247 189134 327256
rect 189092 327146 189120 327247
rect 189080 327140 189132 327146
rect 189080 327082 189132 327088
rect 189736 295934 189764 459575
rect 191196 454164 191248 454170
rect 191196 454106 191248 454112
rect 191102 451480 191158 451489
rect 191102 451415 191158 451424
rect 189816 451376 189868 451382
rect 189816 451318 189868 451324
rect 189828 436762 189856 451318
rect 191010 447808 191066 447817
rect 191010 447743 191066 447752
rect 191024 447166 191052 447743
rect 191012 447160 191064 447166
rect 191012 447102 191064 447108
rect 189816 436756 189868 436762
rect 189816 436698 189868 436704
rect 191116 434042 191144 451415
rect 191208 445738 191236 454106
rect 191654 449168 191710 449177
rect 191654 449103 191710 449112
rect 191668 447914 191696 449103
rect 191656 447908 191708 447914
rect 191656 447850 191708 447856
rect 191654 446448 191710 446457
rect 191654 446383 191710 446392
rect 191668 445806 191696 446383
rect 191656 445800 191708 445806
rect 191656 445742 191708 445748
rect 191196 445732 191248 445738
rect 191196 445674 191248 445680
rect 191654 442096 191710 442105
rect 191654 442031 191710 442040
rect 191668 441697 191696 442031
rect 191654 441688 191710 441697
rect 191654 441623 191710 441632
rect 191378 440736 191434 440745
rect 191378 440671 191434 440680
rect 191392 440298 191420 440671
rect 191380 440292 191432 440298
rect 191380 440234 191432 440240
rect 191378 439376 191434 439385
rect 191378 439311 191434 439320
rect 191392 438938 191420 439311
rect 191380 438932 191432 438938
rect 191380 438874 191432 438880
rect 191564 438184 191616 438190
rect 191564 438126 191616 438132
rect 191576 438025 191604 438126
rect 191562 438016 191618 438025
rect 191562 437951 191618 437960
rect 191564 436076 191616 436082
rect 191564 436018 191616 436024
rect 191576 435305 191604 436018
rect 191562 435296 191618 435305
rect 191562 435231 191618 435240
rect 191104 434036 191156 434042
rect 191104 433978 191156 433984
rect 190644 433220 190696 433226
rect 190644 433162 190696 433168
rect 190656 432313 190684 433162
rect 190642 432304 190698 432313
rect 190642 432239 190698 432248
rect 191196 431248 191248 431254
rect 191196 431190 191248 431196
rect 191102 430944 191158 430953
rect 191102 430879 191158 430888
rect 191116 430574 191144 430879
rect 191104 430568 191156 430574
rect 191104 430510 191156 430516
rect 190642 426864 190698 426873
rect 190642 426799 190698 426808
rect 190656 426494 190684 426799
rect 190644 426488 190696 426494
rect 190644 426430 190696 426436
rect 190642 422512 190698 422521
rect 190642 422447 190698 422456
rect 190656 422346 190684 422447
rect 190644 422340 190696 422346
rect 190644 422282 190696 422288
rect 190366 421016 190422 421025
rect 190366 420951 190422 420960
rect 189816 394732 189868 394738
rect 189816 394674 189868 394680
rect 189828 383654 189856 394674
rect 189816 383648 189868 383654
rect 189816 383590 189868 383596
rect 190380 336054 190408 420951
rect 190644 415948 190696 415954
rect 190644 415890 190696 415896
rect 190656 415449 190684 415890
rect 190642 415440 190698 415449
rect 190642 415375 190698 415384
rect 191010 410000 191066 410009
rect 191010 409935 191066 409944
rect 191024 409902 191052 409935
rect 191012 409896 191064 409902
rect 191012 409838 191064 409844
rect 191010 408640 191066 408649
rect 191010 408575 191066 408584
rect 191024 408542 191052 408575
rect 191012 408536 191064 408542
rect 191012 408478 191064 408484
rect 190826 398576 190882 398585
rect 190826 398511 190882 398520
rect 190840 397526 190868 398511
rect 190828 397520 190880 397526
rect 190828 397462 190880 397468
rect 190826 395856 190882 395865
rect 190826 395791 190882 395800
rect 190840 394806 190868 395791
rect 190828 394800 190880 394806
rect 190828 394742 190880 394748
rect 190826 394496 190882 394505
rect 190826 394431 190882 394440
rect 190458 393408 190514 393417
rect 190840 393378 190868 394431
rect 190458 393343 190514 393352
rect 190828 393372 190880 393378
rect 190472 391785 190500 393343
rect 190828 393314 190880 393320
rect 190458 391776 190514 391785
rect 190458 391711 190514 391720
rect 190368 336048 190420 336054
rect 190368 335990 190420 335996
rect 190366 327312 190422 327321
rect 190366 327247 190422 327256
rect 189906 302288 189962 302297
rect 189906 302223 189962 302232
rect 189080 295928 189132 295934
rect 189080 295870 189132 295876
rect 189724 295928 189776 295934
rect 189724 295870 189776 295876
rect 189092 267034 189120 295870
rect 189814 295352 189870 295361
rect 189814 295287 189870 295296
rect 189828 280809 189856 295287
rect 189920 294642 189948 302223
rect 189908 294636 189960 294642
rect 189908 294578 189960 294584
rect 189814 280800 189870 280809
rect 189814 280735 189870 280744
rect 190276 278044 190328 278050
rect 190276 277986 190328 277992
rect 189080 267028 189132 267034
rect 189080 266970 189132 266976
rect 189816 251864 189868 251870
rect 189816 251806 189868 251812
rect 189722 247072 189778 247081
rect 189722 247007 189778 247016
rect 188988 238740 189040 238746
rect 188988 238682 189040 238688
rect 188436 222896 188488 222902
rect 188436 222838 188488 222844
rect 189736 217297 189764 247007
rect 189828 233073 189856 251806
rect 189906 245712 189962 245721
rect 189906 245647 189962 245656
rect 189920 235249 189948 245647
rect 190288 245614 190316 277986
rect 190380 251870 190408 327247
rect 190460 316736 190512 316742
rect 190460 316678 190512 316684
rect 190472 315246 190500 316678
rect 190460 315240 190512 315246
rect 190460 315182 190512 315188
rect 191012 298852 191064 298858
rect 191012 298794 191064 298800
rect 191024 298761 191052 298794
rect 191010 298752 191066 298761
rect 191010 298687 191066 298696
rect 191116 286793 191144 430510
rect 191208 429593 191236 431190
rect 191194 429584 191250 429593
rect 191194 429519 191250 429528
rect 191668 429434 191696 441623
rect 191484 429406 191696 429434
rect 191484 422294 191512 429406
rect 191760 429298 191788 703394
rect 202800 702642 202828 703520
rect 214564 703316 214616 703322
rect 214564 703258 214616 703264
rect 213184 702908 213236 702914
rect 213184 702850 213236 702856
rect 202788 702636 202840 702642
rect 202788 702578 202840 702584
rect 202144 477556 202196 477562
rect 202144 477498 202196 477504
rect 194598 466576 194654 466585
rect 194598 466511 194654 466520
rect 194612 460934 194640 466511
rect 202156 461378 202184 477498
rect 202880 472116 202932 472122
rect 202880 472058 202932 472064
rect 201500 461372 201552 461378
rect 201500 461314 201552 461320
rect 202144 461372 202196 461378
rect 202144 461314 202196 461320
rect 201512 460934 201540 461314
rect 202156 460970 202184 461314
rect 202144 460964 202196 460970
rect 194612 460906 195192 460934
rect 201512 460906 201816 460934
rect 202144 460906 202196 460912
rect 202892 460934 202920 472058
rect 213196 463690 213224 702850
rect 212632 463684 212684 463690
rect 212632 463626 212684 463632
rect 213184 463684 213236 463690
rect 213184 463626 213236 463632
rect 212644 462466 212672 463626
rect 212632 462460 212684 462466
rect 212632 462402 212684 462408
rect 202892 460906 203656 460934
rect 193404 456884 193456 456890
rect 193404 456826 193456 456832
rect 192666 455696 192722 455705
rect 192666 455631 192722 455640
rect 192484 452668 192536 452674
rect 192484 452610 192536 452616
rect 191840 451308 191892 451314
rect 191840 451250 191892 451256
rect 191852 446418 191880 451250
rect 191840 446412 191892 446418
rect 191840 446354 191892 446360
rect 192496 442950 192524 452610
rect 192576 450560 192628 450566
rect 192576 450502 192628 450508
rect 192484 442944 192536 442950
rect 192484 442886 192536 442892
rect 192482 436656 192538 436665
rect 192482 436591 192538 436600
rect 191668 429270 191788 429298
rect 191668 428074 191696 429270
rect 191748 429140 191800 429146
rect 191748 429082 191800 429088
rect 191760 428233 191788 429082
rect 191746 428224 191802 428233
rect 191746 428159 191802 428168
rect 191668 428046 191788 428074
rect 191760 425746 191788 428046
rect 191748 425740 191800 425746
rect 191748 425682 191800 425688
rect 191760 425513 191788 425682
rect 191746 425504 191802 425513
rect 191746 425439 191802 425448
rect 191484 422266 191696 422294
rect 191668 402974 191696 422266
rect 191746 419792 191802 419801
rect 191746 419727 191802 419736
rect 191760 419558 191788 419727
rect 191748 419552 191800 419558
rect 191748 419494 191800 419500
rect 191746 418432 191802 418441
rect 191746 418367 191802 418376
rect 191760 418198 191788 418367
rect 191748 418192 191800 418198
rect 191748 418134 191800 418140
rect 191748 417444 191800 417450
rect 191748 417386 191800 417392
rect 191760 417081 191788 417386
rect 191746 417072 191802 417081
rect 191746 417007 191802 417016
rect 191746 414080 191802 414089
rect 191746 414015 191748 414024
rect 191800 414015 191802 414024
rect 191748 413986 191800 413992
rect 191748 411936 191800 411942
rect 191748 411878 191800 411884
rect 191760 411369 191788 411878
rect 191746 411360 191802 411369
rect 191746 411295 191802 411304
rect 191746 407008 191802 407017
rect 191746 406943 191802 406952
rect 191760 405754 191788 406943
rect 191748 405748 191800 405754
rect 191748 405690 191800 405696
rect 191746 405648 191802 405657
rect 191746 405583 191802 405592
rect 191760 404394 191788 405583
rect 191748 404388 191800 404394
rect 191748 404330 191800 404336
rect 191746 404288 191802 404297
rect 191746 404223 191802 404232
rect 191760 403034 191788 404223
rect 191484 402946 191696 402974
rect 191748 403028 191800 403034
rect 191748 402970 191800 402976
rect 191484 396522 191512 402946
rect 191654 402384 191710 402393
rect 191654 402319 191710 402328
rect 191668 396658 191696 402319
rect 191746 400208 191802 400217
rect 191746 400143 191802 400152
rect 191760 398886 191788 400143
rect 191748 398880 191800 398886
rect 191748 398822 191800 398828
rect 191746 397216 191802 397225
rect 191746 397151 191802 397160
rect 191760 396778 191788 397151
rect 191748 396772 191800 396778
rect 191748 396714 191800 396720
rect 191668 396630 191788 396658
rect 191484 396494 191696 396522
rect 191562 393136 191618 393145
rect 191562 393071 191618 393080
rect 191576 392086 191604 393071
rect 191564 392080 191616 392086
rect 191564 392022 191616 392028
rect 191564 315240 191616 315246
rect 191564 315182 191616 315188
rect 191380 305108 191432 305114
rect 191380 305050 191432 305056
rect 191392 296714 191420 305050
rect 191472 300824 191524 300830
rect 191472 300766 191524 300772
rect 191484 299713 191512 300766
rect 191470 299704 191526 299713
rect 191470 299639 191526 299648
rect 191392 296686 191512 296714
rect 191288 295384 191340 295390
rect 191288 295326 191340 295332
rect 191196 293956 191248 293962
rect 191196 293898 191248 293904
rect 191208 293321 191236 293898
rect 191194 293312 191250 293321
rect 191194 293247 191250 293256
rect 191300 292233 191328 295326
rect 191286 292224 191342 292233
rect 191286 292159 191342 292168
rect 191102 286784 191158 286793
rect 191102 286719 191158 286728
rect 190458 282432 190514 282441
rect 190458 282367 190514 282376
rect 190472 281586 190500 282367
rect 190460 281580 190512 281586
rect 190460 281522 190512 281528
rect 190550 281344 190606 281353
rect 190550 281279 190606 281288
rect 190564 280906 190592 281279
rect 190552 280900 190604 280906
rect 190552 280842 190604 280848
rect 190460 280084 190512 280090
rect 190460 280026 190512 280032
rect 190472 279177 190500 280026
rect 190458 279168 190514 279177
rect 190458 279103 190514 279112
rect 190458 278080 190514 278089
rect 190458 278015 190460 278024
rect 190512 278015 190514 278024
rect 190460 277986 190512 277992
rect 190458 276992 190514 277001
rect 190458 276927 190514 276936
rect 190472 276078 190500 276927
rect 190460 276072 190512 276078
rect 190460 276014 190512 276020
rect 190458 275904 190514 275913
rect 190458 275839 190514 275848
rect 190472 274718 190500 275839
rect 190550 274816 190606 274825
rect 190550 274751 190552 274760
rect 190604 274751 190606 274760
rect 190552 274722 190604 274728
rect 190460 274712 190512 274718
rect 190460 274654 190512 274660
rect 190458 273728 190514 273737
rect 190458 273663 190514 273672
rect 190472 273290 190500 273663
rect 190460 273284 190512 273290
rect 190460 273226 190512 273232
rect 190826 272640 190882 272649
rect 190826 272575 190882 272584
rect 190840 271930 190868 272575
rect 190828 271924 190880 271930
rect 190828 271866 190880 271872
rect 190826 270464 190882 270473
rect 190826 270399 190882 270408
rect 190840 269142 190868 270399
rect 190828 269136 190880 269142
rect 190828 269078 190880 269084
rect 190828 265056 190880 265062
rect 190826 265024 190828 265033
rect 190880 265024 190882 265033
rect 190826 264959 190882 264968
rect 190460 258120 190512 258126
rect 190458 258088 190460 258097
rect 190512 258088 190514 258097
rect 190458 258023 190514 258032
rect 190642 256320 190698 256329
rect 190642 256255 190698 256264
rect 190656 255338 190684 256255
rect 190644 255332 190696 255338
rect 190644 255274 190696 255280
rect 190368 251864 190420 251870
rect 190368 251806 190420 251812
rect 190642 250880 190698 250889
rect 190642 250815 190698 250824
rect 190656 249830 190684 250815
rect 190644 249824 190696 249830
rect 190644 249766 190696 249772
rect 190826 249792 190882 249801
rect 190826 249727 190882 249736
rect 190840 248470 190868 249727
rect 190828 248464 190880 248470
rect 190828 248406 190880 248412
rect 190276 245608 190328 245614
rect 190276 245550 190328 245556
rect 189998 242992 190054 243001
rect 189998 242927 190054 242936
rect 190012 236609 190040 242927
rect 189998 236600 190054 236609
rect 189998 236535 190054 236544
rect 189906 235240 189962 235249
rect 189906 235175 189962 235184
rect 189814 233064 189870 233073
rect 189814 232999 189870 233008
rect 189722 217288 189778 217297
rect 189722 217223 189778 217232
rect 189724 171896 189776 171902
rect 189724 171838 189776 171844
rect 188434 166424 188490 166433
rect 188434 166359 188490 166368
rect 188448 143585 188476 166359
rect 189736 164218 189764 171838
rect 189080 164212 189132 164218
rect 189080 164154 189132 164160
rect 189724 164212 189776 164218
rect 189724 164154 189776 164160
rect 189092 163538 189120 164154
rect 189080 163532 189132 163538
rect 189080 163474 189132 163480
rect 188618 155272 188674 155281
rect 188618 155207 188674 155216
rect 188526 145072 188582 145081
rect 188526 145007 188582 145016
rect 188434 143576 188490 143585
rect 188434 143511 188490 143520
rect 188448 133890 188476 143511
rect 188540 135182 188568 145007
rect 188632 144265 188660 155207
rect 188618 144256 188674 144265
rect 188618 144191 188674 144200
rect 188528 135176 188580 135182
rect 188528 135118 188580 135124
rect 188436 133884 188488 133890
rect 188436 133826 188488 133832
rect 189092 128450 189120 163474
rect 190366 155272 190422 155281
rect 190366 155207 190422 155216
rect 190274 134192 190330 134201
rect 190274 134127 190330 134136
rect 190288 129849 190316 134127
rect 190274 129840 190330 129849
rect 190274 129775 190330 129784
rect 189080 128444 189132 128450
rect 189080 128386 189132 128392
rect 188988 120216 189040 120222
rect 188988 120158 189040 120164
rect 188344 117224 188396 117230
rect 188344 117166 188396 117172
rect 188252 113212 188304 113218
rect 188252 113154 188304 113160
rect 187700 110492 187752 110498
rect 187700 110434 187752 110440
rect 187712 108322 187740 110434
rect 188264 109750 188292 113154
rect 188896 110560 188948 110566
rect 188896 110502 188948 110508
rect 188252 109744 188304 109750
rect 188252 109686 188304 109692
rect 187700 108316 187752 108322
rect 187700 108258 187752 108264
rect 188066 96928 188122 96937
rect 188066 96863 188122 96872
rect 188080 92041 188108 96863
rect 188344 95260 188396 95266
rect 188344 95202 188396 95208
rect 188066 92032 188122 92041
rect 188066 91967 188122 91976
rect 188356 84153 188384 95202
rect 188342 84144 188398 84153
rect 188342 84079 188398 84088
rect 188908 75886 188936 110502
rect 189000 78577 189028 120158
rect 189078 110800 189134 110809
rect 189078 110735 189134 110744
rect 189092 109002 189120 110735
rect 189080 108996 189132 109002
rect 189080 108938 189132 108944
rect 190276 105596 190328 105602
rect 190276 105538 190328 105544
rect 190182 94480 190238 94489
rect 190182 94415 190238 94424
rect 188986 78568 189042 78577
rect 188986 78503 189042 78512
rect 190196 77994 190224 94415
rect 190184 77988 190236 77994
rect 190184 77930 190236 77936
rect 188896 75880 188948 75886
rect 188896 75822 188948 75828
rect 187608 65544 187660 65550
rect 187608 65486 187660 65492
rect 186964 51740 187016 51746
rect 186964 51682 187016 51688
rect 190288 44878 190316 105538
rect 190380 85513 190408 155207
rect 191116 152522 191144 286719
rect 191300 279478 191328 292159
rect 191484 280265 191512 296686
rect 191576 296585 191604 315182
rect 191562 296576 191618 296585
rect 191562 296511 191618 296520
rect 191576 296070 191604 296511
rect 191564 296064 191616 296070
rect 191564 296006 191616 296012
rect 191668 290057 191696 396494
rect 191760 381546 191788 396630
rect 191748 381540 191800 381546
rect 191748 381482 191800 381488
rect 191746 378992 191802 379001
rect 191746 378927 191802 378936
rect 191760 373289 191788 378927
rect 191746 373280 191802 373289
rect 191746 373215 191802 373224
rect 191746 372872 191802 372881
rect 191746 372807 191802 372816
rect 191760 367713 191788 372807
rect 191746 367704 191802 367713
rect 191746 367639 191802 367648
rect 192496 327758 192524 436591
rect 192588 380322 192616 450502
rect 192680 447953 192708 455631
rect 193312 452804 193364 452810
rect 193312 452746 193364 452752
rect 192666 447944 192722 447953
rect 192666 447879 192722 447888
rect 193126 445088 193182 445097
rect 193126 445023 193182 445032
rect 192668 398948 192720 398954
rect 192668 398890 192720 398896
rect 192680 387122 192708 398890
rect 192668 387116 192720 387122
rect 192668 387058 192720 387064
rect 192576 380316 192628 380322
rect 192576 380258 192628 380264
rect 193140 370569 193168 445023
rect 193324 439550 193352 452746
rect 193416 449206 193444 456826
rect 194690 453112 194746 453121
rect 194690 453047 194746 453056
rect 194704 450228 194732 453047
rect 195164 450242 195192 460906
rect 195796 458312 195848 458318
rect 195794 458280 195796 458289
rect 195848 458280 195850 458289
rect 195794 458215 195850 458224
rect 197360 455524 197412 455530
rect 197360 455466 197412 455472
rect 195980 453348 196032 453354
rect 195980 453290 196032 453296
rect 195992 452985 196020 453290
rect 195978 452976 196034 452985
rect 195978 452911 196034 452920
rect 196532 452668 196584 452674
rect 196532 452610 196584 452616
rect 195164 450214 195638 450242
rect 196544 450228 196572 452610
rect 197372 450242 197400 455466
rect 197910 454200 197966 454209
rect 197910 454135 197966 454144
rect 197924 450242 197952 454135
rect 200120 454096 200172 454102
rect 200120 454038 200172 454044
rect 199292 451308 199344 451314
rect 199292 451250 199344 451256
rect 197372 450214 197478 450242
rect 197924 450214 198398 450242
rect 199304 450228 199332 451250
rect 200132 450242 200160 454038
rect 201788 450242 201816 460906
rect 203154 453112 203210 453121
rect 203154 453047 203210 453056
rect 200132 450214 200422 450242
rect 201788 450214 202262 450242
rect 203168 450228 203196 453047
rect 203628 450242 203656 460906
rect 208400 459604 208452 459610
rect 208400 459546 208452 459552
rect 207570 457056 207626 457065
rect 207570 456991 207626 457000
rect 204536 456816 204588 456822
rect 204536 456758 204588 456764
rect 204548 450242 204576 456758
rect 207110 454336 207166 454345
rect 207110 454271 207166 454280
rect 205914 452840 205970 452849
rect 205914 452775 205970 452784
rect 203628 450214 204102 450242
rect 204548 450214 205022 450242
rect 205928 450228 205956 452775
rect 207124 450242 207152 454271
rect 207046 450214 207152 450242
rect 207584 450242 207612 456991
rect 208412 450242 208440 459546
rect 210422 458416 210478 458425
rect 210422 458351 210478 458360
rect 209778 451480 209834 451489
rect 209778 451415 209834 451424
rect 207584 450214 207966 450242
rect 208412 450214 208886 450242
rect 209792 450228 209820 451415
rect 210436 451314 210464 458351
rect 212448 453348 212500 453354
rect 212448 453290 212500 453296
rect 212460 452713 212488 453290
rect 212446 452704 212502 452713
rect 211252 452668 211304 452674
rect 212446 452639 212502 452648
rect 211252 452610 211304 452616
rect 210424 451308 210476 451314
rect 210424 451250 210476 451256
rect 210436 450242 210464 451250
rect 211264 450566 211292 452610
rect 211618 451888 211674 451897
rect 211618 451823 211674 451832
rect 211252 450560 211304 450566
rect 211252 450502 211304 450508
rect 210436 450214 210726 450242
rect 211632 450228 211660 451823
rect 212644 450242 212672 462402
rect 212722 455696 212778 455705
rect 212722 455631 212778 455640
rect 212736 453422 212764 455631
rect 214576 455569 214604 703258
rect 215944 702636 215996 702642
rect 215944 702578 215996 702584
rect 215956 462330 215984 702578
rect 218992 698970 219020 703520
rect 235184 702710 235212 703520
rect 240784 703248 240836 703254
rect 240784 703190 240836 703196
rect 235172 702704 235224 702710
rect 235172 702646 235224 702652
rect 220084 700324 220136 700330
rect 220084 700266 220136 700272
rect 218980 698964 219032 698970
rect 218980 698906 219032 698912
rect 215392 462324 215444 462330
rect 215392 462266 215444 462272
rect 215944 462324 215996 462330
rect 215944 462266 215996 462272
rect 215404 461038 215432 462266
rect 215392 461032 215444 461038
rect 215392 460974 215444 460980
rect 215404 460934 215432 460974
rect 215404 460906 215984 460934
rect 214562 455560 214618 455569
rect 214562 455495 214618 455504
rect 212724 453416 212776 453422
rect 212724 453358 212776 453364
rect 213644 452804 213696 452810
rect 213644 452746 213696 452752
rect 212644 450214 212750 450242
rect 213656 450228 213684 452746
rect 214576 451274 214604 455495
rect 215484 453416 215536 453422
rect 215484 453358 215536 453364
rect 214116 451246 214604 451274
rect 214116 450242 214144 451246
rect 214116 450214 214590 450242
rect 215496 450228 215524 453358
rect 215956 450242 215984 460906
rect 220096 459649 220124 700266
rect 238024 474768 238076 474774
rect 238024 474710 238076 474716
rect 226984 473408 227036 473414
rect 226984 473350 227036 473356
rect 216862 459640 216918 459649
rect 216862 459575 216918 459584
rect 220082 459640 220138 459649
rect 226996 459610 227024 473350
rect 231860 472048 231912 472054
rect 231860 471990 231912 471996
rect 227812 467968 227864 467974
rect 227812 467910 227864 467916
rect 220082 459575 220138 459584
rect 226984 459604 227036 459610
rect 216876 450242 216904 459575
rect 226984 459546 227036 459552
rect 227628 459604 227680 459610
rect 227628 459546 227680 459552
rect 219806 457056 219862 457065
rect 219806 456991 219862 457000
rect 218980 456884 219032 456890
rect 218980 456826 219032 456832
rect 218152 454164 218204 454170
rect 218152 454106 218204 454112
rect 218164 450242 218192 454106
rect 218992 450242 219020 456826
rect 219820 450242 219848 456991
rect 220818 455560 220874 455569
rect 220818 455495 220874 455504
rect 225512 455524 225564 455530
rect 215956 450214 216430 450242
rect 216876 450214 217350 450242
rect 218164 450214 218454 450242
rect 218992 450214 219374 450242
rect 219820 450214 220294 450242
rect 220832 449993 220860 455495
rect 225512 455466 225564 455472
rect 222568 454096 222620 454102
rect 222568 454038 222620 454044
rect 222108 452736 222160 452742
rect 222108 452678 222160 452684
rect 222120 450228 222148 452678
rect 222580 450242 222608 454038
rect 225050 453248 225106 453257
rect 225050 453183 225106 453192
rect 224130 452704 224186 452713
rect 224130 452639 224186 452648
rect 222580 450214 223054 450242
rect 224144 450228 224172 452639
rect 225064 450228 225092 453183
rect 225524 450242 225552 455466
rect 227640 454034 227668 459546
rect 227720 458312 227772 458318
rect 227720 458254 227772 458260
rect 227628 454028 227680 454034
rect 227628 453970 227680 453976
rect 227732 452674 227760 458254
rect 226892 452668 226944 452674
rect 226892 452610 226944 452616
rect 227720 452668 227772 452674
rect 227720 452610 227772 452616
rect 225524 450214 225998 450242
rect 226904 450228 226932 452610
rect 227824 450242 227852 467910
rect 230480 456816 230532 456822
rect 230480 456758 230532 456764
rect 228732 454028 228784 454034
rect 228732 453970 228784 453976
rect 228086 450392 228142 450401
rect 228086 450327 228142 450336
rect 228100 450242 228128 450327
rect 227824 450228 228128 450242
rect 228744 450228 228772 453970
rect 229652 452668 229704 452674
rect 229652 452610 229704 452616
rect 229664 450228 229692 452610
rect 230492 450265 230520 456758
rect 231214 454200 231270 454209
rect 231214 454135 231270 454144
rect 230478 450256 230534 450265
rect 227838 450214 228128 450228
rect 231228 450242 231256 454135
rect 230534 450214 230782 450242
rect 231228 450214 231702 450242
rect 230478 450191 230534 450200
rect 231872 450022 231900 471990
rect 237380 458312 237432 458318
rect 237380 458254 237432 458260
rect 233238 455696 233294 455705
rect 233238 455631 233294 455640
rect 233252 455462 233280 455631
rect 233240 455456 233292 455462
rect 233240 455398 233292 455404
rect 233252 450242 233280 455398
rect 234894 454064 234950 454073
rect 234894 453999 234950 454008
rect 234434 452704 234490 452713
rect 234434 452639 234490 452648
rect 233252 450214 233542 450242
rect 234448 450228 234476 452639
rect 234908 450242 234936 453999
rect 237392 453257 237420 458254
rect 238036 456074 238064 474710
rect 240796 471986 240824 703190
rect 249064 703180 249116 703186
rect 249064 703122 249116 703128
rect 241520 698964 241572 698970
rect 241520 698906 241572 698912
rect 240140 471980 240192 471986
rect 240140 471922 240192 471928
rect 240784 471980 240836 471986
rect 240784 471922 240836 471928
rect 240152 471306 240180 471922
rect 240140 471300 240192 471306
rect 240140 471242 240192 471248
rect 240152 460193 240180 471242
rect 241532 469878 241560 698906
rect 249076 476134 249104 703122
rect 258724 702704 258776 702710
rect 258724 702646 258776 702652
rect 258736 481642 258764 702646
rect 267660 700330 267688 703520
rect 283852 703458 283880 703520
rect 283840 703452 283892 703458
rect 283840 703394 283892 703400
rect 282828 703384 282880 703390
rect 282828 703326 282880 703332
rect 273904 703112 273956 703118
rect 273904 703054 273956 703060
rect 271144 702976 271196 702982
rect 271144 702918 271196 702924
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 258172 481636 258224 481642
rect 258172 481578 258224 481584
rect 258724 481636 258776 481642
rect 258724 481578 258776 481584
rect 258184 480282 258212 481578
rect 258172 480276 258224 480282
rect 258172 480218 258224 480224
rect 251824 478916 251876 478922
rect 251824 478858 251876 478864
rect 249064 476128 249116 476134
rect 249064 476070 249116 476076
rect 241520 469872 241572 469878
rect 241520 469814 241572 469820
rect 241532 469334 241560 469814
rect 241520 469328 241572 469334
rect 241520 469270 241572 469276
rect 242164 469328 242216 469334
rect 242164 469270 242216 469276
rect 240138 460184 240194 460193
rect 240138 460119 240194 460128
rect 240152 459649 240180 460119
rect 238758 459640 238814 459649
rect 238758 459575 238814 459584
rect 240138 459640 240194 459649
rect 240138 459575 240194 459584
rect 238024 456068 238076 456074
rect 238024 456010 238076 456016
rect 237378 453248 237434 453257
rect 237378 453183 237434 453192
rect 237380 452668 237432 452674
rect 237380 452610 237432 452616
rect 236734 451888 236790 451897
rect 236734 451823 236790 451832
rect 236748 450242 236776 451823
rect 234908 450214 235382 450242
rect 236486 450214 236776 450242
rect 237392 450228 237420 452610
rect 238772 450242 238800 459575
rect 241520 456068 241572 456074
rect 241520 456010 241572 456016
rect 240232 451444 240284 451450
rect 240232 451386 240284 451392
rect 240244 450242 240272 451386
rect 241060 451376 241112 451382
rect 241060 451318 241112 451324
rect 238772 450214 239246 450242
rect 240166 450214 240272 450242
rect 241072 450228 241100 451318
rect 231860 450016 231912 450022
rect 220818 449984 220874 449993
rect 200960 449942 201342 449970
rect 200960 449886 200988 449942
rect 220874 449942 221214 449970
rect 232872 450016 232924 450022
rect 231860 449958 231912 449964
rect 232622 449964 232872 449970
rect 238482 449984 238538 449993
rect 232622 449958 232924 449964
rect 232622 449942 232912 449958
rect 238326 449942 238482 449970
rect 220818 449919 220874 449928
rect 240244 449954 240272 450214
rect 241532 449970 241560 456010
rect 242176 453937 242204 469270
rect 242900 466540 242952 466546
rect 242900 466482 242952 466488
rect 242162 453928 242218 453937
rect 242162 453863 242218 453872
rect 242912 450242 242940 466482
rect 245660 465112 245712 465118
rect 245660 465054 245712 465060
rect 245672 460934 245700 465054
rect 249076 460934 249104 476070
rect 251180 470620 251232 470626
rect 251180 470562 251232 470568
rect 245672 460906 246344 460934
rect 249076 460906 249288 460934
rect 244002 453928 244058 453937
rect 244002 453863 244058 453872
rect 244016 452985 244044 453863
rect 244002 452976 244058 452985
rect 244002 452911 244058 452920
rect 242912 450214 243110 450242
rect 244016 450228 244044 452911
rect 246316 450242 246344 460906
rect 249260 458289 249288 460906
rect 249246 458280 249302 458289
rect 249246 458215 249302 458224
rect 247866 451344 247922 451353
rect 247866 451279 247922 451288
rect 246316 450214 246790 450242
rect 247880 450228 247908 451279
rect 249260 450242 249288 458215
rect 250626 456920 250682 456929
rect 250626 456855 250682 456864
rect 250640 452713 250668 456855
rect 251192 456142 251220 470562
rect 251180 456136 251232 456142
rect 251180 456078 251232 456084
rect 251836 452810 251864 478858
rect 255412 469260 255464 469266
rect 255412 469202 255464 469208
rect 252560 466472 252612 466478
rect 252560 466414 252612 466420
rect 252572 460934 252600 466414
rect 255320 463820 255372 463826
rect 255320 463762 255372 463768
rect 253938 461000 253994 461009
rect 253938 460935 253994 460944
rect 252572 460906 252968 460934
rect 252100 456136 252152 456142
rect 252100 456078 252152 456084
rect 251824 452804 251876 452810
rect 251824 452746 251876 452752
rect 251456 452736 251508 452742
rect 250626 452704 250682 452713
rect 251456 452678 251508 452684
rect 250626 452639 250682 452648
rect 249260 450214 249734 450242
rect 250640 450228 250668 452639
rect 244554 450120 244610 450129
rect 244610 450078 244950 450106
rect 244554 450055 244610 450064
rect 248510 449984 248566 449993
rect 241532 449954 242480 449970
rect 238482 449919 238538 449928
rect 240232 449948 240284 449954
rect 241532 449948 242492 449954
rect 241532 449942 242440 449948
rect 240232 449890 240284 449896
rect 248566 449942 248814 449970
rect 248510 449919 248566 449928
rect 242440 449890 242492 449896
rect 200948 449880 201000 449886
rect 200948 449822 201000 449828
rect 251468 449750 251496 452678
rect 251836 450242 251864 452746
rect 251574 450214 251864 450242
rect 252112 450242 252140 456078
rect 252940 450242 252968 460906
rect 252112 450214 252494 450242
rect 252940 450214 253414 450242
rect 251456 449744 251508 449750
rect 193494 449712 193550 449721
rect 245750 449712 245806 449721
rect 193550 449670 193614 449698
rect 193494 449647 193550 449656
rect 245806 449670 245870 449698
rect 251456 449686 251508 449692
rect 245750 449647 245806 449656
rect 193404 449200 193456 449206
rect 193404 449142 193456 449148
rect 253952 446185 253980 460935
rect 254584 449948 254636 449954
rect 254584 449890 254636 449896
rect 253938 446176 253994 446185
rect 253938 446111 253994 446120
rect 253938 440464 253994 440473
rect 253938 440399 253994 440408
rect 193312 439544 193364 439550
rect 193312 439486 193364 439492
rect 253570 402112 253626 402121
rect 253570 402047 253626 402056
rect 253584 393314 253612 402047
rect 253492 393286 253612 393314
rect 193404 392012 193456 392018
rect 193404 391954 193456 391960
rect 193416 380798 193444 391954
rect 193494 390960 193550 390969
rect 252558 390960 252614 390969
rect 193550 390918 193614 390946
rect 193494 390895 193550 390904
rect 252558 390895 252614 390904
rect 223486 390824 223542 390833
rect 223486 390759 223542 390768
rect 196912 390658 197294 390674
rect 196900 390652 197294 390658
rect 196952 390646 197294 390652
rect 196900 390594 196952 390600
rect 223500 390402 223528 390759
rect 194520 389065 194548 390388
rect 195440 389201 195468 390388
rect 195992 390374 196374 390402
rect 197372 390374 198214 390402
rect 198752 390374 199134 390402
rect 200132 390374 200238 390402
rect 195426 389192 195482 389201
rect 195426 389127 195482 389136
rect 194506 389056 194562 389065
rect 194506 388991 194562 389000
rect 194600 381608 194652 381614
rect 194600 381550 194652 381556
rect 193404 380792 193456 380798
rect 193404 380734 193456 380740
rect 193126 370560 193182 370569
rect 193126 370495 193182 370504
rect 193404 363792 193456 363798
rect 193404 363734 193456 363740
rect 193416 363662 193444 363734
rect 193404 363656 193456 363662
rect 193404 363598 193456 363604
rect 193312 355360 193364 355366
rect 193312 355302 193364 355308
rect 192576 328568 192628 328574
rect 192576 328510 192628 328516
rect 192484 327752 192536 327758
rect 192484 327694 192536 327700
rect 192484 316124 192536 316130
rect 192484 316066 192536 316072
rect 192496 300966 192524 316066
rect 192588 315081 192616 328510
rect 193128 320952 193180 320958
rect 193128 320894 193180 320900
rect 192574 315072 192630 315081
rect 192574 315007 192630 315016
rect 192666 313984 192722 313993
rect 192666 313919 192722 313928
rect 192680 302938 192708 313919
rect 192668 302932 192720 302938
rect 192668 302874 192720 302880
rect 192576 302320 192628 302326
rect 192576 302262 192628 302268
rect 192484 300960 192536 300966
rect 192484 300902 192536 300908
rect 191746 299840 191802 299849
rect 191746 299775 191802 299784
rect 191760 299538 191788 299775
rect 191748 299532 191800 299538
rect 191748 299474 191800 299480
rect 191748 298104 191800 298110
rect 191748 298046 191800 298052
rect 191760 297673 191788 298046
rect 191746 297664 191802 297673
rect 191746 297599 191802 297608
rect 191746 291136 191802 291145
rect 191746 291071 191802 291080
rect 191654 290048 191710 290057
rect 191654 289983 191710 289992
rect 191760 289882 191788 291071
rect 191748 289876 191800 289882
rect 191748 289818 191800 289824
rect 191656 289808 191708 289814
rect 191656 289750 191708 289756
rect 191668 288969 191696 289750
rect 191654 288960 191710 288969
rect 191654 288895 191710 288904
rect 191838 288416 191894 288425
rect 191838 288351 191894 288360
rect 191746 287872 191802 287881
rect 191746 287807 191802 287816
rect 191760 287774 191788 287807
rect 191748 287768 191800 287774
rect 191748 287710 191800 287716
rect 191746 284608 191802 284617
rect 191746 284543 191802 284552
rect 191760 284374 191788 284543
rect 191748 284368 191800 284374
rect 191748 284310 191800 284316
rect 191748 284232 191800 284238
rect 191748 284174 191800 284180
rect 191760 283529 191788 284174
rect 191746 283520 191802 283529
rect 191746 283455 191802 283464
rect 191852 282198 191880 288351
rect 191840 282192 191892 282198
rect 191840 282134 191892 282140
rect 191746 281344 191802 281353
rect 191746 281279 191802 281288
rect 191470 280256 191526 280265
rect 191470 280191 191526 280200
rect 191288 279472 191340 279478
rect 191288 279414 191340 279420
rect 191484 273254 191512 280191
rect 191208 273226 191512 273254
rect 191208 167686 191236 273226
rect 191654 271552 191710 271561
rect 191654 271487 191710 271496
rect 191668 270638 191696 271487
rect 191656 270632 191708 270638
rect 191656 270574 191708 270580
rect 191562 269376 191618 269385
rect 191562 269311 191618 269320
rect 191576 269210 191604 269311
rect 191564 269204 191616 269210
rect 191564 269146 191616 269152
rect 191654 268288 191710 268297
rect 191654 268223 191710 268232
rect 191668 267782 191696 268223
rect 191656 267776 191708 267782
rect 191656 267718 191708 267724
rect 191654 266112 191710 266121
rect 191654 266047 191710 266056
rect 191668 264994 191696 266047
rect 191656 264988 191708 264994
rect 191656 264930 191708 264936
rect 191654 263936 191710 263945
rect 191654 263871 191710 263880
rect 191668 263634 191696 263871
rect 191656 263628 191708 263634
rect 191656 263570 191708 263576
rect 191654 262848 191710 262857
rect 191654 262783 191710 262792
rect 191668 262274 191696 262783
rect 191656 262268 191708 262274
rect 191656 262210 191708 262216
rect 191654 261760 191710 261769
rect 191654 261695 191710 261704
rect 191668 260914 191696 261695
rect 191656 260908 191708 260914
rect 191656 260850 191708 260856
rect 191654 260672 191710 260681
rect 191654 260607 191710 260616
rect 191668 259554 191696 260607
rect 191656 259548 191708 259554
rect 191656 259490 191708 259496
rect 191654 257408 191710 257417
rect 191654 257343 191710 257352
rect 191668 256766 191696 257343
rect 191656 256760 191708 256766
rect 191656 256702 191708 256708
rect 191654 255232 191710 255241
rect 191654 255167 191710 255176
rect 191562 254144 191618 254153
rect 191562 254079 191618 254088
rect 191576 253978 191604 254079
rect 191668 254046 191696 255167
rect 191656 254040 191708 254046
rect 191656 253982 191708 253988
rect 191564 253972 191616 253978
rect 191564 253914 191616 253920
rect 191654 253056 191710 253065
rect 191654 252991 191710 253000
rect 191668 252618 191696 252991
rect 191656 252612 191708 252618
rect 191656 252554 191708 252560
rect 191654 251968 191710 251977
rect 191654 251903 191710 251912
rect 191668 251258 191696 251903
rect 191656 251252 191708 251258
rect 191656 251194 191708 251200
rect 191288 245676 191340 245682
rect 191288 245618 191340 245624
rect 191300 235958 191328 245618
rect 191760 238105 191788 281279
rect 191840 245608 191892 245614
rect 191840 245550 191892 245556
rect 191746 238096 191802 238105
rect 191746 238031 191802 238040
rect 191288 235952 191340 235958
rect 191288 235894 191340 235900
rect 191196 167680 191248 167686
rect 191196 167622 191248 167628
rect 191656 160132 191708 160138
rect 191656 160074 191708 160080
rect 191564 155916 191616 155922
rect 191564 155858 191616 155864
rect 190460 152516 190512 152522
rect 190460 152458 190512 152464
rect 191104 152516 191156 152522
rect 191104 152458 191156 152464
rect 191196 152516 191248 152522
rect 191196 152458 191248 152464
rect 190472 132494 190500 152458
rect 190472 132466 190592 132494
rect 190564 118697 190592 132466
rect 191208 132462 191236 152458
rect 191196 132456 191248 132462
rect 191196 132398 191248 132404
rect 191010 130112 191066 130121
rect 191010 130047 191066 130056
rect 191024 129810 191052 130047
rect 191012 129804 191064 129810
rect 191012 129746 191064 129752
rect 191208 129305 191236 132398
rect 191194 129296 191250 129305
rect 191194 129231 191250 129240
rect 191472 129056 191524 129062
rect 191472 128998 191524 129004
rect 191194 128480 191250 128489
rect 191194 128415 191196 128424
rect 191248 128415 191250 128424
rect 191196 128386 191248 128392
rect 191012 124160 191064 124166
rect 191012 124102 191064 124108
rect 191024 123049 191052 124102
rect 191484 123865 191512 128998
rect 191576 126585 191604 155858
rect 191668 139913 191696 160074
rect 191748 157412 191800 157418
rect 191748 157354 191800 157360
rect 191760 155922 191788 157354
rect 191748 155916 191800 155922
rect 191748 155858 191800 155864
rect 191852 148374 191880 245550
rect 192496 242962 192524 300902
rect 192588 291009 192616 302262
rect 192574 291000 192630 291009
rect 192574 290935 192630 290944
rect 193140 285705 193168 320894
rect 193218 315072 193274 315081
rect 193218 315007 193274 315016
rect 193232 303686 193260 315007
rect 193324 305114 193352 355302
rect 193312 305108 193364 305114
rect 193312 305050 193364 305056
rect 193220 303680 193272 303686
rect 193220 303622 193272 303628
rect 193312 301096 193364 301102
rect 193310 301064 193312 301073
rect 193364 301064 193366 301073
rect 193310 300999 193366 301008
rect 193416 295390 193444 363598
rect 194612 352578 194640 381550
rect 195992 363798 196020 390374
rect 196072 390312 196124 390318
rect 196072 390254 196124 390260
rect 196084 369238 196112 390254
rect 197372 385121 197400 390374
rect 198004 385688 198056 385694
rect 198004 385630 198056 385636
rect 197358 385112 197414 385121
rect 197358 385047 197414 385056
rect 197372 383625 197400 385047
rect 197358 383616 197414 383625
rect 197358 383551 197414 383560
rect 198016 372502 198044 385630
rect 198752 380934 198780 390374
rect 198740 380928 198792 380934
rect 198740 380870 198792 380876
rect 198752 380769 198780 380870
rect 198738 380760 198794 380769
rect 198738 380695 198794 380704
rect 200132 380225 200160 390374
rect 201144 388521 201172 390388
rect 201512 390374 202078 390402
rect 202892 390374 202998 390402
rect 201130 388512 201186 388521
rect 201130 388447 201186 388456
rect 200210 385792 200266 385801
rect 200210 385727 200266 385736
rect 200224 380905 200252 385727
rect 200210 380896 200266 380905
rect 200210 380831 200266 380840
rect 200118 380216 200174 380225
rect 200118 380151 200174 380160
rect 198004 372496 198056 372502
rect 198004 372438 198056 372444
rect 196072 369232 196124 369238
rect 196072 369174 196124 369180
rect 201512 367810 201540 390374
rect 202142 380760 202198 380769
rect 202142 380695 202198 380704
rect 201500 367804 201552 367810
rect 201500 367746 201552 367752
rect 195980 363792 196032 363798
rect 195980 363734 196032 363740
rect 194600 352572 194652 352578
rect 194600 352514 194652 352520
rect 195244 349920 195296 349926
rect 195244 349862 195296 349868
rect 195256 315246 195284 349862
rect 196624 348424 196676 348430
rect 196624 348366 196676 348372
rect 195244 315240 195296 315246
rect 195244 315182 195296 315188
rect 193496 305108 193548 305114
rect 193496 305050 193548 305056
rect 193508 299033 193536 305050
rect 196256 303748 196308 303754
rect 196256 303690 196308 303696
rect 193588 303680 193640 303686
rect 193588 303622 193640 303628
rect 193600 301594 193628 303622
rect 193600 301566 193890 301594
rect 196268 301580 196296 303690
rect 196636 303657 196664 348366
rect 202156 344321 202184 380695
rect 202892 355366 202920 390374
rect 203904 385694 203932 390388
rect 204272 390374 204838 390402
rect 205652 390374 205942 390402
rect 203892 385688 203944 385694
rect 203892 385630 203944 385636
rect 204272 372065 204300 390374
rect 205546 389328 205602 389337
rect 205546 389263 205602 389272
rect 205560 387841 205588 389263
rect 205546 387832 205602 387841
rect 205546 387767 205602 387776
rect 204350 381576 204406 381585
rect 204350 381511 204406 381520
rect 204258 372056 204314 372065
rect 204258 371991 204314 372000
rect 204272 367062 204300 371991
rect 204260 367056 204312 367062
rect 204260 366998 204312 367004
rect 202880 355360 202932 355366
rect 202880 355302 202932 355308
rect 202142 344312 202198 344321
rect 202142 344247 202198 344256
rect 204260 343664 204312 343670
rect 204260 343606 204312 343612
rect 199382 331256 199438 331265
rect 199382 331191 199438 331200
rect 198830 322960 198886 322969
rect 198830 322895 198886 322904
rect 197452 317552 197504 317558
rect 197452 317494 197504 317500
rect 197358 306776 197414 306785
rect 197358 306711 197414 306720
rect 197372 306406 197400 306711
rect 197360 306400 197412 306406
rect 197360 306342 197412 306348
rect 197358 305280 197414 305289
rect 197358 305215 197414 305224
rect 196622 303648 196678 303657
rect 196622 303583 196678 303592
rect 197372 302938 197400 305215
rect 197360 302932 197412 302938
rect 197360 302874 197412 302880
rect 196806 302288 196862 302297
rect 196806 302223 196862 302232
rect 196820 301580 196848 302223
rect 197464 301580 197492 317494
rect 197910 306504 197966 306513
rect 197910 306439 197966 306448
rect 197924 302841 197952 306439
rect 197910 302832 197966 302841
rect 197910 302767 197966 302776
rect 198004 302252 198056 302258
rect 198004 302194 198056 302200
rect 198016 301580 198044 302194
rect 198844 301594 198872 322895
rect 199396 307086 199424 331191
rect 201682 329896 201738 329905
rect 201682 329831 201738 329840
rect 201696 325694 201724 329831
rect 201696 325666 201816 325694
rect 201590 307864 201646 307873
rect 201590 307799 201646 307808
rect 199384 307080 199436 307086
rect 199384 307022 199436 307028
rect 201038 302560 201094 302569
rect 201038 302495 201094 302504
rect 200394 302424 200450 302433
rect 200394 302359 200450 302368
rect 198844 301566 199226 301594
rect 200408 301580 200436 302359
rect 201052 301580 201080 302495
rect 201604 301580 201632 307799
rect 201788 301594 201816 325666
rect 203062 310584 203118 310593
rect 203062 310519 203118 310528
rect 202788 305108 202840 305114
rect 202788 305050 202840 305056
rect 201788 301566 202262 301594
rect 202800 301580 202828 305050
rect 203076 301594 203104 310519
rect 203984 307080 204036 307086
rect 203984 307022 204036 307028
rect 203076 301566 203458 301594
rect 203996 301580 204024 307022
rect 204272 301594 204300 343606
rect 204364 313993 204392 381511
rect 205560 345681 205588 387767
rect 205652 377466 205680 390374
rect 206848 387841 206876 390388
rect 207032 390374 207782 390402
rect 208412 390374 208702 390402
rect 208872 390374 209622 390402
rect 209792 390374 210542 390402
rect 211172 390374 211646 390402
rect 206834 387832 206890 387841
rect 206834 387767 206890 387776
rect 207032 379438 207060 390374
rect 207020 379432 207072 379438
rect 207020 379374 207072 379380
rect 205640 377460 205692 377466
rect 205640 377402 205692 377408
rect 205546 345672 205602 345681
rect 205546 345607 205602 345616
rect 208412 341562 208440 390374
rect 208872 373994 208900 390374
rect 208504 373966 208900 373994
rect 208504 373318 208532 373966
rect 208492 373312 208544 373318
rect 208492 373254 208544 373260
rect 209792 371890 209820 390374
rect 209780 371884 209832 371890
rect 209780 371826 209832 371832
rect 211172 354686 211200 390374
rect 211160 354680 211212 354686
rect 211160 354622 211212 354628
rect 211172 346526 211200 354622
rect 212552 354006 212580 390388
rect 213472 388385 213500 390388
rect 213932 390374 214406 390402
rect 213458 388376 213514 388385
rect 213458 388311 213514 388320
rect 213932 366382 213960 390374
rect 214562 387832 214618 387841
rect 214562 387767 214618 387776
rect 214012 387116 214064 387122
rect 214012 387058 214064 387064
rect 213920 366376 213972 366382
rect 213920 366318 213972 366324
rect 213826 363624 213882 363633
rect 213826 363559 213882 363568
rect 213840 361593 213868 363559
rect 213826 361584 213882 361593
rect 213826 361519 213882 361528
rect 212540 354000 212592 354006
rect 212540 353942 212592 353948
rect 211160 346520 211212 346526
rect 211160 346462 211212 346468
rect 211804 346520 211856 346526
rect 211804 346462 211856 346468
rect 208400 341556 208452 341562
rect 208400 341498 208452 341504
rect 205638 340912 205694 340921
rect 205638 340847 205694 340856
rect 204350 313984 204406 313993
rect 204350 313919 204406 313928
rect 204718 313440 204774 313449
rect 204718 313375 204774 313384
rect 204732 301594 204760 313375
rect 205652 301594 205680 340847
rect 205730 339552 205786 339561
rect 205730 339487 205786 339496
rect 205744 325694 205772 339487
rect 205744 325666 206048 325694
rect 206020 301594 206048 325666
rect 207110 321736 207166 321745
rect 207110 321671 207166 321680
rect 207124 301594 207152 321671
rect 209042 317792 209098 317801
rect 209042 317727 209098 317736
rect 208400 313404 208452 313410
rect 208400 313346 208452 313352
rect 208412 301594 208440 313346
rect 209056 302977 209084 317727
rect 211816 315353 211844 346462
rect 213182 334112 213238 334121
rect 213182 334047 213238 334056
rect 211802 315344 211858 315353
rect 211802 315279 211858 315288
rect 209778 314936 209834 314945
rect 209778 314871 209834 314880
rect 209042 302968 209098 302977
rect 209042 302903 209098 302912
rect 209792 301594 209820 314871
rect 211344 313336 211396 313342
rect 211344 313278 211396 313284
rect 210238 309496 210294 309505
rect 210238 309431 210294 309440
rect 210252 301594 210280 309431
rect 211356 303686 211384 313278
rect 211434 310720 211490 310729
rect 211434 310655 211490 310664
rect 211344 303680 211396 303686
rect 211344 303622 211396 303628
rect 211252 302932 211304 302938
rect 211252 302874 211304 302880
rect 204272 301566 204654 301594
rect 204732 301566 205206 301594
rect 205652 301566 205850 301594
rect 206020 301566 206402 301594
rect 207124 301566 207598 301594
rect 208412 301566 208886 301594
rect 209792 301566 210082 301594
rect 210252 301566 210634 301594
rect 211264 301580 211292 302874
rect 211448 301594 211476 310655
rect 213196 304298 213224 334047
rect 213274 330032 213330 330041
rect 213274 329967 213330 329976
rect 213288 305794 213316 329967
rect 214024 316810 214052 387058
rect 214576 365673 214604 387767
rect 214562 365664 214618 365673
rect 214562 365599 214618 365608
rect 215206 365664 215262 365673
rect 215206 365599 215262 365608
rect 215220 364993 215248 365599
rect 215206 364984 215262 364993
rect 215206 364919 215262 364928
rect 215220 363633 215248 364919
rect 215206 363624 215262 363633
rect 215206 363559 215262 363568
rect 215312 358766 215340 390388
rect 215404 390374 216246 390402
rect 216692 390374 217350 390402
rect 215404 359514 215432 390374
rect 216692 361554 216720 390374
rect 218256 387841 218284 390388
rect 218532 390374 219190 390402
rect 219452 390374 220110 390402
rect 218242 387832 218298 387841
rect 218242 387767 218298 387776
rect 218532 373994 218560 390374
rect 219452 383654 219480 390374
rect 221016 387190 221044 390388
rect 221292 390374 221950 390402
rect 222212 390374 222870 390402
rect 223500 390374 223974 390402
rect 224236 390374 224894 390402
rect 224972 390374 225814 390402
rect 226444 390374 226734 390402
rect 227272 390374 227654 390402
rect 227732 390374 228574 390402
rect 229112 390374 229678 390402
rect 230492 390374 230598 390402
rect 231228 390374 231518 390402
rect 231872 390374 232438 390402
rect 233252 390374 233358 390402
rect 221004 387184 221056 387190
rect 221004 387126 221056 387132
rect 219452 383626 219572 383654
rect 218072 373966 218560 373994
rect 216680 361548 216732 361554
rect 216680 361490 216732 361496
rect 215392 359508 215444 359514
rect 215392 359450 215444 359456
rect 215300 358760 215352 358766
rect 215300 358702 215352 358708
rect 215944 358760 215996 358766
rect 215944 358702 215996 358708
rect 215956 335354 215984 358702
rect 215864 335326 215984 335354
rect 215864 324465 215892 335326
rect 216034 327176 216090 327185
rect 216034 327111 216090 327120
rect 215942 325952 215998 325961
rect 215942 325887 215998 325896
rect 215850 324456 215906 324465
rect 215850 324391 215906 324400
rect 215300 319456 215352 319462
rect 215300 319398 215352 319404
rect 214012 316804 214064 316810
rect 214012 316746 214064 316752
rect 214564 316804 214616 316810
rect 214564 316746 214616 316752
rect 214576 316130 214604 316746
rect 215312 316742 215340 319398
rect 215300 316736 215352 316742
rect 215300 316678 215352 316684
rect 214564 316124 214616 316130
rect 214564 316066 214616 316072
rect 213642 308000 213698 308009
rect 213642 307935 213698 307944
rect 213276 305788 213328 305794
rect 213276 305730 213328 305736
rect 213184 304292 213236 304298
rect 213184 304234 213236 304240
rect 212998 303920 213054 303929
rect 212998 303855 213054 303864
rect 212172 303680 212224 303686
rect 212172 303622 212224 303628
rect 212184 301594 212212 303622
rect 211448 301566 211830 301594
rect 212184 301566 212474 301594
rect 213012 301580 213040 303855
rect 213656 301580 213684 307935
rect 214196 306468 214248 306474
rect 214196 306410 214248 306416
rect 214208 301580 214236 306410
rect 207938 301472 207994 301481
rect 207994 301430 208242 301458
rect 207938 301407 207994 301416
rect 198370 301336 198426 301345
rect 198426 301294 198674 301322
rect 198370 301271 198426 301280
rect 194230 301200 194286 301209
rect 194286 301158 194442 301186
rect 194230 301135 194286 301144
rect 195244 301096 195296 301102
rect 195296 301044 195638 301050
rect 195244 301038 195638 301044
rect 195256 301022 195638 301038
rect 206940 301034 207046 301050
rect 206928 301028 207046 301034
rect 206980 301022 207046 301028
rect 206928 300970 206980 300976
rect 214576 300966 214604 316066
rect 214838 305144 214894 305153
rect 214838 305079 214894 305088
rect 214852 301580 214880 305079
rect 215390 305008 215446 305017
rect 215390 304943 215446 304952
rect 215404 301580 215432 304943
rect 215956 303686 215984 325887
rect 216048 313954 216076 327111
rect 216692 320958 216720 361490
rect 216680 320952 216732 320958
rect 216680 320894 216732 320900
rect 216036 313948 216088 313954
rect 216036 313890 216088 313896
rect 218072 311166 218100 373966
rect 219544 362846 219572 383626
rect 221292 373994 221320 390374
rect 220924 373966 221320 373994
rect 220726 365800 220782 365809
rect 220726 365735 220782 365744
rect 220740 365702 220768 365735
rect 220728 365696 220780 365702
rect 220728 365638 220780 365644
rect 219532 362840 219584 362846
rect 219532 362782 219584 362788
rect 220084 362840 220136 362846
rect 220084 362782 220136 362788
rect 219438 332616 219494 332625
rect 219438 332551 219494 332560
rect 219452 325694 219480 332551
rect 220096 330449 220124 362782
rect 220924 356046 220952 373966
rect 220912 356040 220964 356046
rect 220912 355982 220964 355988
rect 221556 356040 221608 356046
rect 221556 355982 221608 355988
rect 221464 336796 221516 336802
rect 221464 336738 221516 336744
rect 220082 330440 220138 330449
rect 220082 330375 220138 330384
rect 219452 325666 219848 325694
rect 218702 314800 218758 314809
rect 218702 314735 218758 314744
rect 218060 311160 218112 311166
rect 218060 311102 218112 311108
rect 217416 310548 217468 310554
rect 217416 310490 217468 310496
rect 216036 307828 216088 307834
rect 216036 307770 216088 307776
rect 215944 303680 215996 303686
rect 215944 303622 215996 303628
rect 216048 301580 216076 307770
rect 216588 305040 216640 305046
rect 216588 304982 216640 304988
rect 216600 301580 216628 304982
rect 217232 303680 217284 303686
rect 217232 303622 217284 303628
rect 217244 301580 217272 303622
rect 217428 301594 217456 310490
rect 218518 309360 218574 309369
rect 218518 309295 218574 309304
rect 218428 302320 218480 302326
rect 218428 302262 218480 302268
rect 217428 301566 217810 301594
rect 218440 301580 218468 302262
rect 218532 301594 218560 309295
rect 218716 304978 218744 314735
rect 219622 306776 219678 306785
rect 219622 306711 219678 306720
rect 218704 304972 218756 304978
rect 218704 304914 218756 304920
rect 218532 301566 219006 301594
rect 219636 301580 219664 306711
rect 219820 301594 219848 325666
rect 220910 312080 220966 312089
rect 220910 312015 220966 312024
rect 220820 304972 220872 304978
rect 220820 304914 220872 304920
rect 219820 301566 220202 301594
rect 220832 301580 220860 304914
rect 220924 303686 220952 312015
rect 221002 311944 221058 311953
rect 221002 311879 221058 311888
rect 220912 303680 220964 303686
rect 220912 303622 220964 303628
rect 221016 301594 221044 311879
rect 221476 303754 221504 336738
rect 221568 333305 221596 355982
rect 222212 353326 222240 390374
rect 222200 353320 222252 353326
rect 222200 353262 222252 353268
rect 222844 352572 222896 352578
rect 222844 352514 222896 352520
rect 222290 335472 222346 335481
rect 222290 335407 222346 335416
rect 221554 333296 221610 333305
rect 221554 333231 221610 333240
rect 221464 303748 221516 303754
rect 221464 303690 221516 303696
rect 221740 303680 221792 303686
rect 221740 303622 221792 303628
rect 221752 301594 221780 303622
rect 222304 301594 222332 335407
rect 222856 305658 222884 352514
rect 223500 337414 223528 390374
rect 224236 373994 224264 390374
rect 224972 375290 225000 390374
rect 226340 387048 226392 387054
rect 226340 386990 226392 386996
rect 224960 375284 225012 375290
rect 224960 375226 225012 375232
rect 223592 373966 224264 373994
rect 223488 337408 223540 337414
rect 223488 337350 223540 337356
rect 222934 323096 222990 323105
rect 222934 323031 222990 323040
rect 222844 305652 222896 305658
rect 222844 305594 222896 305600
rect 222948 303686 222976 323031
rect 223592 308446 223620 373966
rect 226352 358834 226380 386990
rect 226444 361486 226472 390374
rect 227272 387054 227300 390374
rect 227260 387048 227312 387054
rect 227260 386990 227312 386996
rect 226432 361480 226484 361486
rect 226432 361422 226484 361428
rect 226444 360262 226472 361422
rect 226432 360256 226484 360262
rect 226432 360198 226484 360204
rect 226984 360256 227036 360262
rect 226984 360198 227036 360204
rect 226340 358828 226392 358834
rect 226340 358770 226392 358776
rect 226352 356726 226380 358770
rect 226340 356720 226392 356726
rect 226340 356662 226392 356668
rect 224224 342916 224276 342922
rect 224224 342858 224276 342864
rect 223670 325816 223726 325825
rect 223670 325751 223726 325760
rect 223580 308440 223632 308446
rect 223580 308382 223632 308388
rect 223212 304292 223264 304298
rect 223212 304234 223264 304240
rect 222936 303680 222988 303686
rect 222936 303622 222988 303628
rect 221016 301566 221398 301594
rect 221752 301566 222042 301594
rect 222304 301566 222594 301594
rect 223224 301580 223252 304234
rect 223684 301594 223712 325751
rect 224236 307057 224264 342858
rect 225142 328536 225198 328545
rect 225142 328471 225198 328480
rect 224222 307048 224278 307057
rect 224222 306983 224278 306992
rect 224408 303748 224460 303754
rect 224408 303690 224460 303696
rect 223684 301566 223882 301594
rect 224420 301580 224448 303690
rect 225050 302968 225106 302977
rect 225050 302903 225106 302912
rect 225064 301580 225092 302903
rect 225156 301594 225184 328471
rect 226996 320958 227024 360198
rect 227732 342922 227760 390374
rect 228362 388376 228418 388385
rect 228362 388311 228418 388320
rect 228376 356697 228404 388311
rect 229112 365022 229140 390374
rect 229100 365016 229152 365022
rect 229100 364958 229152 364964
rect 228362 356688 228418 356697
rect 228362 356623 228418 356632
rect 227720 342916 227772 342922
rect 227720 342858 227772 342864
rect 227718 336832 227774 336841
rect 227718 336767 227774 336776
rect 227076 326392 227128 326398
rect 227076 326334 227128 326340
rect 226984 320952 227036 320958
rect 226984 320894 227036 320900
rect 226982 316296 227038 316305
rect 226982 316231 227038 316240
rect 226340 314696 226392 314702
rect 226340 314638 226392 314644
rect 226352 307086 226380 314638
rect 226340 307080 226392 307086
rect 226340 307022 226392 307028
rect 226522 306640 226578 306649
rect 226522 306575 226578 306584
rect 226536 303822 226564 306575
rect 226996 304366 227024 316231
rect 227088 309777 227116 326334
rect 227732 325694 227760 336767
rect 227732 325666 228312 325694
rect 227074 309768 227130 309777
rect 227074 309703 227130 309712
rect 226984 304360 227036 304366
rect 226984 304302 227036 304308
rect 227442 304056 227498 304065
rect 227442 303991 227498 304000
rect 226524 303816 226576 303822
rect 226524 303758 226576 303764
rect 226248 303680 226300 303686
rect 226248 303622 226300 303628
rect 225156 301566 225630 301594
rect 226260 301580 226288 303622
rect 226798 302832 226854 302841
rect 226798 302767 226854 302776
rect 226812 301580 226840 302767
rect 227456 301580 227484 303991
rect 227718 301608 227774 301617
rect 228284 301594 228312 325666
rect 228376 315314 228404 356623
rect 229100 338224 229152 338230
rect 229100 338166 229152 338172
rect 228454 331392 228510 331401
rect 228454 331327 228510 331336
rect 228364 315308 228416 315314
rect 228364 315250 228416 315256
rect 228468 304201 228496 331327
rect 229112 325694 229140 338166
rect 229112 325666 229324 325694
rect 229296 306374 229324 325666
rect 229926 317656 229982 317665
rect 229926 317591 229982 317600
rect 229296 306346 229416 306374
rect 228454 304192 228510 304201
rect 228454 304127 228510 304136
rect 229190 303784 229246 303793
rect 229190 303719 229246 303728
rect 227774 301566 228022 301594
rect 228284 301566 228666 301594
rect 229204 301580 229232 303719
rect 229388 301594 229416 306346
rect 229940 301594 229968 317591
rect 230492 305697 230520 390374
rect 231228 386442 231256 390374
rect 231216 386436 231268 386442
rect 231216 386378 231268 386384
rect 231122 386336 231178 386345
rect 231122 386271 231178 386280
rect 231136 368490 231164 386271
rect 231228 380866 231256 386378
rect 231872 382294 231900 390374
rect 232504 385076 232556 385082
rect 232504 385018 232556 385024
rect 231860 382288 231912 382294
rect 231860 382230 231912 382236
rect 231216 380860 231268 380866
rect 231216 380802 231268 380808
rect 231872 378826 231900 382230
rect 231860 378820 231912 378826
rect 231860 378762 231912 378768
rect 232516 369170 232544 385018
rect 232504 369164 232556 369170
rect 232504 369106 232556 369112
rect 231124 368484 231176 368490
rect 231124 368426 231176 368432
rect 231136 359417 231164 368426
rect 232504 367872 232556 367878
rect 232504 367814 232556 367820
rect 231122 359408 231178 359417
rect 231122 359343 231178 359352
rect 231124 353320 231176 353326
rect 231124 353262 231176 353268
rect 230478 305688 230534 305697
rect 230478 305623 230534 305632
rect 231136 304298 231164 353262
rect 231214 342272 231270 342281
rect 231214 342207 231270 342216
rect 231124 304292 231176 304298
rect 231124 304234 231176 304240
rect 231032 303816 231084 303822
rect 231032 303758 231084 303764
rect 229388 301566 229862 301594
rect 229940 301566 230414 301594
rect 231044 301580 231072 303758
rect 231228 303657 231256 342207
rect 232516 333266 232544 367814
rect 232596 360868 232648 360874
rect 232596 360810 232648 360816
rect 232608 337482 232636 360810
rect 232596 337476 232648 337482
rect 232596 337418 232648 337424
rect 232504 333260 232556 333266
rect 232504 333202 232556 333208
rect 233148 332648 233200 332654
rect 233148 332590 233200 332596
rect 232504 329928 232556 329934
rect 232504 329870 232556 329876
rect 231860 311908 231912 311914
rect 231860 311850 231912 311856
rect 231584 305788 231636 305794
rect 231584 305730 231636 305736
rect 231214 303648 231270 303657
rect 231214 303583 231270 303592
rect 231596 301580 231624 305730
rect 231872 301594 231900 311850
rect 232516 301753 232544 329870
rect 232778 304192 232834 304201
rect 232778 304127 232834 304136
rect 232502 301744 232558 301753
rect 232502 301679 232558 301688
rect 231872 301566 232254 301594
rect 232792 301580 232820 304127
rect 233160 302938 233188 332590
rect 233252 307154 233280 390374
rect 234264 386345 234292 390388
rect 234632 390374 235382 390402
rect 236012 390374 236302 390402
rect 236656 390374 237222 390402
rect 234250 386336 234306 386345
rect 234250 386271 234306 386280
rect 234632 385665 234660 390374
rect 234618 385656 234674 385665
rect 234618 385591 234674 385600
rect 234632 380225 234660 385591
rect 234618 380216 234674 380225
rect 234618 380151 234674 380160
rect 236012 373998 236040 390374
rect 236656 385014 236684 390374
rect 238022 389872 238078 389881
rect 238022 389807 238078 389816
rect 236644 385008 236696 385014
rect 236644 384950 236696 384956
rect 236656 384334 236684 384950
rect 236644 384328 236696 384334
rect 236644 384270 236696 384276
rect 236000 373992 236052 373998
rect 236000 373934 236052 373940
rect 236012 372638 236040 373934
rect 236000 372632 236052 372638
rect 236000 372574 236052 372580
rect 236644 372632 236696 372638
rect 236644 372574 236696 372580
rect 233882 366344 233938 366353
rect 233882 366279 233938 366288
rect 233896 332654 233924 366279
rect 234804 346452 234856 346458
rect 234804 346394 234856 346400
rect 234712 345160 234764 345166
rect 234712 345102 234764 345108
rect 233976 342304 234028 342310
rect 233976 342246 234028 342252
rect 233884 332648 233936 332654
rect 233884 332590 233936 332596
rect 233988 319462 234016 342246
rect 233976 319456 234028 319462
rect 233976 319398 234028 319404
rect 233330 318880 233386 318889
rect 233330 318815 233386 318824
rect 233240 307148 233292 307154
rect 233240 307090 233292 307096
rect 233148 302932 233200 302938
rect 233148 302874 233200 302880
rect 233344 301594 233372 318815
rect 233974 308136 234030 308145
rect 233974 308071 234030 308080
rect 233344 301566 233450 301594
rect 233988 301580 234016 308071
rect 234618 303648 234674 303657
rect 234618 303583 234674 303592
rect 234632 301580 234660 303583
rect 234724 301594 234752 345102
rect 234816 325694 234844 346394
rect 236656 326398 236684 372574
rect 238036 348430 238064 389807
rect 238128 388385 238156 390388
rect 238760 389224 238812 389230
rect 238760 389166 238812 389172
rect 238114 388376 238170 388385
rect 238114 388311 238170 388320
rect 238666 366480 238722 366489
rect 238666 366415 238722 366424
rect 238024 348424 238076 348430
rect 238024 348366 238076 348372
rect 236644 326392 236696 326398
rect 236644 326334 236696 326340
rect 234816 325666 235488 325694
rect 235460 301594 235488 325666
rect 236552 313948 236604 313954
rect 236552 313890 236604 313896
rect 236368 304360 236420 304366
rect 236368 304302 236420 304308
rect 234724 301566 235198 301594
rect 235460 301566 235842 301594
rect 236380 301580 236408 304302
rect 236564 301594 236592 313890
rect 238680 313342 238708 366415
rect 238772 338162 238800 389166
rect 239048 385082 239076 390388
rect 239968 389230 239996 390388
rect 240152 390374 241086 390402
rect 242006 390374 242296 390402
rect 239956 389224 240008 389230
rect 239956 389166 240008 389172
rect 239036 385076 239088 385082
rect 239036 385018 239088 385024
rect 240046 361720 240102 361729
rect 240046 361655 240102 361664
rect 238760 338156 238812 338162
rect 238760 338098 238812 338104
rect 239404 338156 239456 338162
rect 239404 338098 239456 338104
rect 239416 324970 239444 338098
rect 239404 324964 239456 324970
rect 239404 324906 239456 324912
rect 239402 320376 239458 320385
rect 239402 320311 239458 320320
rect 239416 313954 239444 320311
rect 239404 313948 239456 313954
rect 239404 313890 239456 313896
rect 238668 313336 238720 313342
rect 238720 313284 238800 313290
rect 238668 313278 238800 313284
rect 238680 313262 238800 313278
rect 238680 313213 238708 313262
rect 237378 309224 237434 309233
rect 237378 309159 237434 309168
rect 237392 301594 237420 309159
rect 238206 306912 238262 306921
rect 238206 306847 238262 306856
rect 236564 301566 237038 301594
rect 237392 301566 237590 301594
rect 238220 301580 238248 306847
rect 238772 306374 238800 313262
rect 238772 306346 238984 306374
rect 238850 303920 238906 303929
rect 238850 303855 238906 303864
rect 238864 301580 238892 303855
rect 238956 301594 238984 306346
rect 240060 305046 240088 361655
rect 240152 357406 240180 390374
rect 242268 389065 242296 390374
rect 242254 389056 242310 389065
rect 242254 388991 242310 389000
rect 240784 386300 240836 386306
rect 240784 386242 240836 386248
rect 240232 369232 240284 369238
rect 240232 369174 240284 369180
rect 240140 357400 240192 357406
rect 240140 357342 240192 357348
rect 240244 329866 240272 369174
rect 240796 365702 240824 386242
rect 242162 371920 242218 371929
rect 242162 371855 242218 371864
rect 240784 365696 240836 365702
rect 240784 365638 240836 365644
rect 240784 357400 240836 357406
rect 240784 357342 240836 357348
rect 240232 329860 240284 329866
rect 240232 329802 240284 329808
rect 240244 325694 240272 329802
rect 240796 325694 240824 357342
rect 240244 325666 240732 325694
rect 240796 325666 240916 325694
rect 240704 306374 240732 325666
rect 240704 306346 240824 306374
rect 240048 305040 240100 305046
rect 240048 304982 240100 304988
rect 240598 305008 240654 305017
rect 238956 301566 239430 301594
rect 240060 301580 240088 304982
rect 240598 304943 240654 304952
rect 240612 301580 240640 304943
rect 240796 301594 240824 306346
rect 240888 301714 240916 325666
rect 242176 302297 242204 371855
rect 242268 361593 242296 388991
rect 242912 385665 242940 390388
rect 243096 390374 243846 390402
rect 244292 390374 244766 390402
rect 245686 390374 245792 390402
rect 242898 385656 242954 385665
rect 242898 385591 242954 385600
rect 243096 379506 243124 390374
rect 243084 379500 243136 379506
rect 243084 379442 243136 379448
rect 243096 379030 243124 379442
rect 243084 379024 243136 379030
rect 243084 378966 243136 378972
rect 243544 379024 243596 379030
rect 243544 378966 243596 378972
rect 243556 370569 243584 378966
rect 242990 370560 243046 370569
rect 242990 370495 243046 370504
rect 243542 370560 243598 370569
rect 243542 370495 243598 370504
rect 242254 361584 242310 361593
rect 242254 361519 242310 361528
rect 242900 359508 242952 359514
rect 242900 359450 242952 359456
rect 242912 331362 242940 359450
rect 242900 331356 242952 331362
rect 242900 331298 242952 331304
rect 242808 328092 242860 328098
rect 242808 328034 242860 328040
rect 242820 308417 242848 328034
rect 242806 308408 242862 308417
rect 242806 308343 242862 308352
rect 242438 303784 242494 303793
rect 242438 303719 242494 303728
rect 241794 302288 241850 302297
rect 241794 302223 241850 302232
rect 242162 302288 242218 302297
rect 242162 302223 242218 302232
rect 240876 301708 240928 301714
rect 240876 301650 240928 301656
rect 240796 301566 241270 301594
rect 241808 301580 241836 302223
rect 242452 301580 242480 303719
rect 242912 301594 242940 331298
rect 243004 325718 243032 370495
rect 244292 340202 244320 390374
rect 245764 375358 245792 390374
rect 246592 389162 246620 390388
rect 247604 390374 247710 390402
rect 248340 390374 248630 390402
rect 246396 389156 246448 389162
rect 246396 389098 246448 389104
rect 246580 389156 246632 389162
rect 246580 389098 246632 389104
rect 245752 375352 245804 375358
rect 245752 375294 245804 375300
rect 245764 374610 245792 375294
rect 245752 374604 245804 374610
rect 245752 374546 245804 374552
rect 246304 374604 246356 374610
rect 246304 374546 246356 374552
rect 244922 371376 244978 371385
rect 244922 371311 244978 371320
rect 244372 341556 244424 341562
rect 244372 341498 244424 341504
rect 244384 340950 244412 341498
rect 244372 340944 244424 340950
rect 244372 340886 244424 340892
rect 244280 340196 244332 340202
rect 244280 340138 244332 340144
rect 244384 328098 244412 340886
rect 244372 328092 244424 328098
rect 244372 328034 244424 328040
rect 242992 325712 243044 325718
rect 243044 325666 243216 325694
rect 242992 325654 243044 325660
rect 243082 313984 243138 313993
rect 243082 313919 243138 313928
rect 243096 303686 243124 313919
rect 243084 303680 243136 303686
rect 243084 303622 243136 303628
rect 243188 301594 243216 325666
rect 244936 309233 244964 371311
rect 245660 331288 245712 331294
rect 245660 331230 245712 331236
rect 245672 325694 245700 331230
rect 245672 325666 246160 325694
rect 244922 309224 244978 309233
rect 244922 309159 244978 309168
rect 243820 303680 243872 303686
rect 243820 303622 243872 303628
rect 243832 301594 243860 303622
rect 244936 301594 244964 309159
rect 246028 305652 246080 305658
rect 246028 305594 246080 305600
rect 242912 301566 243018 301594
rect 243188 301566 243662 301594
rect 243832 301566 244214 301594
rect 244858 301566 244964 301594
rect 246040 301580 246068 305594
rect 246132 301594 246160 325666
rect 246316 302841 246344 374546
rect 246408 330546 246436 389098
rect 247604 388929 247632 390374
rect 247684 389836 247736 389842
rect 247684 389778 247736 389784
rect 247038 388920 247094 388929
rect 247038 388855 247094 388864
rect 247590 388920 247646 388929
rect 247590 388855 247646 388864
rect 247052 386306 247080 388855
rect 247040 386300 247092 386306
rect 247040 386242 247092 386248
rect 247696 376718 247724 389778
rect 248340 389298 248368 390374
rect 248328 389292 248380 389298
rect 248328 389234 248380 389240
rect 249156 389224 249208 389230
rect 249156 389166 249208 389172
rect 249062 384976 249118 384985
rect 249062 384911 249118 384920
rect 247040 376712 247092 376718
rect 247040 376654 247092 376660
rect 247684 376712 247736 376718
rect 247684 376654 247736 376660
rect 247052 334014 247080 376654
rect 247040 334008 247092 334014
rect 247040 333950 247092 333956
rect 247684 334008 247736 334014
rect 247684 333950 247736 333956
rect 246396 330540 246448 330546
rect 246396 330482 246448 330488
rect 246394 327720 246450 327729
rect 246394 327655 246450 327664
rect 246302 302832 246358 302841
rect 246302 302767 246358 302776
rect 246408 301753 246436 327655
rect 246488 318844 246540 318850
rect 246488 318786 246540 318792
rect 246500 312594 246528 318786
rect 246488 312588 246540 312594
rect 246488 312530 246540 312536
rect 247696 302258 247724 333950
rect 249076 311273 249104 384911
rect 249168 349926 249196 389166
rect 249248 387864 249300 387870
rect 249248 387806 249300 387812
rect 249260 353258 249288 387806
rect 249536 384985 249564 390388
rect 249812 390374 250470 390402
rect 249522 384976 249578 384985
rect 249522 384911 249578 384920
rect 249708 353320 249760 353326
rect 249708 353262 249760 353268
rect 249248 353252 249300 353258
rect 249248 353194 249300 353200
rect 249156 349920 249208 349926
rect 249156 349862 249208 349868
rect 249062 311264 249118 311273
rect 249062 311199 249118 311208
rect 249616 311160 249668 311166
rect 249616 311102 249668 311108
rect 249628 306513 249656 311102
rect 249614 306504 249670 306513
rect 249614 306439 249670 306448
rect 249248 305108 249300 305114
rect 249248 305050 249300 305056
rect 248970 304600 249026 304609
rect 248970 304535 249026 304544
rect 248984 303686 249012 304535
rect 248420 303680 248472 303686
rect 247866 303648 247922 303657
rect 248420 303622 248472 303628
rect 248972 303680 249024 303686
rect 248972 303622 249024 303628
rect 247866 303583 247922 303592
rect 247684 302252 247736 302258
rect 247684 302194 247736 302200
rect 246394 301744 246450 301753
rect 246394 301679 246450 301688
rect 247222 301744 247278 301753
rect 247222 301679 247278 301688
rect 246132 301566 246606 301594
rect 247236 301580 247264 301679
rect 247696 301594 247724 302194
rect 247880 301753 247908 303583
rect 247866 301744 247922 301753
rect 247866 301679 247922 301688
rect 247696 301566 247802 301594
rect 248432 301580 248460 303622
rect 249260 301594 249288 305050
rect 248998 301566 249288 301594
rect 249628 301580 249656 306439
rect 249720 305114 249748 353262
rect 249812 351898 249840 390374
rect 251376 387870 251404 390388
rect 251836 390374 252310 390402
rect 251836 389094 251864 390374
rect 251824 389088 251876 389094
rect 251824 389030 251876 389036
rect 251364 387864 251416 387870
rect 251364 387806 251416 387812
rect 251836 382974 251864 389030
rect 251824 382968 251876 382974
rect 251824 382910 251876 382916
rect 251824 382220 251876 382226
rect 251824 382162 251876 382168
rect 249800 351892 249852 351898
rect 249800 351834 249852 351840
rect 251836 335374 251864 382162
rect 252468 370524 252520 370530
rect 252468 370466 252520 370472
rect 251824 335368 251876 335374
rect 251824 335310 251876 335316
rect 249800 324964 249852 324970
rect 249800 324906 249852 324912
rect 249708 305108 249760 305114
rect 249708 305050 249760 305056
rect 249812 301594 249840 324906
rect 250810 307864 250866 307873
rect 251836 307834 251864 335310
rect 250810 307799 250866 307808
rect 251824 307828 251876 307834
rect 249812 301566 250194 301594
rect 250824 301580 250852 307799
rect 251824 307770 251876 307776
rect 251362 303648 251418 303657
rect 251362 303583 251418 303592
rect 251376 301580 251404 303583
rect 251836 301594 251864 307770
rect 252480 302190 252508 370466
rect 252572 362914 252600 390895
rect 252664 390374 253414 390402
rect 252664 372570 252692 390374
rect 253492 387122 253520 393286
rect 253480 387116 253532 387122
rect 253480 387058 253532 387064
rect 252744 383648 252796 383654
rect 252744 383590 252796 383596
rect 252756 382294 252784 383590
rect 252744 382288 252796 382294
rect 252744 382230 252796 382236
rect 252652 372564 252704 372570
rect 252652 372506 252704 372512
rect 253848 363792 253900 363798
rect 253848 363734 253900 363740
rect 252560 362908 252612 362914
rect 252560 362850 252612 362856
rect 252572 353326 252600 362850
rect 252560 353320 252612 353326
rect 252560 353262 252612 353268
rect 253204 342916 253256 342922
rect 253204 342858 253256 342864
rect 252560 307148 252612 307154
rect 252560 307090 252612 307096
rect 252468 302184 252520 302190
rect 252468 302126 252520 302132
rect 251836 301566 252034 301594
rect 227718 301543 227774 301552
rect 245108 301096 245160 301102
rect 242070 301064 242126 301073
rect 245160 301044 245410 301050
rect 245108 301038 245410 301044
rect 245120 301022 245410 301038
rect 242070 300999 242072 301008
rect 242124 300999 242126 301008
rect 242072 300970 242124 300976
rect 199476 300960 199528 300966
rect 194690 300928 194746 300937
rect 194746 300886 195086 300914
rect 214564 300960 214616 300966
rect 209134 300928 209190 300937
rect 199528 300908 199870 300914
rect 199476 300902 199870 300908
rect 199488 300886 199870 300902
rect 194690 300863 194746 300872
rect 209190 300886 209438 300914
rect 214564 300902 214616 300908
rect 209134 300863 209190 300872
rect 252468 300824 252520 300830
rect 252466 300792 252468 300801
rect 252520 300792 252522 300801
rect 252466 300727 252522 300736
rect 193494 299024 193550 299033
rect 193494 298959 193550 298968
rect 193404 295384 193456 295390
rect 193404 295326 193456 295332
rect 192574 285696 192630 285705
rect 192574 285631 192630 285640
rect 193126 285696 193182 285705
rect 193126 285631 193182 285640
rect 192588 243574 192616 285631
rect 192668 256216 192720 256222
rect 192668 256158 192720 256164
rect 192576 243568 192628 243574
rect 192576 243510 192628 243516
rect 192116 242956 192168 242962
rect 192116 242898 192168 242904
rect 192484 242956 192536 242962
rect 192484 242898 192536 242904
rect 192128 241466 192156 242898
rect 192116 241460 192168 241466
rect 192116 241402 192168 241408
rect 192588 236609 192616 243510
rect 192680 240038 192708 256158
rect 193220 251864 193272 251870
rect 193220 251806 193272 251812
rect 192668 240032 192720 240038
rect 192668 239974 192720 239980
rect 193126 239864 193182 239873
rect 193126 239799 193182 239808
rect 192574 236600 192630 236609
rect 192574 236535 192630 236544
rect 193140 199442 193168 239799
rect 193128 199436 193180 199442
rect 193128 199378 193180 199384
rect 193232 166297 193260 251806
rect 193588 246356 193640 246362
rect 193588 246298 193640 246304
rect 193600 238754 193628 246298
rect 193678 242856 193734 242865
rect 193678 242791 193734 242800
rect 193692 242026 193720 242791
rect 252376 242344 252428 242350
rect 252376 242286 252428 242292
rect 195336 242072 195388 242078
rect 193770 242040 193826 242049
rect 193692 241998 193770 242026
rect 193770 241975 193826 241984
rect 194506 242040 194562 242049
rect 195796 242072 195848 242078
rect 195336 242014 195388 242020
rect 195794 242040 195796 242049
rect 248512 242072 248564 242078
rect 195848 242040 195850 242049
rect 194506 241975 194562 241984
rect 193600 238726 193812 238754
rect 193784 237318 193812 238726
rect 193772 237312 193824 237318
rect 193772 237254 193824 237260
rect 194520 188358 194548 241975
rect 194810 241590 195284 241618
rect 195256 239737 195284 241590
rect 195242 239728 195298 239737
rect 195242 239663 195298 239672
rect 195256 196654 195284 239663
rect 195348 227050 195376 242014
rect 195794 241975 195850 241984
rect 248510 242040 248512 242049
rect 250444 242072 250496 242078
rect 248564 242040 248566 242049
rect 250444 242014 250496 242020
rect 248510 241975 248566 241984
rect 196164 240032 196216 240038
rect 196164 239974 196216 239980
rect 196176 239426 196204 239974
rect 196164 239420 196216 239426
rect 196164 239362 196216 239368
rect 195336 227044 195388 227050
rect 195336 226986 195388 226992
rect 195244 196648 195296 196654
rect 195244 196590 195296 196596
rect 195244 193860 195296 193866
rect 195244 193802 195296 193808
rect 194508 188352 194560 188358
rect 194508 188294 194560 188300
rect 193496 184204 193548 184210
rect 193496 184146 193548 184152
rect 193218 166288 193274 166297
rect 193218 166223 193274 166232
rect 191930 164384 191986 164393
rect 191930 164319 191986 164328
rect 191944 161430 191972 164319
rect 191932 161424 191984 161430
rect 191932 161366 191984 161372
rect 191944 160138 191972 161366
rect 191932 160132 191984 160138
rect 191932 160074 191984 160080
rect 193128 158772 193180 158778
rect 193128 158714 193180 158720
rect 193140 154562 193168 158714
rect 193128 154556 193180 154562
rect 193128 154498 193180 154504
rect 191840 148368 191892 148374
rect 191840 148310 191892 148316
rect 192484 147076 192536 147082
rect 192484 147018 192536 147024
rect 191654 139904 191710 139913
rect 191654 139839 191710 139848
rect 191654 137456 191710 137465
rect 191654 137391 191710 137400
rect 191668 136678 191696 137391
rect 191656 136672 191708 136678
rect 191656 136614 191708 136620
rect 191748 136604 191800 136610
rect 191748 136546 191800 136552
rect 191760 136377 191788 136546
rect 191746 136368 191802 136377
rect 191746 136303 191802 136312
rect 191746 135552 191802 135561
rect 191746 135487 191802 135496
rect 191760 135318 191788 135487
rect 191748 135312 191800 135318
rect 191748 135254 191800 135260
rect 192496 135250 192524 147018
rect 192576 145580 192628 145586
rect 192576 145522 192628 145528
rect 192484 135244 192536 135250
rect 192484 135186 192536 135192
rect 191748 133884 191800 133890
rect 191748 133826 191800 133832
rect 191760 132841 191788 133826
rect 191746 132832 191802 132841
rect 191746 132767 191802 132776
rect 191748 128308 191800 128314
rect 191748 128250 191800 128256
rect 191760 127673 191788 128250
rect 191746 127664 191802 127673
rect 191746 127599 191802 127608
rect 191562 126576 191618 126585
rect 191562 126511 191618 126520
rect 191656 126268 191708 126274
rect 191656 126210 191708 126216
rect 191470 123856 191526 123865
rect 191470 123791 191526 123800
rect 191010 123040 191066 123049
rect 191010 122975 191066 122984
rect 190550 118688 190606 118697
rect 190550 118623 190606 118632
rect 191010 118688 191066 118697
rect 191010 118623 191066 118632
rect 191024 117978 191052 118623
rect 191012 117972 191064 117978
rect 191012 117914 191064 117920
rect 191668 117609 191696 126210
rect 191746 122224 191802 122233
rect 191746 122159 191802 122168
rect 191760 122126 191788 122159
rect 191748 122120 191800 122126
rect 191748 122062 191800 122068
rect 191748 121440 191800 121446
rect 191746 121408 191748 121417
rect 191800 121408 191802 121417
rect 191746 121343 191802 121352
rect 191746 120320 191802 120329
rect 191746 120255 191802 120264
rect 191760 120222 191788 120255
rect 191748 120216 191800 120222
rect 191748 120158 191800 120164
rect 191748 120080 191800 120086
rect 191748 120022 191800 120028
rect 191760 119513 191788 120022
rect 191746 119504 191802 119513
rect 191746 119439 191802 119448
rect 191654 117600 191710 117609
rect 191654 117535 191710 117544
rect 191012 117224 191064 117230
rect 191012 117166 191064 117172
rect 191024 115977 191052 117166
rect 191010 115968 191066 115977
rect 190828 115932 190880 115938
rect 191010 115903 191066 115912
rect 190828 115874 190880 115880
rect 190840 115161 190868 115874
rect 190826 115152 190882 115161
rect 190826 115087 190882 115096
rect 191102 109712 191158 109721
rect 191102 109647 191158 109656
rect 191116 100094 191144 109647
rect 191196 106276 191248 106282
rect 191196 106218 191248 106224
rect 191208 106185 191236 106218
rect 191194 106176 191250 106185
rect 191194 106111 191250 106120
rect 191472 101448 191524 101454
rect 191472 101390 191524 101396
rect 191104 100088 191156 100094
rect 191104 100030 191156 100036
rect 190552 98048 190604 98054
rect 190550 98016 190552 98025
rect 190604 98016 190606 98025
rect 190460 97980 190512 97986
rect 190550 97951 190606 97960
rect 190460 97922 190512 97928
rect 190472 97209 190500 97922
rect 190458 97200 190514 97209
rect 190458 97135 190514 97144
rect 191378 95432 191434 95441
rect 191378 95367 191434 95376
rect 190458 93664 190514 93673
rect 190458 93599 190514 93608
rect 190472 93226 190500 93599
rect 190460 93220 190512 93226
rect 190460 93162 190512 93168
rect 190366 85504 190422 85513
rect 190366 85439 190422 85448
rect 191392 84833 191420 95367
rect 191484 94586 191512 101390
rect 191562 100736 191618 100745
rect 191562 100671 191618 100680
rect 191472 94580 191524 94586
rect 191472 94522 191524 94528
rect 191378 84824 191434 84833
rect 191378 84759 191434 84768
rect 191576 78674 191604 100671
rect 191564 78668 191616 78674
rect 191564 78610 191616 78616
rect 190276 44872 190328 44878
rect 190276 44814 190328 44820
rect 191668 43450 191696 117535
rect 191748 117292 191800 117298
rect 191748 117234 191800 117240
rect 191760 116793 191788 117234
rect 191746 116784 191802 116793
rect 191746 116719 191802 116728
rect 191838 114064 191894 114073
rect 191838 113999 191894 114008
rect 191746 113248 191802 113257
rect 191746 113183 191748 113192
rect 191800 113183 191802 113192
rect 191748 113154 191800 113160
rect 191748 112464 191800 112470
rect 191746 112432 191748 112441
rect 191800 112432 191802 112441
rect 191746 112367 191802 112376
rect 191852 110566 191880 113999
rect 191840 110560 191892 110566
rect 191746 110528 191802 110537
rect 191840 110502 191892 110508
rect 191746 110463 191748 110472
rect 191800 110463 191802 110472
rect 191748 110434 191800 110440
rect 192022 108352 192078 108361
rect 192022 108287 192078 108296
rect 192036 107681 192064 108287
rect 192022 107672 192078 107681
rect 191748 107636 191800 107642
rect 192022 107607 192078 107616
rect 191748 107578 191800 107584
rect 191760 107001 191788 107578
rect 191746 106992 191802 107001
rect 191746 106927 191802 106936
rect 191748 105596 191800 105602
rect 191748 105538 191800 105544
rect 191760 105097 191788 105538
rect 191746 105088 191802 105097
rect 191746 105023 191802 105032
rect 192496 104281 192524 135186
rect 192588 129062 192616 145522
rect 193036 140480 193088 140486
rect 193036 140422 193088 140428
rect 193048 138281 193076 140422
rect 193034 138272 193090 138281
rect 193034 138207 193090 138216
rect 192942 132016 192998 132025
rect 192942 131951 192998 131960
rect 192956 131510 192984 131951
rect 192944 131504 192996 131510
rect 192944 131446 192996 131452
rect 192576 129056 192628 129062
rect 192576 128998 192628 129004
rect 192482 104272 192538 104281
rect 192482 104207 192538 104216
rect 191746 103456 191802 103465
rect 191746 103391 191802 103400
rect 191760 102270 191788 103391
rect 191748 102264 191800 102270
rect 191748 102206 191800 102212
rect 191746 101552 191802 101561
rect 191746 101487 191802 101496
rect 191760 101454 191788 101487
rect 191748 101448 191800 101454
rect 191748 101390 191800 101396
rect 191748 100700 191800 100706
rect 191748 100642 191800 100648
rect 191760 99929 191788 100642
rect 191746 99920 191802 99929
rect 191746 99855 191802 99864
rect 191748 94580 191800 94586
rect 191748 94522 191800 94528
rect 191656 43444 191708 43450
rect 191656 43386 191708 43392
rect 185676 19984 185728 19990
rect 185676 19926 185728 19932
rect 173164 9036 173216 9042
rect 173164 8978 173216 8984
rect 191760 7614 191788 94522
rect 191840 94512 191892 94518
rect 191840 94454 191892 94460
rect 191852 93430 191880 94454
rect 192850 93800 192906 93809
rect 192850 93735 192906 93744
rect 191840 93424 191892 93430
rect 191840 93366 191892 93372
rect 192864 68338 192892 93735
rect 192956 86193 192984 131446
rect 193140 124953 193168 154498
rect 193312 140820 193364 140826
rect 193312 140762 193364 140768
rect 193324 140049 193352 140762
rect 193310 140040 193366 140049
rect 193310 139975 193366 139984
rect 193404 138712 193456 138718
rect 193402 138680 193404 138689
rect 193456 138680 193458 138689
rect 193402 138615 193458 138624
rect 193508 132494 193536 184146
rect 194784 172508 194836 172514
rect 194784 172450 194836 172456
rect 194796 171834 194824 172450
rect 194784 171828 194836 171834
rect 194784 171770 194836 171776
rect 194690 147928 194746 147937
rect 194690 147863 194746 147872
rect 193586 144256 193642 144265
rect 193586 144191 193642 144200
rect 193600 140964 193628 144191
rect 194140 143676 194192 143682
rect 194140 143618 194192 143624
rect 194152 140964 194180 143618
rect 194704 143449 194732 147863
rect 194690 143440 194746 143449
rect 194690 143375 194746 143384
rect 194704 140964 194732 143375
rect 194796 140486 194824 171770
rect 195256 141137 195284 193802
rect 195336 192500 195388 192506
rect 195336 192442 195388 192448
rect 195348 172514 195376 192442
rect 195336 172508 195388 172514
rect 195336 172450 195388 172456
rect 195980 168428 196032 168434
rect 195980 168370 196032 168376
rect 195886 152008 195942 152017
rect 195886 151943 195942 151952
rect 195900 142154 195928 151943
rect 195808 142126 195928 142154
rect 195242 141128 195298 141137
rect 195242 141063 195298 141072
rect 195808 140978 195836 142126
rect 195454 140950 195836 140978
rect 195992 140964 196020 168370
rect 196070 152144 196126 152153
rect 196070 152079 196126 152088
rect 196084 140978 196112 152079
rect 196176 143449 196204 239362
rect 197188 235278 197216 241604
rect 199594 241590 200068 241618
rect 197358 237960 197414 237969
rect 197358 237895 197414 237904
rect 197176 235272 197228 235278
rect 197176 235214 197228 235220
rect 196624 232552 196676 232558
rect 196624 232494 196676 232500
rect 196636 223582 196664 232494
rect 196624 223576 196676 223582
rect 196624 223518 196676 223524
rect 196624 213988 196676 213994
rect 196624 213930 196676 213936
rect 196636 206990 196664 213930
rect 196624 206984 196676 206990
rect 196624 206926 196676 206932
rect 197268 206984 197320 206990
rect 197268 206926 197320 206932
rect 196624 198008 196676 198014
rect 196624 197950 196676 197956
rect 196636 168434 196664 197950
rect 197280 175953 197308 206926
rect 197266 175944 197322 175953
rect 197266 175879 197322 175888
rect 196624 168428 196676 168434
rect 196624 168370 196676 168376
rect 196622 143576 196678 143585
rect 196622 143511 196678 143520
rect 196162 143440 196218 143449
rect 196162 143375 196218 143384
rect 196084 140950 196558 140978
rect 196636 140826 196664 143511
rect 197372 140978 197400 237895
rect 200040 203590 200068 241590
rect 201972 241534 202000 241604
rect 201500 241528 201552 241534
rect 201500 241470 201552 241476
rect 201960 241528 202012 241534
rect 201960 241470 202012 241476
rect 201406 205728 201462 205737
rect 201406 205663 201462 205672
rect 200028 203584 200080 203590
rect 200028 203526 200080 203532
rect 201420 202774 201448 205663
rect 201408 202768 201460 202774
rect 201408 202710 201460 202716
rect 198096 181484 198148 181490
rect 198096 181426 198148 181432
rect 198002 167648 198058 167657
rect 198002 167583 198058 167592
rect 198016 149841 198044 167583
rect 198108 166394 198136 181426
rect 201420 167657 201448 202710
rect 201512 181558 201540 241470
rect 204364 241466 204392 241604
rect 204352 241460 204404 241466
rect 204352 241402 204404 241408
rect 206756 239426 206784 241604
rect 206744 239420 206796 239426
rect 206744 239362 206796 239368
rect 209148 238678 209176 241604
rect 211554 241590 211844 241618
rect 211816 240106 211844 241590
rect 211804 240100 211856 240106
rect 211804 240042 211856 240048
rect 209136 238672 209188 238678
rect 209136 238614 209188 238620
rect 202878 233880 202934 233889
rect 202878 233815 202934 233824
rect 202234 214568 202290 214577
rect 202234 214503 202290 214512
rect 202248 202842 202276 214503
rect 201592 202836 201644 202842
rect 201592 202778 201644 202784
rect 202236 202836 202288 202842
rect 202236 202778 202288 202784
rect 201500 181552 201552 181558
rect 201500 181494 201552 181500
rect 201500 172576 201552 172582
rect 201500 172518 201552 172524
rect 201512 171086 201540 172518
rect 201500 171080 201552 171086
rect 201500 171022 201552 171028
rect 201406 167648 201462 167657
rect 201406 167583 201462 167592
rect 198096 166388 198148 166394
rect 198096 166330 198148 166336
rect 200120 163940 200172 163946
rect 200120 163882 200172 163888
rect 199292 151088 199344 151094
rect 199292 151030 199344 151036
rect 198002 149832 198058 149841
rect 198002 149767 198058 149776
rect 199304 149190 199332 151030
rect 199292 149184 199344 149190
rect 199292 149126 199344 149132
rect 198830 148472 198886 148481
rect 198830 148407 198886 148416
rect 197912 147008 197964 147014
rect 197912 146950 197964 146956
rect 197924 140978 197952 146950
rect 198844 140978 198872 148407
rect 199304 140978 199332 149126
rect 200132 140978 200160 163882
rect 201512 151814 201540 171022
rect 201604 155281 201632 202778
rect 201590 155272 201646 155281
rect 201590 155207 201646 155216
rect 201512 151786 202276 151814
rect 201408 149728 201460 149734
rect 201408 149670 201460 149676
rect 201420 147801 201448 149670
rect 200302 147792 200358 147801
rect 200302 147727 200358 147736
rect 201406 147792 201462 147801
rect 201406 147727 201462 147736
rect 200316 140978 200344 147727
rect 201590 145616 201646 145625
rect 201590 145551 201646 145560
rect 201314 144120 201370 144129
rect 201314 144055 201370 144064
rect 197372 140950 197846 140978
rect 197924 140950 198398 140978
rect 198844 140950 198950 140978
rect 199304 140950 199686 140978
rect 200132 140950 200238 140978
rect 200316 140950 200790 140978
rect 201328 140964 201356 144055
rect 201604 140978 201632 145551
rect 202248 140978 202276 151786
rect 202892 141001 202920 233815
rect 204904 232552 204956 232558
rect 204904 232494 204956 232500
rect 204444 229764 204496 229770
rect 204444 229706 204496 229712
rect 204456 223514 204484 229706
rect 204444 223508 204496 223514
rect 204444 223450 204496 223456
rect 204916 177342 204944 232494
rect 206282 222864 206338 222873
rect 206282 222799 206338 222808
rect 204996 221468 205048 221474
rect 204996 221410 205048 221416
rect 205008 209001 205036 221410
rect 204994 208992 205050 209001
rect 204994 208927 205050 208936
rect 204996 195288 205048 195294
rect 204996 195230 205048 195236
rect 204904 177336 204956 177342
rect 204904 177278 204956 177284
rect 203524 174548 203576 174554
rect 203524 174490 203576 174496
rect 203536 170406 203564 174490
rect 202972 170400 203024 170406
rect 202972 170342 203024 170348
rect 203524 170400 203576 170406
rect 203524 170342 203576 170348
rect 202984 151814 203012 170342
rect 204916 151814 204944 177278
rect 205008 163946 205036 195230
rect 206296 180130 206324 222799
rect 210422 217288 210478 217297
rect 210422 217223 210478 217232
rect 209042 202328 209098 202337
rect 209042 202263 209098 202272
rect 206284 180124 206336 180130
rect 206284 180066 206336 180072
rect 205638 174584 205694 174593
rect 205638 174519 205694 174528
rect 204996 163940 205048 163946
rect 204996 163882 205048 163888
rect 204994 153776 205050 153785
rect 204994 153711 205050 153720
rect 202984 151786 203472 151814
rect 202878 140992 202934 141001
rect 201604 140950 202078 140978
rect 202248 140950 202630 140978
rect 203444 140978 203472 151786
rect 204548 151786 204944 151814
rect 204548 149122 204576 151786
rect 204536 149116 204588 149122
rect 204536 149058 204588 149064
rect 204350 147656 204406 147665
rect 204350 147591 204406 147600
rect 204364 140978 204392 147591
rect 204548 140978 204576 149058
rect 205008 143682 205036 153711
rect 204996 143676 205048 143682
rect 204996 143618 205048 143624
rect 205454 140992 205510 141001
rect 203444 140950 203918 140978
rect 204364 140950 204470 140978
rect 204548 140950 205022 140978
rect 202878 140927 202934 140936
rect 205454 140927 205510 140936
rect 202892 140842 202920 140927
rect 202892 140826 203472 140842
rect 196624 140820 196676 140826
rect 202892 140820 203484 140826
rect 202892 140814 203432 140820
rect 196624 140762 196676 140768
rect 203432 140762 203484 140768
rect 205468 140570 205496 140927
rect 205192 140554 205574 140570
rect 205180 140548 205574 140554
rect 205232 140542 205574 140548
rect 205180 140490 205232 140496
rect 194784 140480 194836 140486
rect 194784 140422 194836 140428
rect 196806 140448 196862 140457
rect 205652 140434 205680 174519
rect 209056 167793 209084 202263
rect 209964 177336 210016 177342
rect 209964 177278 210016 177284
rect 209042 167784 209098 167793
rect 209042 167719 209098 167728
rect 207664 166320 207716 166326
rect 207664 166262 207716 166268
rect 207020 152584 207072 152590
rect 207020 152526 207072 152532
rect 207032 151814 207060 152526
rect 207032 151786 207428 151814
rect 207110 149832 207166 149841
rect 207110 149767 207166 149776
rect 206928 147756 206980 147762
rect 206928 147698 206980 147704
rect 206558 140584 206614 140593
rect 206940 140570 206968 147698
rect 207124 140978 207152 149767
rect 207400 142154 207428 151786
rect 207676 147626 207704 166262
rect 208584 159384 208636 159390
rect 208584 159326 208636 159332
rect 208596 157457 208624 159326
rect 208398 157448 208454 157457
rect 208398 157383 208454 157392
rect 208582 157448 208638 157457
rect 208582 157383 208638 157392
rect 207664 147620 207716 147626
rect 207664 147562 207716 147568
rect 208412 147014 208440 157383
rect 209872 156460 209924 156466
rect 209872 156402 209924 156408
rect 208490 153776 208546 153785
rect 208490 153711 208546 153720
rect 208504 151881 208532 153711
rect 208490 151872 208546 151881
rect 208490 151807 208546 151816
rect 208400 147008 208452 147014
rect 208400 146950 208452 146956
rect 207400 142126 207796 142154
rect 207768 140978 207796 142126
rect 208504 140978 208532 151807
rect 209884 147014 209912 156402
rect 209976 151814 210004 177278
rect 210436 169153 210464 217223
rect 211816 189145 211844 240042
rect 213932 235958 213960 241604
rect 215300 238060 215352 238066
rect 215300 238002 215352 238008
rect 213920 235952 213972 235958
rect 213920 235894 213972 235900
rect 213932 234666 213960 235894
rect 213920 234660 213972 234666
rect 213920 234602 213972 234608
rect 214656 234660 214708 234666
rect 214656 234602 214708 234608
rect 213828 231124 213880 231130
rect 213828 231066 213880 231072
rect 213840 227633 213868 231066
rect 213826 227624 213882 227633
rect 213826 227559 213882 227568
rect 213184 189780 213236 189786
rect 213184 189722 213236 189728
rect 211802 189136 211858 189145
rect 211802 189071 211858 189080
rect 211802 186960 211858 186969
rect 211802 186895 211858 186904
rect 210422 169144 210478 169153
rect 210422 169079 210478 169088
rect 210436 156466 210464 169079
rect 210424 156460 210476 156466
rect 210424 156402 210476 156408
rect 210436 155990 210464 156402
rect 210424 155984 210476 155990
rect 210424 155926 210476 155932
rect 209976 151786 210096 151814
rect 208860 147008 208912 147014
rect 208860 146950 208912 146956
rect 209872 147008 209924 147014
rect 209872 146950 209924 146956
rect 208872 140978 208900 146950
rect 209780 143676 209832 143682
rect 209780 143618 209832 143624
rect 207124 140950 207414 140978
rect 207768 140950 208150 140978
rect 208504 140950 208702 140978
rect 208872 140950 209254 140978
rect 206614 140542 206968 140570
rect 209792 140570 209820 143618
rect 210068 140978 210096 151786
rect 211816 147665 211844 186895
rect 213196 148481 213224 189722
rect 213276 175296 213328 175302
rect 213276 175238 213328 175244
rect 213182 148472 213238 148481
rect 213182 148407 213238 148416
rect 212354 147792 212410 147801
rect 212354 147727 212410 147736
rect 211802 147656 211858 147665
rect 211160 147620 211212 147626
rect 211802 147591 211858 147600
rect 211160 147562 211212 147568
rect 210700 147008 210752 147014
rect 210700 146950 210752 146956
rect 210712 140978 210740 146950
rect 211172 140978 211200 147562
rect 212368 142497 212396 147727
rect 213288 144809 213316 175238
rect 213840 149705 213868 227559
rect 214562 226944 214618 226953
rect 214562 226879 214618 226888
rect 214576 222193 214604 226879
rect 214562 222184 214618 222193
rect 214562 222119 214618 222128
rect 214010 175400 214066 175409
rect 214010 175335 214066 175344
rect 214024 151814 214052 175335
rect 214576 171193 214604 222119
rect 214668 202162 214696 234602
rect 215312 233209 215340 238002
rect 215484 237312 215536 237318
rect 215484 237254 215536 237260
rect 215496 236638 215524 237254
rect 216324 236638 216352 241604
rect 218072 241590 218730 241618
rect 217966 240816 218022 240825
rect 217966 240751 218022 240760
rect 217980 236638 218008 240751
rect 215484 236632 215536 236638
rect 215484 236574 215536 236580
rect 216312 236632 216364 236638
rect 216312 236574 216364 236580
rect 217968 236632 218020 236638
rect 217968 236574 218020 236580
rect 215298 233200 215354 233209
rect 215298 233135 215354 233144
rect 215206 232520 215262 232529
rect 215206 232455 215262 232464
rect 214656 202156 214708 202162
rect 214656 202098 214708 202104
rect 214562 171184 214618 171193
rect 214562 171119 214618 171128
rect 214576 157418 214604 171119
rect 214564 157412 214616 157418
rect 214564 157354 214616 157360
rect 215116 157412 215168 157418
rect 215116 157354 215168 157360
rect 214024 151786 214328 151814
rect 213826 149696 213882 149705
rect 213826 149631 213882 149640
rect 213460 146940 213512 146946
rect 213460 146882 213512 146888
rect 213274 144800 213330 144809
rect 213274 144735 213330 144744
rect 212354 142488 212410 142497
rect 212354 142423 212410 142432
rect 210068 140950 210542 140978
rect 210712 140950 211094 140978
rect 211172 140950 211646 140978
rect 212368 140964 212396 142423
rect 213288 140978 213316 144735
rect 213472 142254 213500 146882
rect 214012 143268 214064 143274
rect 214012 143210 214064 143216
rect 213460 142248 213512 142254
rect 213460 142190 213512 142196
rect 212934 140950 213316 140978
rect 213472 140964 213500 142190
rect 214024 140964 214052 143210
rect 214300 140978 214328 151786
rect 215128 143274 215156 157354
rect 215220 148345 215248 232455
rect 215392 167680 215444 167686
rect 215392 167622 215444 167628
rect 215300 167068 215352 167074
rect 215300 167010 215352 167016
rect 215312 164898 215340 167010
rect 215300 164892 215352 164898
rect 215300 164834 215352 164840
rect 215404 162926 215432 167622
rect 215392 162920 215444 162926
rect 215392 162862 215444 162868
rect 215206 148336 215262 148345
rect 215206 148271 215262 148280
rect 215220 147801 215248 148271
rect 215206 147792 215262 147801
rect 215206 147727 215262 147736
rect 215404 147014 215432 162862
rect 215496 147082 215524 236574
rect 215944 233912 215996 233918
rect 215944 233854 215996 233860
rect 215956 231810 215984 233854
rect 215944 231804 215996 231810
rect 215944 231746 215996 231752
rect 215956 164286 215984 231746
rect 215944 164280 215996 164286
rect 215944 164222 215996 164228
rect 215956 161474 215984 164222
rect 215588 161446 215984 161474
rect 215484 147076 215536 147082
rect 215484 147018 215536 147024
rect 215392 147008 215444 147014
rect 215392 146950 215444 146956
rect 215116 143268 215168 143274
rect 215116 143210 215168 143216
rect 215300 142180 215352 142186
rect 215300 142122 215352 142128
rect 214300 140950 214774 140978
rect 209792 140556 210096 140570
rect 209806 140554 210096 140556
rect 209806 140548 210108 140554
rect 209806 140542 210056 140548
rect 206558 140519 206614 140528
rect 210056 140490 210108 140496
rect 206558 140448 206614 140457
rect 196862 140406 197110 140434
rect 205652 140406 206558 140434
rect 196806 140383 196862 140392
rect 215312 140434 215340 142122
rect 215588 140978 215616 161446
rect 218072 154562 218100 241590
rect 218702 240816 218758 240825
rect 218702 240751 218758 240760
rect 218150 235240 218206 235249
rect 218150 235175 218206 235184
rect 218060 154556 218112 154562
rect 218060 154498 218112 154504
rect 218058 153096 218114 153105
rect 218058 153031 218114 153040
rect 216680 150476 216732 150482
rect 216680 150418 216732 150424
rect 216220 147008 216272 147014
rect 216220 146950 216272 146956
rect 216232 140978 216260 146950
rect 216692 140978 216720 150418
rect 218072 149326 218100 153031
rect 218164 151814 218192 235175
rect 218716 224777 218744 240751
rect 221108 239698 221136 241604
rect 219440 239692 219492 239698
rect 219440 239634 219492 239640
rect 221096 239692 221148 239698
rect 221096 239634 221148 239640
rect 219452 238814 219480 239634
rect 219440 238808 219492 238814
rect 219440 238750 219492 238756
rect 218702 224768 218758 224777
rect 218702 224703 218758 224712
rect 218716 214606 218744 224703
rect 218704 214600 218756 214606
rect 218704 214542 218756 214548
rect 219452 169017 219480 238750
rect 220912 236632 220964 236638
rect 222108 236632 222160 236638
rect 220912 236574 220964 236580
rect 222106 236600 222108 236609
rect 222160 236600 222162 236609
rect 219530 235240 219586 235249
rect 219530 235175 219586 235184
rect 219544 169833 219572 235175
rect 220818 217424 220874 217433
rect 220818 217359 220874 217368
rect 220832 176730 220860 217359
rect 220820 176724 220872 176730
rect 220820 176666 220872 176672
rect 220084 173936 220136 173942
rect 220084 173878 220136 173884
rect 219530 169824 219586 169833
rect 219530 169759 219586 169768
rect 219438 169008 219494 169017
rect 219438 168943 219494 168952
rect 218242 154592 218298 154601
rect 218242 154527 218298 154536
rect 218256 153105 218284 154527
rect 218242 153096 218298 153105
rect 218242 153031 218298 153040
rect 218164 151786 218284 151814
rect 218060 149320 218112 149326
rect 218060 149262 218112 149268
rect 217232 144968 217284 144974
rect 217232 144910 217284 144916
rect 217244 140978 217272 144910
rect 218256 142497 218284 151786
rect 218612 149320 218664 149326
rect 218612 149262 218664 149268
rect 218242 142488 218298 142497
rect 218242 142423 218298 142432
rect 218256 142322 218284 142423
rect 218244 142316 218296 142322
rect 218244 142258 218296 142264
rect 215588 140950 215878 140978
rect 216232 140950 216614 140978
rect 216692 140950 217166 140978
rect 217244 140950 217718 140978
rect 218256 140964 218284 142258
rect 218624 140978 218652 149262
rect 219532 143540 219584 143546
rect 219532 143482 219584 143488
rect 218624 140950 219006 140978
rect 219544 140964 219572 143482
rect 220096 143478 220124 173878
rect 220924 171134 220952 236574
rect 222106 236535 222162 236544
rect 223500 231849 223528 241604
rect 222842 231840 222898 231849
rect 222842 231775 222898 231784
rect 223486 231840 223542 231849
rect 223486 231775 223542 231784
rect 222292 202156 222344 202162
rect 222292 202098 222344 202104
rect 221464 176724 221516 176730
rect 221464 176666 221516 176672
rect 220924 171106 221044 171134
rect 220266 169824 220322 169833
rect 220266 169759 220322 169768
rect 220176 160744 220228 160750
rect 220176 160686 220228 160692
rect 220188 146266 220216 160686
rect 220280 154601 220308 169759
rect 220358 169008 220414 169017
rect 220358 168943 220414 168952
rect 220372 160138 220400 168943
rect 220360 160132 220412 160138
rect 220360 160074 220412 160080
rect 220266 154592 220322 154601
rect 220266 154527 220322 154536
rect 220176 146260 220228 146266
rect 220176 146202 220228 146208
rect 220280 143546 220308 154527
rect 220372 152590 220400 160074
rect 220820 158024 220872 158030
rect 220820 157966 220872 157972
rect 220360 152584 220412 152590
rect 220360 152526 220412 152532
rect 220268 143540 220320 143546
rect 220268 143482 220320 143488
rect 220084 143472 220136 143478
rect 220084 143414 220136 143420
rect 220096 140964 220124 143414
rect 220832 140964 220860 157966
rect 221016 149161 221044 171106
rect 221002 149152 221058 149161
rect 221002 149087 221058 149096
rect 220912 146260 220964 146266
rect 220912 146202 220964 146208
rect 220924 140978 220952 146202
rect 221476 142154 221504 176666
rect 222200 163532 222252 163538
rect 222200 163474 222252 163480
rect 222212 161537 222240 163474
rect 222198 161528 222254 161537
rect 222198 161463 222254 161472
rect 222014 149152 222070 149161
rect 222014 149087 222070 149096
rect 222028 146305 222056 149087
rect 222014 146296 222070 146305
rect 222014 146231 222070 146240
rect 221922 142216 221978 142225
rect 221922 142154 221978 142160
rect 221476 142151 221978 142154
rect 221476 142126 221964 142151
rect 220924 140950 221398 140978
rect 221936 140964 221964 142126
rect 222212 140978 222240 161463
rect 222304 144673 222332 202098
rect 222856 176390 222884 231775
rect 224316 231124 224368 231130
rect 224316 231066 224368 231072
rect 224224 227044 224276 227050
rect 224224 226986 224276 226992
rect 223580 188352 223632 188358
rect 223580 188294 223632 188300
rect 222844 176384 222896 176390
rect 222844 176326 222896 176332
rect 223592 173058 223620 188294
rect 223580 173052 223632 173058
rect 223580 172994 223632 173000
rect 223592 172650 223620 172994
rect 223580 172644 223632 172650
rect 223580 172586 223632 172592
rect 223670 166288 223726 166297
rect 223670 166223 223726 166232
rect 223580 153264 223632 153270
rect 223580 153206 223632 153212
rect 223592 147014 223620 153206
rect 223580 147008 223632 147014
rect 223580 146950 223632 146956
rect 222290 144664 222346 144673
rect 222290 144599 222346 144608
rect 223026 144664 223082 144673
rect 223026 144599 223082 144608
rect 223040 143721 223068 144599
rect 223026 143712 223082 143721
rect 223026 143647 223082 143656
rect 223040 141030 223068 143647
rect 223684 142866 223712 166223
rect 223672 142860 223724 142866
rect 223672 142802 223724 142808
rect 223684 142594 223712 142802
rect 223212 142588 223264 142594
rect 223212 142530 223264 142536
rect 223672 142588 223724 142594
rect 223672 142530 223724 142536
rect 223028 141024 223080 141030
rect 222212 140950 222502 140978
rect 223028 140966 223080 140972
rect 223224 140964 223252 142530
rect 223488 142180 223540 142186
rect 223488 142122 223540 142128
rect 223500 140758 223528 142122
rect 223578 140856 223634 140865
rect 224236 140842 224264 226986
rect 224328 202774 224356 231066
rect 225788 204944 225840 204950
rect 225788 204886 225840 204892
rect 225800 204406 225828 204886
rect 225144 204400 225196 204406
rect 225144 204342 225196 204348
rect 225788 204400 225840 204406
rect 225788 204342 225840 204348
rect 224316 202768 224368 202774
rect 224316 202710 224368 202716
rect 224960 176384 225012 176390
rect 224960 176326 225012 176332
rect 224316 173052 224368 173058
rect 224316 172994 224368 173000
rect 223634 140814 224264 140842
rect 223578 140791 223634 140800
rect 223488 140752 223540 140758
rect 223488 140694 223540 140700
rect 215392 140480 215444 140486
rect 215312 140428 215392 140434
rect 215312 140422 215444 140428
rect 224328 140434 224356 172994
rect 224972 161498 225000 176326
rect 224960 161492 225012 161498
rect 225012 161446 225092 161474
rect 224960 161434 225012 161440
rect 224960 147688 225012 147694
rect 224960 147630 225012 147636
rect 224500 147008 224552 147014
rect 224500 146950 224552 146956
rect 224512 140978 224540 146950
rect 224512 140950 224894 140978
rect 224498 140448 224554 140457
rect 215312 140420 215432 140422
rect 224328 140420 224498 140434
rect 215326 140406 215432 140420
rect 224342 140406 224498 140420
rect 206558 140383 206614 140392
rect 224498 140383 224554 140392
rect 193416 132466 193536 132494
rect 193416 126274 193444 132466
rect 193404 126268 193456 126274
rect 193404 126210 193456 126216
rect 193126 124944 193182 124953
rect 193126 124879 193182 124888
rect 193036 103488 193088 103494
rect 193036 103430 193088 103436
rect 193048 102649 193076 103430
rect 193034 102640 193090 102649
rect 193034 102575 193090 102584
rect 192942 86184 192998 86193
rect 192942 86119 192998 86128
rect 192852 68332 192904 68338
rect 192852 68274 192904 68280
rect 193048 49026 193076 102575
rect 193140 69698 193168 124879
rect 224972 122834 225000 147630
rect 225064 129033 225092 161446
rect 225050 129024 225106 129033
rect 225050 128959 225106 128968
rect 225156 122834 225184 204342
rect 225984 184210 226012 241604
rect 227076 238808 227128 238814
rect 227076 238750 227128 238756
rect 227088 220794 227116 238750
rect 228376 237046 228404 241604
rect 230768 238814 230796 241604
rect 233160 238814 233188 241604
rect 234620 240848 234672 240854
rect 234620 240790 234672 240796
rect 234632 240106 234660 240790
rect 233884 240100 233936 240106
rect 233884 240042 233936 240048
rect 234620 240100 234672 240106
rect 234620 240042 234672 240048
rect 230756 238808 230808 238814
rect 230756 238750 230808 238756
rect 233148 238808 233200 238814
rect 233148 238750 233200 238756
rect 233160 237386 233188 238750
rect 233148 237380 233200 237386
rect 233148 237322 233200 237328
rect 228364 237040 228416 237046
rect 228364 236982 228416 236988
rect 230480 237040 230532 237046
rect 230480 236982 230532 236988
rect 227718 234016 227774 234025
rect 227718 233951 227774 233960
rect 227076 220788 227128 220794
rect 227076 220730 227128 220736
rect 226984 220108 227036 220114
rect 226984 220050 227036 220056
rect 226432 199436 226484 199442
rect 226432 199378 226484 199384
rect 226340 196648 226392 196654
rect 226340 196590 226392 196596
rect 225972 184204 226024 184210
rect 225972 184146 226024 184152
rect 225236 143608 225288 143614
rect 225236 143550 225288 143556
rect 225248 132494 225276 143550
rect 225326 140176 225382 140185
rect 225326 140111 225382 140120
rect 225340 138990 225368 140111
rect 225328 138984 225380 138990
rect 225328 138926 225380 138932
rect 225248 132466 225460 132494
rect 225432 131102 225460 132466
rect 225420 131096 225472 131102
rect 225420 131038 225472 131044
rect 225432 130937 225460 131038
rect 225418 130928 225474 130937
rect 225418 130863 225474 130872
rect 226154 128480 226210 128489
rect 226154 128415 226210 128424
rect 226168 128382 226196 128415
rect 226156 128376 226208 128382
rect 226156 128318 226208 128324
rect 224972 122806 225092 122834
rect 225156 122806 225368 122834
rect 225064 113801 225092 122806
rect 225234 116784 225290 116793
rect 225234 116719 225290 116728
rect 225050 113792 225106 113801
rect 225050 113727 225106 113736
rect 225142 109712 225198 109721
rect 224972 109670 225142 109698
rect 193218 104136 193274 104145
rect 193218 104071 193274 104080
rect 193232 96393 193260 104071
rect 193218 96384 193274 96393
rect 193218 96319 193274 96328
rect 193232 95441 193260 96319
rect 193218 95432 193274 95441
rect 193218 95367 193274 95376
rect 193404 93900 193456 93906
rect 193404 93842 193456 93848
rect 193220 93832 193272 93838
rect 193220 93774 193272 93780
rect 193232 92313 193260 93774
rect 193416 93362 193444 93842
rect 199108 93424 199160 93430
rect 193784 93362 194166 93378
rect 221648 93424 221700 93430
rect 202234 93392 202290 93401
rect 199160 93372 199502 93378
rect 199108 93366 199502 93372
rect 193404 93356 193456 93362
rect 193404 93298 193456 93304
rect 193772 93356 194166 93362
rect 193824 93350 194166 93356
rect 199120 93364 199502 93366
rect 199120 93350 199516 93364
rect 193772 93298 193824 93304
rect 193324 92806 193614 92834
rect 193218 92304 193274 92313
rect 193218 92239 193274 92248
rect 193220 92132 193272 92138
rect 193220 92074 193272 92080
rect 193128 69692 193180 69698
rect 193128 69634 193180 69640
rect 193232 60042 193260 92074
rect 193324 63510 193352 92806
rect 193784 92138 193812 93298
rect 194718 92806 194824 92834
rect 194506 92712 194562 92721
rect 194506 92647 194562 92656
rect 193772 92132 193824 92138
rect 193772 92074 193824 92080
rect 194520 72457 194548 92647
rect 194692 91044 194744 91050
rect 194692 90986 194744 90992
rect 194506 72448 194562 72457
rect 194506 72383 194562 72392
rect 193312 63504 193364 63510
rect 193312 63446 193364 63452
rect 193220 60036 193272 60042
rect 193220 59978 193272 59984
rect 193324 59362 193352 63446
rect 194704 62014 194732 90986
rect 194796 69018 194824 92806
rect 195256 91050 195284 92820
rect 195244 91044 195296 91050
rect 195244 90986 195296 90992
rect 195992 84114 196020 92820
rect 196544 89593 196572 92820
rect 196530 89584 196586 89593
rect 196530 89519 196586 89528
rect 197096 86873 197124 92820
rect 197372 92806 197662 92834
rect 197082 86864 197138 86873
rect 197082 86799 197138 86808
rect 195980 84108 196032 84114
rect 195980 84050 196032 84056
rect 195992 82890 196020 84050
rect 195980 82884 196032 82890
rect 195980 82826 196032 82832
rect 196624 82884 196676 82890
rect 196624 82826 196676 82832
rect 194784 69012 194836 69018
rect 194784 68954 194836 68960
rect 195336 69012 195388 69018
rect 195336 68954 195388 68960
rect 195348 62014 195376 68954
rect 194692 62008 194744 62014
rect 194692 61950 194744 61956
rect 195336 62008 195388 62014
rect 195336 61950 195388 61956
rect 194704 60790 194732 61950
rect 194692 60784 194744 60790
rect 194692 60726 194744 60732
rect 195244 60784 195296 60790
rect 195244 60726 195296 60732
rect 193312 59356 193364 59362
rect 193312 59298 193364 59304
rect 193864 59356 193916 59362
rect 193864 59298 193916 59304
rect 193036 49020 193088 49026
rect 193036 48962 193088 48968
rect 193876 29646 193904 59298
rect 195256 31074 195284 60726
rect 195244 31068 195296 31074
rect 195244 31010 195296 31016
rect 193864 29640 193916 29646
rect 193864 29582 193916 29588
rect 196636 8974 196664 82826
rect 197372 67590 197400 92806
rect 198384 88233 198412 92820
rect 198950 92806 199424 92834
rect 198370 88224 198426 88233
rect 198370 88159 198426 88168
rect 199396 86970 199424 92806
rect 199384 86964 199436 86970
rect 199384 86906 199436 86912
rect 197360 67584 197412 67590
rect 197360 67526 197412 67532
rect 198004 67584 198056 67590
rect 198004 67526 198056 67532
rect 198016 56506 198044 67526
rect 198004 56500 198056 56506
rect 198004 56442 198056 56448
rect 199396 39370 199424 86906
rect 199488 86290 199516 93350
rect 202290 93350 202630 93378
rect 221398 93372 221648 93378
rect 221398 93366 221700 93372
rect 224774 93392 224830 93401
rect 221398 93350 221688 93366
rect 202234 93327 202290 93336
rect 224830 93350 224894 93378
rect 224774 93327 224830 93336
rect 224498 93256 224554 93265
rect 224342 93214 224498 93242
rect 224498 93191 224554 93200
rect 207664 93152 207716 93158
rect 207664 93094 207716 93100
rect 200302 92848 200358 92857
rect 200132 92806 200238 92834
rect 199476 86284 199528 86290
rect 199476 86226 199528 86232
rect 200132 59226 200160 92806
rect 201038 92848 201094 92857
rect 200302 92783 200358 92792
rect 200316 84194 200344 92783
rect 200776 92177 200804 92820
rect 201094 92806 201342 92834
rect 201512 92806 201894 92834
rect 203182 92806 203564 92834
rect 201038 92783 201094 92792
rect 200762 92168 200818 92177
rect 200762 92103 200818 92112
rect 200224 84166 200344 84194
rect 200224 76566 200252 84166
rect 200212 76560 200264 76566
rect 200212 76502 200264 76508
rect 201512 67590 201540 92806
rect 203536 90409 203564 92806
rect 203720 90681 203748 92820
rect 203706 90672 203762 90681
rect 203706 90607 203762 90616
rect 203522 90400 203578 90409
rect 203522 90335 203578 90344
rect 203536 79558 203564 90335
rect 203720 81297 203748 90607
rect 204456 90545 204484 92820
rect 204442 90536 204498 90545
rect 204442 90471 204498 90480
rect 204352 89820 204404 89826
rect 204352 89762 204404 89768
rect 203706 81288 203762 81297
rect 203706 81223 203762 81232
rect 204168 79960 204220 79966
rect 204168 79902 204220 79908
rect 204180 79558 204208 79902
rect 203524 79552 203576 79558
rect 203524 79494 203576 79500
rect 204168 79552 204220 79558
rect 204168 79494 204220 79500
rect 201500 67584 201552 67590
rect 201500 67526 201552 67532
rect 202144 67584 202196 67590
rect 202144 67526 202196 67532
rect 200120 59220 200172 59226
rect 200120 59162 200172 59168
rect 200132 57866 200160 59162
rect 200120 57860 200172 57866
rect 200120 57802 200172 57808
rect 200764 57860 200816 57866
rect 200764 57802 200816 57808
rect 199384 39364 199436 39370
rect 199384 39306 199436 39312
rect 200776 33794 200804 57802
rect 202156 56574 202184 67526
rect 202144 56568 202196 56574
rect 202144 56510 202196 56516
rect 200764 33788 200816 33794
rect 200764 33730 200816 33736
rect 202156 10334 202184 56510
rect 204180 21418 204208 79494
rect 204364 60654 204392 89762
rect 204456 87553 204484 90471
rect 204904 89752 204956 89758
rect 204904 89694 204956 89700
rect 204442 87544 204498 87553
rect 204442 87479 204498 87488
rect 204916 81326 204944 89694
rect 205008 85474 205036 92820
rect 205560 92177 205588 92820
rect 206112 92449 206140 92820
rect 206098 92440 206154 92449
rect 205640 92404 205692 92410
rect 206098 92375 206154 92384
rect 205640 92346 205692 92352
rect 205546 92168 205602 92177
rect 205546 92103 205602 92112
rect 205560 89826 205588 92103
rect 205652 92041 205680 92346
rect 205638 92032 205694 92041
rect 205638 91967 205694 91976
rect 205640 91792 205692 91798
rect 205640 91734 205692 91740
rect 205548 89820 205600 89826
rect 205548 89762 205600 89768
rect 205652 88262 205680 91734
rect 205640 88256 205692 88262
rect 205640 88198 205692 88204
rect 206848 87650 206876 92820
rect 207124 92806 207414 92834
rect 206836 87644 206888 87650
rect 206836 87586 206888 87592
rect 204996 85468 205048 85474
rect 204996 85410 205048 85416
rect 206848 84862 206876 87586
rect 206836 84856 206888 84862
rect 206836 84798 206888 84804
rect 204904 81320 204956 81326
rect 204904 81262 204956 81268
rect 204352 60648 204404 60654
rect 204352 60590 204404 60596
rect 204364 60246 204392 60590
rect 204352 60240 204404 60246
rect 204352 60182 204404 60188
rect 204168 21412 204220 21418
rect 204168 21354 204220 21360
rect 202144 10328 202196 10334
rect 202144 10270 202196 10276
rect 196624 8968 196676 8974
rect 196624 8910 196676 8916
rect 191748 7608 191800 7614
rect 191748 7550 191800 7556
rect 204916 4826 204944 81262
rect 204996 60240 205048 60246
rect 204996 60182 205048 60188
rect 205008 14482 205036 60182
rect 207124 59362 207152 92806
rect 207676 77217 207704 93094
rect 210422 92984 210478 92993
rect 210358 92956 210422 92970
rect 210344 92942 210422 92956
rect 208398 92848 208454 92857
rect 207952 89758 207980 92820
rect 208454 92820 208702 92834
rect 208454 92806 208716 92820
rect 208398 92783 208454 92792
rect 208688 90273 208716 92806
rect 208674 90264 208730 90273
rect 208674 90199 208730 90208
rect 207940 89752 207992 89758
rect 207940 89694 207992 89700
rect 209240 87961 209268 92820
rect 209806 92806 209912 92834
rect 209686 90264 209742 90273
rect 209686 90199 209742 90208
rect 209226 87952 209282 87961
rect 209226 87887 209282 87896
rect 207662 77208 207718 77217
rect 207662 77143 207718 77152
rect 207112 59356 207164 59362
rect 207112 59298 207164 59304
rect 207664 59356 207716 59362
rect 207664 59298 207716 59304
rect 207676 24138 207704 59298
rect 209700 25566 209728 90199
rect 209884 84114 209912 92806
rect 210344 89865 210372 92942
rect 210422 92919 210478 92928
rect 224038 92848 224094 92857
rect 210436 92806 211094 92834
rect 210330 89856 210386 89865
rect 210330 89791 210386 89800
rect 210436 84194 210464 92806
rect 211632 89729 211660 92820
rect 212184 92721 212212 92820
rect 212170 92712 212226 92721
rect 212170 92647 212226 92656
rect 212184 90953 212212 92647
rect 212170 90944 212226 90953
rect 212170 90879 212226 90888
rect 212920 90370 212948 92820
rect 213012 92806 213486 92834
rect 213932 92806 214038 92834
rect 212908 90364 212960 90370
rect 212908 90306 212960 90312
rect 211618 89720 211674 89729
rect 211618 89655 211674 89664
rect 212920 86970 212948 90306
rect 212908 86964 212960 86970
rect 212908 86906 212960 86912
rect 213012 84194 213040 92806
rect 213828 86964 213880 86970
rect 213828 86906 213880 86912
rect 210068 84166 210464 84194
rect 212644 84166 213040 84194
rect 209872 84108 209924 84114
rect 209872 84050 209924 84056
rect 210068 79937 210096 84166
rect 210424 84108 210476 84114
rect 210424 84050 210476 84056
rect 210054 79928 210110 79937
rect 210054 79863 210110 79872
rect 210436 74526 210464 84050
rect 212644 74526 212672 84166
rect 210424 74520 210476 74526
rect 210424 74462 210476 74468
rect 212632 74520 212684 74526
rect 212632 74462 212684 74468
rect 212644 73234 212672 74462
rect 212632 73228 212684 73234
rect 212632 73170 212684 73176
rect 213184 73228 213236 73234
rect 213184 73170 213236 73176
rect 213196 64870 213224 73170
rect 213184 64864 213236 64870
rect 213184 64806 213236 64812
rect 213196 28286 213224 64806
rect 213184 28280 213236 28286
rect 213184 28222 213236 28228
rect 209688 25560 209740 25566
rect 209688 25502 209740 25508
rect 207664 24132 207716 24138
rect 207664 24074 207716 24080
rect 213840 22778 213868 86906
rect 213932 84182 213960 92806
rect 214576 92449 214604 92820
rect 215326 92806 215432 92834
rect 215878 92806 216076 92834
rect 214562 92440 214618 92449
rect 214562 92375 214618 92384
rect 215298 90264 215354 90273
rect 215298 90199 215354 90208
rect 213920 84176 213972 84182
rect 213920 84118 213972 84124
rect 214656 77988 214708 77994
rect 214656 77930 214708 77936
rect 214564 65544 214616 65550
rect 214564 65486 214616 65492
rect 214576 36582 214604 65486
rect 214668 53106 214696 77930
rect 215312 73166 215340 90199
rect 215404 88330 215432 92806
rect 215392 88324 215444 88330
rect 215392 88266 215444 88272
rect 216048 84250 216076 92806
rect 216416 90273 216444 92820
rect 217166 92806 217364 92834
rect 218348 92820 218822 92834
rect 217336 91050 217364 92806
rect 217324 91044 217376 91050
rect 217324 90986 217376 90992
rect 216402 90264 216458 90273
rect 216402 90199 216458 90208
rect 216036 84244 216088 84250
rect 216036 84186 216088 84192
rect 215300 73160 215352 73166
rect 215300 73102 215352 73108
rect 215312 71806 215340 73102
rect 215300 71800 215352 71806
rect 215300 71742 215352 71748
rect 215944 71800 215996 71806
rect 215944 71742 215996 71748
rect 214656 53100 214708 53106
rect 214656 53042 214708 53048
rect 214564 36576 214616 36582
rect 214564 36518 214616 36524
rect 213828 22772 213880 22778
rect 213828 22714 213880 22720
rect 204996 14476 205048 14482
rect 204996 14418 205048 14424
rect 215956 11762 215984 71742
rect 216048 62082 216076 84186
rect 217336 63442 217364 90986
rect 217704 89690 217732 92820
rect 217692 89684 217744 89690
rect 217692 89626 217744 89632
rect 218256 89622 218284 92820
rect 218348 92806 218836 92820
rect 219558 92806 220032 92834
rect 218244 89616 218296 89622
rect 218244 89558 218296 89564
rect 218348 84194 218376 92806
rect 218808 92585 218836 92806
rect 218794 92576 218850 92585
rect 218794 92511 218850 92520
rect 220004 89690 220032 92806
rect 219992 89684 220044 89690
rect 219992 89626 220044 89632
rect 220004 85354 220032 89626
rect 220096 85513 220124 92820
rect 220648 85542 220676 92820
rect 221936 86737 221964 92820
rect 222212 92806 222502 92834
rect 222672 92806 223054 92834
rect 223790 92820 224038 92834
rect 223776 92806 224038 92820
rect 221922 86728 221978 86737
rect 221922 86663 221978 86672
rect 220636 85536 220688 85542
rect 220082 85504 220138 85513
rect 220636 85478 220688 85484
rect 220082 85439 220138 85448
rect 220004 85326 220216 85354
rect 220084 84856 220136 84862
rect 220084 84798 220136 84804
rect 218072 84166 218376 84194
rect 218072 71670 218100 84166
rect 218060 71664 218112 71670
rect 218060 71606 218112 71612
rect 218336 71664 218388 71670
rect 218336 71606 218388 71612
rect 218348 71058 218376 71606
rect 218336 71052 218388 71058
rect 218336 70994 218388 71000
rect 217324 63436 217376 63442
rect 217324 63378 217376 63384
rect 216036 62076 216088 62082
rect 216036 62018 216088 62024
rect 217336 46238 217364 63378
rect 217324 46232 217376 46238
rect 217324 46174 217376 46180
rect 215944 11756 215996 11762
rect 215944 11698 215996 11704
rect 204904 4820 204956 4826
rect 204904 4762 204956 4768
rect 220096 3466 220124 84798
rect 220188 80073 220216 85326
rect 220174 80064 220230 80073
rect 220174 79999 220230 80008
rect 222212 57934 222240 92806
rect 222672 84194 222700 92806
rect 223776 90302 223804 92806
rect 224038 92783 224094 92792
rect 223764 90296 223816 90302
rect 223764 90238 223816 90244
rect 224868 90296 224920 90302
rect 224868 90238 224920 90244
rect 222304 84166 222700 84194
rect 222304 70378 222332 84166
rect 222292 70372 222344 70378
rect 222292 70314 222344 70320
rect 222844 70372 222896 70378
rect 222844 70314 222896 70320
rect 222200 57928 222252 57934
rect 222200 57870 222252 57876
rect 222856 18630 222884 70314
rect 222936 57928 222988 57934
rect 222936 57870 222988 57876
rect 222948 35222 222976 57870
rect 222936 35216 222988 35222
rect 222936 35158 222988 35164
rect 222844 18624 222896 18630
rect 222844 18566 222896 18572
rect 224880 6186 224908 90238
rect 224972 82822 225000 109670
rect 225142 109647 225198 109656
rect 225248 108338 225276 116719
rect 225064 108310 225276 108338
rect 225064 93158 225092 108310
rect 225340 103514 225368 122806
rect 225156 103486 225368 103514
rect 225156 93430 225184 103486
rect 226248 97980 226300 97986
rect 226248 97922 226300 97928
rect 226260 97209 226288 97922
rect 225234 97200 225290 97209
rect 225234 97135 225290 97144
rect 226246 97200 226302 97209
rect 226246 97135 226302 97144
rect 225144 93424 225196 93430
rect 225144 93366 225196 93372
rect 225052 93152 225104 93158
rect 225052 93094 225104 93100
rect 225248 92410 225276 97135
rect 226352 95169 226380 196590
rect 226444 137170 226472 199378
rect 226996 191146 227024 220050
rect 226984 191140 227036 191146
rect 226984 191082 227036 191088
rect 226524 180124 226576 180130
rect 226524 180066 226576 180072
rect 226536 137442 226564 180066
rect 227732 156097 227760 233951
rect 230386 225584 230442 225593
rect 230386 225519 230442 225528
rect 230400 223553 230428 225519
rect 229098 223544 229154 223553
rect 229098 223479 229154 223488
rect 230386 223544 230442 223553
rect 230386 223479 230442 223488
rect 227812 221468 227864 221474
rect 227812 221410 227864 221416
rect 227824 220833 227852 221410
rect 227810 220824 227866 220833
rect 227810 220759 227866 220768
rect 227824 162897 227852 220759
rect 227810 162888 227866 162897
rect 227810 162823 227866 162832
rect 227718 156088 227774 156097
rect 227718 156023 227774 156032
rect 227732 147098 227760 156023
rect 227824 147218 227852 162823
rect 229112 158817 229140 223479
rect 229098 158808 229154 158817
rect 229098 158743 229154 158752
rect 227994 150512 228050 150521
rect 227994 150447 228050 150456
rect 227812 147212 227864 147218
rect 227812 147154 227864 147160
rect 227732 147070 227852 147098
rect 227720 147008 227772 147014
rect 227720 146950 227772 146956
rect 226798 146568 226854 146577
rect 226798 146503 226854 146512
rect 226536 137414 226748 137442
rect 226522 137184 226578 137193
rect 226444 137142 226522 137170
rect 226522 137119 226578 137128
rect 226536 135930 226564 137119
rect 226524 135924 226576 135930
rect 226524 135866 226576 135872
rect 226524 135652 226576 135658
rect 226524 135594 226576 135600
rect 226536 135561 226564 135594
rect 226522 135552 226578 135561
rect 226522 135487 226578 135496
rect 226720 134745 226748 137414
rect 226812 136377 226840 146503
rect 227626 139088 227682 139097
rect 227732 139074 227760 146950
rect 227682 139046 227760 139074
rect 227626 139023 227682 139032
rect 227720 138984 227772 138990
rect 227720 138926 227772 138932
rect 226798 136368 226854 136377
rect 226798 136303 226854 136312
rect 226706 134736 226762 134745
rect 226706 134671 226762 134680
rect 226982 134736 227038 134745
rect 226982 134671 227038 134680
rect 226708 133884 226760 133890
rect 226708 133826 226760 133832
rect 226720 133657 226748 133826
rect 226892 133816 226944 133822
rect 226892 133758 226944 133764
rect 226706 133648 226762 133657
rect 226706 133583 226762 133592
rect 226904 132841 226932 133758
rect 226890 132832 226946 132841
rect 226890 132767 226946 132776
rect 226708 132456 226760 132462
rect 226708 132398 226760 132404
rect 226720 132025 226748 132398
rect 226706 132016 226762 132025
rect 226706 131951 226762 131960
rect 226616 131028 226668 131034
rect 226616 130970 226668 130976
rect 226628 130121 226656 130970
rect 226614 130112 226670 130121
rect 226614 130047 226670 130056
rect 226616 128308 226668 128314
rect 226616 128250 226668 128256
rect 226628 127401 226656 128250
rect 226614 127392 226670 127401
rect 226614 127327 226670 127336
rect 226432 126948 226484 126954
rect 226432 126890 226484 126896
rect 226444 125769 226472 126890
rect 226892 126880 226944 126886
rect 226892 126822 226944 126828
rect 226904 126585 226932 126822
rect 226890 126576 226946 126585
rect 226890 126511 226946 126520
rect 226430 125760 226486 125769
rect 226430 125695 226486 125704
rect 226616 125588 226668 125594
rect 226616 125530 226668 125536
rect 226628 124681 226656 125530
rect 226614 124672 226670 124681
rect 226614 124607 226670 124616
rect 226708 124160 226760 124166
rect 226708 124102 226760 124108
rect 226524 123888 226576 123894
rect 226522 123856 226524 123865
rect 226576 123856 226578 123865
rect 226522 123791 226578 123800
rect 226720 123049 226748 124102
rect 226706 123040 226762 123049
rect 226706 122975 226762 122984
rect 226524 122800 226576 122806
rect 226524 122742 226576 122748
rect 226536 122233 226564 122742
rect 226522 122224 226578 122233
rect 226522 122159 226578 122168
rect 226996 122126 227024 134671
rect 227168 129328 227220 129334
rect 227166 129296 227168 129305
rect 227220 129296 227222 129305
rect 227166 129231 227222 129240
rect 227536 126880 227588 126886
rect 227536 126822 227588 126828
rect 226984 122120 227036 122126
rect 226984 122062 227036 122068
rect 226708 121440 226760 121446
rect 226708 121382 226760 121388
rect 226720 120329 226748 121382
rect 226706 120320 226762 120329
rect 226706 120255 226762 120264
rect 226706 118416 226762 118425
rect 226706 118351 226762 118360
rect 226614 117600 226670 117609
rect 226614 117535 226670 117544
rect 226628 117366 226656 117535
rect 226616 117360 226668 117366
rect 226616 117302 226668 117308
rect 226720 117026 226748 118351
rect 227548 117978 227576 126822
rect 227536 117972 227588 117978
rect 227536 117914 227588 117920
rect 226708 117020 226760 117026
rect 226708 116962 226760 116968
rect 226708 116000 226760 116006
rect 226706 115968 226708 115977
rect 226760 115968 226762 115977
rect 226706 115903 226762 115912
rect 226706 114880 226762 114889
rect 226706 114815 226762 114824
rect 226720 114578 226748 114815
rect 226708 114572 226760 114578
rect 226708 114514 226760 114520
rect 226616 114504 226668 114510
rect 226616 114446 226668 114452
rect 226628 114073 226656 114446
rect 226614 114064 226670 114073
rect 226614 113999 226670 114008
rect 226706 112160 226762 112169
rect 226706 112095 226762 112104
rect 226720 111858 226748 112095
rect 226708 111852 226760 111858
rect 226708 111794 226760 111800
rect 227732 111110 227760 138926
rect 227824 138689 227852 147070
rect 228008 142154 228036 150447
rect 227916 142126 228036 142154
rect 227810 138680 227866 138689
rect 227810 138615 227866 138624
rect 227916 133822 227944 142126
rect 227996 141024 228048 141030
rect 227996 140966 228048 140972
rect 227904 133816 227956 133822
rect 227904 133758 227956 133764
rect 228008 129334 228036 140966
rect 229112 132462 229140 158743
rect 230492 155922 230520 236982
rect 232502 222864 232558 222873
rect 232502 222799 232558 222808
rect 231124 188352 231176 188358
rect 231124 188294 231176 188300
rect 230480 155916 230532 155922
rect 230480 155858 230532 155864
rect 229190 146432 229246 146441
rect 229190 146367 229246 146376
rect 229100 132456 229152 132462
rect 229100 132398 229152 132404
rect 227996 129328 228048 129334
rect 227996 129270 228048 129276
rect 228008 127702 228036 129270
rect 227996 127696 228048 127702
rect 227996 127638 228048 127644
rect 229204 123894 229232 146367
rect 231136 144945 231164 188294
rect 232516 187678 232544 222799
rect 232596 218816 232648 218822
rect 232596 218758 232648 218764
rect 232608 209778 232636 218758
rect 232596 209772 232648 209778
rect 232596 209714 232648 209720
rect 232504 187672 232556 187678
rect 232504 187614 232556 187620
rect 231860 164892 231912 164898
rect 231860 164834 231912 164840
rect 231768 155916 231820 155922
rect 231768 155858 231820 155864
rect 231780 155310 231808 155858
rect 231768 155304 231820 155310
rect 231768 155246 231820 155252
rect 231766 148472 231822 148481
rect 231766 148407 231822 148416
rect 230478 144936 230534 144945
rect 230478 144871 230534 144880
rect 231122 144936 231178 144945
rect 231122 144871 231178 144880
rect 229282 143576 229338 143585
rect 229282 143511 229338 143520
rect 229296 133890 229324 143511
rect 230492 135658 230520 144871
rect 231780 143585 231808 148407
rect 231766 143576 231822 143585
rect 231766 143511 231822 143520
rect 230480 135652 230532 135658
rect 230480 135594 230532 135600
rect 229284 133884 229336 133890
rect 229284 133826 229336 133832
rect 230388 129056 230440 129062
rect 230388 128998 230440 129004
rect 230400 126886 230428 128998
rect 231872 128314 231900 164834
rect 233240 164348 233292 164354
rect 233240 164290 233292 164296
rect 232504 147756 232556 147762
rect 232504 147698 232556 147704
rect 232516 135250 232544 147698
rect 232504 135244 232556 135250
rect 232504 135186 232556 135192
rect 231860 128308 231912 128314
rect 231860 128250 231912 128256
rect 233148 128308 233200 128314
rect 233148 128250 233200 128256
rect 233160 127634 233188 128250
rect 233148 127628 233200 127634
rect 233148 127570 233200 127576
rect 230388 126880 230440 126886
rect 230388 126822 230440 126828
rect 233252 124166 233280 164290
rect 233240 124160 233292 124166
rect 233240 124102 233292 124108
rect 229192 123888 229244 123894
rect 229192 123830 229244 123836
rect 230480 117020 230532 117026
rect 230480 116962 230532 116968
rect 231124 117020 231176 117026
rect 231124 116962 231176 116968
rect 230388 116680 230440 116686
rect 230388 116622 230440 116628
rect 230400 116006 230428 116622
rect 229100 116000 229152 116006
rect 229100 115942 229152 115948
rect 230388 116000 230440 116006
rect 230388 115942 230440 115948
rect 227076 111104 227128 111110
rect 227076 111046 227128 111052
rect 227720 111104 227772 111110
rect 227720 111046 227772 111052
rect 227088 110537 227116 111046
rect 227718 110800 227774 110809
rect 227718 110735 227774 110744
rect 227074 110528 227130 110537
rect 227074 110463 227130 110472
rect 227732 110430 227760 110735
rect 227720 110424 227772 110430
rect 227720 110366 227772 110372
rect 228364 110424 228416 110430
rect 228364 110366 228416 110372
rect 226432 108996 226484 109002
rect 226432 108938 226484 108944
rect 226444 108633 226472 108938
rect 226430 108624 226486 108633
rect 226430 108559 226486 108568
rect 226706 107808 226762 107817
rect 226706 107743 226762 107752
rect 226720 107710 226748 107743
rect 226708 107704 226760 107710
rect 226708 107646 226760 107652
rect 226800 107636 226852 107642
rect 226800 107578 226852 107584
rect 226812 107001 226840 107578
rect 226798 106992 226854 107001
rect 226798 106927 226854 106936
rect 226706 105904 226762 105913
rect 226706 105839 226762 105848
rect 226720 105602 226748 105839
rect 226708 105596 226760 105602
rect 226708 105538 226760 105544
rect 226430 105088 226486 105097
rect 226430 105023 226486 105032
rect 226338 95160 226394 95169
rect 226338 95095 226394 95104
rect 226352 94489 226380 95095
rect 226338 94480 226394 94489
rect 226338 94415 226394 94424
rect 225236 92404 225288 92410
rect 225236 92346 225288 92352
rect 226444 88262 226472 105023
rect 226706 104272 226762 104281
rect 226706 104207 226762 104216
rect 226720 103562 226748 104207
rect 226708 103556 226760 103562
rect 226708 103498 226760 103504
rect 226614 103456 226670 103465
rect 226614 103391 226670 103400
rect 226628 102270 226656 103391
rect 226706 102368 226762 102377
rect 226706 102303 226762 102312
rect 226616 102264 226668 102270
rect 226616 102206 226668 102212
rect 226720 102202 226748 102303
rect 226708 102196 226760 102202
rect 226708 102138 226760 102144
rect 226524 102128 226576 102134
rect 226524 102070 226576 102076
rect 226536 101561 226564 102070
rect 226522 101552 226578 101561
rect 226522 101487 226578 101496
rect 226706 100736 226762 100745
rect 226706 100671 226762 100680
rect 226614 99648 226670 99657
rect 226614 99583 226670 99592
rect 226628 99414 226656 99583
rect 226720 99482 226748 100671
rect 226708 99476 226760 99482
rect 226708 99418 226760 99424
rect 226616 99408 226668 99414
rect 226616 99350 226668 99356
rect 226628 92478 226656 99350
rect 227352 98660 227404 98666
rect 227352 98602 227404 98608
rect 227364 98025 227392 98602
rect 227350 98016 227406 98025
rect 227350 97951 227406 97960
rect 227718 98016 227774 98025
rect 227718 97951 227774 97960
rect 226708 96620 226760 96626
rect 226708 96562 226760 96568
rect 226720 96121 226748 96562
rect 226706 96112 226762 96121
rect 226706 96047 226762 96056
rect 226892 95940 226944 95946
rect 226892 95882 226944 95888
rect 226904 93673 226932 95882
rect 227534 95160 227590 95169
rect 227534 95095 227590 95104
rect 226890 93664 226946 93673
rect 226890 93599 226946 93608
rect 226616 92472 226668 92478
rect 226616 92414 226668 92420
rect 226432 88256 226484 88262
rect 226432 88198 226484 88204
rect 227548 87650 227576 95095
rect 227536 87644 227588 87650
rect 227536 87586 227588 87592
rect 224960 82816 225012 82822
rect 224960 82758 225012 82764
rect 227732 64802 227760 97951
rect 227810 95840 227866 95849
rect 227810 95775 227866 95784
rect 227824 84153 227852 95775
rect 227810 84144 227866 84153
rect 227810 84079 227866 84088
rect 228376 71738 228404 110366
rect 229112 75857 229140 115942
rect 229192 99476 229244 99482
rect 229192 99418 229244 99424
rect 229204 77246 229232 99418
rect 230492 80034 230520 116962
rect 231136 116618 231164 116962
rect 231124 116612 231176 116618
rect 231124 116554 231176 116560
rect 233240 115252 233292 115258
rect 233240 115194 233292 115200
rect 233252 114578 233280 115194
rect 233240 114572 233292 114578
rect 233240 114514 233292 114520
rect 231952 111852 232004 111858
rect 231952 111794 232004 111800
rect 231768 108316 231820 108322
rect 231768 108258 231820 108264
rect 231780 107710 231808 108258
rect 230572 107704 230624 107710
rect 230572 107646 230624 107652
rect 231768 107704 231820 107710
rect 231768 107646 231820 107652
rect 230480 80028 230532 80034
rect 230480 79970 230532 79976
rect 229192 77240 229244 77246
rect 229192 77182 229244 77188
rect 229098 75848 229154 75857
rect 229098 75783 229154 75792
rect 230584 75721 230612 107646
rect 231860 102264 231912 102270
rect 231860 102206 231912 102212
rect 230570 75712 230626 75721
rect 230570 75647 230626 75656
rect 228364 71732 228416 71738
rect 228364 71674 228416 71680
rect 231872 67522 231900 102206
rect 231964 92313 231992 111794
rect 233148 102808 233200 102814
rect 233148 102750 233200 102756
rect 233160 102270 233188 102750
rect 233148 102264 233200 102270
rect 233148 102206 233200 102212
rect 231950 92304 232006 92313
rect 231950 92239 232006 92248
rect 233252 77081 233280 114514
rect 233896 110430 233924 240042
rect 235552 223582 235580 241604
rect 237380 238808 237432 238814
rect 237380 238750 237432 238756
rect 235908 229764 235960 229770
rect 235908 229706 235960 229712
rect 234620 223576 234672 223582
rect 234620 223518 234672 223524
rect 235540 223576 235592 223582
rect 235540 223518 235592 223524
rect 234632 158001 234660 223518
rect 234618 157992 234674 158001
rect 234618 157927 234674 157936
rect 235264 113824 235316 113830
rect 235264 113766 235316 113772
rect 233884 110424 233936 110430
rect 233884 110366 233936 110372
rect 233332 104168 233384 104174
rect 233332 104110 233384 104116
rect 233344 103562 233372 104110
rect 233332 103556 233384 103562
rect 233332 103498 233384 103504
rect 233344 81394 233372 103498
rect 235276 86970 235304 113766
rect 235920 104174 235948 229706
rect 236000 218748 236052 218754
rect 236000 218690 236052 218696
rect 236012 217977 236040 218690
rect 235998 217968 236054 217977
rect 235998 217903 236054 217912
rect 237286 217968 237342 217977
rect 237286 217903 237342 217912
rect 236644 212288 236696 212294
rect 236644 212230 236696 212236
rect 236000 162852 236052 162858
rect 236000 162794 236052 162800
rect 236012 161566 236040 162794
rect 236000 161560 236052 161566
rect 236000 161502 236052 161508
rect 236012 122806 236040 161502
rect 236000 122800 236052 122806
rect 236000 122742 236052 122748
rect 235908 104168 235960 104174
rect 235908 104110 235960 104116
rect 236656 98666 236684 212230
rect 237300 178702 237328 217903
rect 236736 178696 236788 178702
rect 236736 178638 236788 178644
rect 237288 178696 237340 178702
rect 237288 178638 237340 178644
rect 236748 162858 236776 178638
rect 236736 162852 236788 162858
rect 236736 162794 236788 162800
rect 236736 109744 236788 109750
rect 236736 109686 236788 109692
rect 236644 98660 236696 98666
rect 236644 98602 236696 98608
rect 236748 89729 236776 109686
rect 236734 89720 236790 89729
rect 236734 89655 236790 89664
rect 235264 86964 235316 86970
rect 235264 86906 235316 86912
rect 233332 81388 233384 81394
rect 233332 81330 233384 81336
rect 237392 79966 237420 238750
rect 237944 223582 237972 241604
rect 240152 241590 240350 241618
rect 240152 238754 240180 241590
rect 242728 240106 242756 241604
rect 242164 240100 242216 240106
rect 242164 240042 242216 240048
rect 242716 240100 242768 240106
rect 242716 240042 242768 240048
rect 240060 238726 240180 238754
rect 237472 223576 237524 223582
rect 237472 223518 237524 223524
rect 237932 223576 237984 223582
rect 237932 223518 237984 223524
rect 237484 212294 237512 223518
rect 237656 214600 237708 214606
rect 237656 214542 237708 214548
rect 237472 212288 237524 212294
rect 237472 212230 237524 212236
rect 237564 102196 237616 102202
rect 237564 102138 237616 102144
rect 237380 79960 237432 79966
rect 237380 79902 237432 79908
rect 233238 77072 233294 77081
rect 233238 77007 233294 77016
rect 237576 73098 237604 102138
rect 237668 97986 237696 214542
rect 240060 161474 240088 238726
rect 240138 220144 240194 220153
rect 240138 220079 240194 220088
rect 239968 161446 240088 161474
rect 239968 153270 239996 161446
rect 239956 153264 240008 153270
rect 240152 153241 240180 220079
rect 239956 153206 240008 153212
rect 240138 153232 240194 153241
rect 239968 152522 239996 153206
rect 240138 153167 240194 153176
rect 239956 152516 240008 152522
rect 239956 152458 240008 152464
rect 239404 135924 239456 135930
rect 239404 135866 239456 135872
rect 239416 120766 239444 135866
rect 240152 121446 240180 153167
rect 240784 144220 240836 144226
rect 240784 144162 240836 144168
rect 240796 143546 240824 144162
rect 240784 143540 240836 143546
rect 240784 143482 240836 143488
rect 240140 121440 240192 121446
rect 240140 121382 240192 121388
rect 239404 120760 239456 120766
rect 239404 120702 239456 120708
rect 239404 111172 239456 111178
rect 239404 111114 239456 111120
rect 237656 97980 237708 97986
rect 237656 97922 237708 97928
rect 239416 90953 239444 111114
rect 239402 90944 239458 90953
rect 239402 90879 239458 90888
rect 237564 73092 237616 73098
rect 237564 73034 237616 73040
rect 237576 71806 237604 73034
rect 237564 71800 237616 71806
rect 237564 71742 237616 71748
rect 238024 71800 238076 71806
rect 238024 71742 238076 71748
rect 231860 67516 231912 67522
rect 231860 67458 231912 67464
rect 227720 64796 227772 64802
rect 227720 64738 227772 64744
rect 227732 63578 227760 64738
rect 227720 63572 227772 63578
rect 227720 63514 227772 63520
rect 228364 63572 228416 63578
rect 228364 63514 228416 63520
rect 226984 47592 227036 47598
rect 226984 47534 227036 47540
rect 224868 6180 224920 6186
rect 224868 6122 224920 6128
rect 220084 3460 220136 3466
rect 220084 3402 220136 3408
rect 226996 2106 227024 47534
rect 228376 17270 228404 63514
rect 233884 39364 233936 39370
rect 233884 39306 233936 39312
rect 228364 17264 228416 17270
rect 228364 17206 228416 17212
rect 233896 4078 233924 39306
rect 238036 4418 238064 71742
rect 239416 40730 239444 90879
rect 239404 40724 239456 40730
rect 239404 40666 239456 40672
rect 240796 15910 240824 143482
rect 242176 113830 242204 240042
rect 243636 235272 243688 235278
rect 243636 235214 243688 235220
rect 242808 225616 242860 225622
rect 242808 225558 242860 225564
rect 242820 225010 242848 225558
rect 242256 225004 242308 225010
rect 242256 224946 242308 224952
rect 242808 225004 242860 225010
rect 242808 224946 242860 224952
rect 242268 114510 242296 224946
rect 243544 202156 243596 202162
rect 243544 202098 243596 202104
rect 242256 114504 242308 114510
rect 242256 114446 242308 114452
rect 242164 113824 242216 113830
rect 242164 113766 242216 113772
rect 242164 111104 242216 111110
rect 242164 111046 242216 111052
rect 242176 90370 242204 111046
rect 242164 90364 242216 90370
rect 242164 90306 242216 90312
rect 241520 87644 241572 87650
rect 241520 87586 241572 87592
rect 241532 66230 241560 87586
rect 243556 85474 243584 202098
rect 243648 192506 243676 235214
rect 244924 200796 244976 200802
rect 244924 200738 244976 200744
rect 243636 192500 243688 192506
rect 243636 192442 243688 192448
rect 244936 181490 244964 200738
rect 244924 181484 244976 181490
rect 244924 181426 244976 181432
rect 243636 155304 243688 155310
rect 243636 155246 243688 155252
rect 243648 135930 243676 155246
rect 244924 149116 244976 149122
rect 244924 149058 244976 149064
rect 243636 135924 243688 135930
rect 243636 135866 243688 135872
rect 244280 86284 244332 86290
rect 244280 86226 244332 86232
rect 242808 85468 242860 85474
rect 242808 85410 242860 85416
rect 243544 85468 243596 85474
rect 243544 85410 243596 85416
rect 242820 84250 242848 85410
rect 242808 84244 242860 84250
rect 242808 84186 242860 84192
rect 241520 66224 241572 66230
rect 241520 66166 241572 66172
rect 241532 16574 241560 66166
rect 242820 20058 242848 84186
rect 242808 20052 242860 20058
rect 242808 19994 242860 20000
rect 242992 19984 243044 19990
rect 242992 19926 243044 19932
rect 243004 16574 243032 19926
rect 244292 16574 244320 86226
rect 244936 38010 244964 149058
rect 245120 145586 245148 241604
rect 247052 241590 247526 241618
rect 247052 240145 247080 241590
rect 247038 240136 247094 240145
rect 247038 240071 247094 240080
rect 246302 239456 246358 239465
rect 246302 239391 246358 239400
rect 246316 226273 246344 239391
rect 246302 226264 246358 226273
rect 246302 226199 246358 226208
rect 245568 225684 245620 225690
rect 245568 225626 245620 225632
rect 245580 217938 245608 225626
rect 246316 225049 246344 226199
rect 245658 225040 245714 225049
rect 245658 224975 245714 224984
rect 246302 225040 246358 225049
rect 246302 224975 246358 224984
rect 245568 217932 245620 217938
rect 245568 217874 245620 217880
rect 245580 216714 245608 217874
rect 245568 216708 245620 216714
rect 245568 216650 245620 216656
rect 245108 145580 245160 145586
rect 245108 145522 245160 145528
rect 245016 142860 245068 142866
rect 245016 142802 245068 142808
rect 245028 91798 245056 142802
rect 245672 109002 245700 224975
rect 246304 216708 246356 216714
rect 246304 216650 246356 216656
rect 246316 192506 246344 216650
rect 246304 192500 246356 192506
rect 246304 192442 246356 192448
rect 245660 108996 245712 109002
rect 245660 108938 245712 108944
rect 245660 99476 245712 99482
rect 245660 99418 245712 99424
rect 245672 98666 245700 99418
rect 245660 98660 245712 98666
rect 245660 98602 245712 98608
rect 246316 95849 246344 192442
rect 246302 95840 246358 95849
rect 246302 95775 246358 95784
rect 245016 91792 245068 91798
rect 245016 91734 245068 91740
rect 245660 76560 245712 76566
rect 245660 76502 245712 76508
rect 244924 38004 244976 38010
rect 244924 37946 244976 37952
rect 245672 16574 245700 76502
rect 247052 56506 247080 240071
rect 249064 239420 249116 239426
rect 249064 239362 249116 239368
rect 247682 232656 247738 232665
rect 247682 232591 247738 232600
rect 247696 201482 247724 232591
rect 247684 201476 247736 201482
rect 247684 201418 247736 201424
rect 247132 162172 247184 162178
rect 247132 162114 247184 162120
rect 247144 161430 247172 162114
rect 247132 161424 247184 161430
rect 247132 161366 247184 161372
rect 247682 147928 247738 147937
rect 247682 147863 247738 147872
rect 247696 134570 247724 147863
rect 249076 135250 249104 239362
rect 249156 236020 249208 236026
rect 249156 235962 249208 235968
rect 249168 212498 249196 235962
rect 249904 235890 249932 241604
rect 249892 235884 249944 235890
rect 249892 235826 249944 235832
rect 249156 212492 249208 212498
rect 249156 212434 249208 212440
rect 249800 155236 249852 155242
rect 249800 155178 249852 155184
rect 249064 135244 249116 135250
rect 249064 135186 249116 135192
rect 247684 134564 247736 134570
rect 247684 134506 247736 134512
rect 248420 78668 248472 78674
rect 248420 78610 248472 78616
rect 247040 56500 247092 56506
rect 247040 56442 247092 56448
rect 247592 56500 247644 56506
rect 247592 56442 247644 56448
rect 247604 55894 247632 56442
rect 247592 55888 247644 55894
rect 247592 55830 247644 55836
rect 246304 24132 246356 24138
rect 246304 24074 246356 24080
rect 241532 16546 241744 16574
rect 243004 16546 244136 16574
rect 244292 16546 245240 16574
rect 245672 16546 245976 16574
rect 240784 15904 240836 15910
rect 240784 15846 240836 15852
rect 238024 4412 238076 4418
rect 238024 4354 238076 4360
rect 239312 4412 239364 4418
rect 239312 4354 239364 4360
rect 233884 4072 233936 4078
rect 233884 4014 233936 4020
rect 160744 2100 160796 2106
rect 160744 2042 160796 2048
rect 226984 2100 227036 2106
rect 226984 2042 227036 2048
rect 239324 480 239352 4354
rect 240508 4072 240560 4078
rect 240508 4014 240560 4020
rect 240520 480 240548 4014
rect 241716 480 241744 16546
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242912 480 242940 3402
rect 244108 480 244136 16546
rect 245212 480 245240 16546
rect 245948 490 245976 16546
rect 246316 2990 246344 24074
rect 246304 2984 246356 2990
rect 246304 2926 246356 2932
rect 247592 2984 247644 2990
rect 247592 2926 247644 2932
rect 246224 598 246436 626
rect 246224 490 246252 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 462 246252 490
rect 246408 480 246436 598
rect 247604 480 247632 2926
rect 248432 490 248460 78610
rect 249076 13122 249104 135186
rect 249812 129062 249840 155178
rect 249800 129056 249852 129062
rect 249800 128998 249852 129004
rect 249156 93220 249208 93226
rect 249156 93162 249208 93168
rect 249168 78674 249196 93162
rect 250456 92177 250484 242014
rect 251824 240780 251876 240786
rect 251824 240722 251876 240728
rect 250536 235884 250588 235890
rect 250536 235826 250588 235832
rect 250548 155242 250576 235826
rect 250536 155236 250588 155242
rect 250536 155178 250588 155184
rect 251836 140758 251864 240722
rect 251914 240136 251970 240145
rect 251914 240071 251970 240080
rect 251928 220114 251956 240071
rect 252296 240009 252324 241604
rect 252282 240000 252338 240009
rect 252282 239935 252338 239944
rect 252296 237386 252324 239935
rect 252284 237380 252336 237386
rect 252284 237322 252336 237328
rect 252296 229094 252324 237322
rect 252388 236026 252416 242286
rect 252376 236020 252428 236026
rect 252376 235962 252428 235968
rect 252296 229066 252508 229094
rect 251916 220108 251968 220114
rect 251916 220050 251968 220056
rect 252480 146334 252508 229066
rect 252468 146328 252520 146334
rect 252468 146270 252520 146276
rect 252480 145625 252508 146270
rect 252466 145616 252522 145625
rect 252466 145551 252522 145560
rect 251824 140752 251876 140758
rect 251824 140694 251876 140700
rect 251836 139806 251864 140694
rect 251272 139800 251324 139806
rect 251272 139742 251324 139748
rect 251824 139800 251876 139806
rect 251824 139742 251876 139748
rect 250536 114504 250588 114510
rect 250536 114446 250588 114452
rect 250442 92168 250498 92177
rect 250442 92103 250498 92112
rect 249156 78668 249208 78674
rect 249156 78610 249208 78616
rect 249800 37936 249852 37942
rect 249800 37878 249852 37884
rect 249812 16574 249840 37878
rect 249812 16546 250024 16574
rect 249064 13116 249116 13122
rect 249064 13058 249116 13064
rect 249800 7608 249852 7614
rect 249800 7550 249852 7556
rect 249812 3330 249840 7550
rect 249800 3324 249852 3330
rect 249800 3266 249852 3272
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 250548 7682 250576 114446
rect 251284 16574 251312 139742
rect 252572 92585 252600 307090
rect 253216 306610 253244 342858
rect 253860 327826 253888 363734
rect 253952 347041 253980 440399
rect 254030 415168 254086 415177
rect 254030 415103 254086 415112
rect 254044 389842 254072 415103
rect 254122 412448 254178 412457
rect 254122 412383 254178 412392
rect 254136 390561 254164 412383
rect 254596 407114 254624 449890
rect 254674 446176 254730 446185
rect 254674 446111 254730 446120
rect 254688 431225 254716 446111
rect 255332 439550 255360 463762
rect 255424 447846 255452 469202
rect 256792 459672 256844 459678
rect 256792 459614 256844 459620
rect 255502 454472 255558 454481
rect 255502 454407 255558 454416
rect 255516 449274 255544 454407
rect 256700 451376 256752 451382
rect 256700 451318 256752 451324
rect 255962 450120 256018 450129
rect 255962 450055 256018 450064
rect 255504 449268 255556 449274
rect 255504 449210 255556 449216
rect 255516 448905 255544 449210
rect 255502 448896 255558 448905
rect 255502 448831 255558 448840
rect 255412 447840 255464 447846
rect 255412 447782 255464 447788
rect 255424 447545 255452 447782
rect 255410 447536 255466 447545
rect 255410 447471 255466 447480
rect 255410 444816 255466 444825
rect 255410 444751 255466 444760
rect 255424 444446 255452 444751
rect 255412 444440 255464 444446
rect 255412 444382 255464 444388
rect 255410 443456 255466 443465
rect 255410 443391 255412 443400
rect 255464 443391 255466 443400
rect 255412 443362 255464 443368
rect 255410 442096 255466 442105
rect 255410 442031 255412 442040
rect 255464 442031 255466 442040
rect 255412 442002 255464 442008
rect 255320 439544 255372 439550
rect 255320 439486 255372 439492
rect 255332 439113 255360 439486
rect 255318 439104 255374 439113
rect 255318 439039 255374 439048
rect 255412 438184 255464 438190
rect 255412 438126 255464 438132
rect 255424 437753 255452 438126
rect 255410 437744 255466 437753
rect 255410 437679 255466 437688
rect 255412 436756 255464 436762
rect 255412 436698 255464 436704
rect 255424 436393 255452 436698
rect 255410 436384 255466 436393
rect 255410 436319 255466 436328
rect 255412 435396 255464 435402
rect 255412 435338 255464 435344
rect 255424 435033 255452 435338
rect 255410 435024 255466 435033
rect 255410 434959 255466 434968
rect 255412 434716 255464 434722
rect 255412 434658 255464 434664
rect 255424 433673 255452 434658
rect 255410 433664 255466 433673
rect 255410 433599 255466 433608
rect 255410 432032 255466 432041
rect 255410 431967 255412 431976
rect 255464 431967 255466 431976
rect 255412 431938 255464 431944
rect 254674 431216 254730 431225
rect 254674 431151 254730 431160
rect 255410 430672 255466 430681
rect 255410 430607 255466 430616
rect 255424 428466 255452 430607
rect 255504 429548 255556 429554
rect 255504 429490 255556 429496
rect 255516 429321 255544 429490
rect 255502 429312 255558 429321
rect 255502 429247 255558 429256
rect 255412 428460 255464 428466
rect 255412 428402 255464 428408
rect 255410 427952 255466 427961
rect 255410 427887 255466 427896
rect 255424 427854 255452 427887
rect 255412 427848 255464 427854
rect 255412 427790 255464 427796
rect 255504 427780 255556 427786
rect 255504 427722 255556 427728
rect 255516 426601 255544 427722
rect 255502 426592 255558 426601
rect 255502 426527 255558 426536
rect 255872 425740 255924 425746
rect 255872 425682 255924 425688
rect 255884 425241 255912 425682
rect 255870 425232 255926 425241
rect 255870 425167 255926 425176
rect 255502 423600 255558 423609
rect 255502 423535 255558 423544
rect 255516 422346 255544 423535
rect 255504 422340 255556 422346
rect 255504 422282 255556 422288
rect 255502 422240 255558 422249
rect 255502 422175 255558 422184
rect 255516 420986 255544 422175
rect 255976 421598 256004 450055
rect 255964 421592 256016 421598
rect 255964 421534 256016 421540
rect 255504 420980 255556 420986
rect 255504 420922 255556 420928
rect 255502 420880 255558 420889
rect 255502 420815 255558 420824
rect 255516 419558 255544 420815
rect 255504 419552 255556 419558
rect 255410 419520 255466 419529
rect 255504 419494 255556 419500
rect 255410 419455 255466 419464
rect 255424 418198 255452 419455
rect 255412 418192 255464 418198
rect 255412 418134 255464 418140
rect 255502 418160 255558 418169
rect 255502 418095 255558 418104
rect 255412 416900 255464 416906
rect 255412 416842 255464 416848
rect 255424 416809 255452 416842
rect 255516 416838 255544 418095
rect 255504 416832 255556 416838
rect 255410 416800 255466 416809
rect 255504 416774 255556 416780
rect 255410 416735 255466 416744
rect 255410 413808 255466 413817
rect 255410 413743 255466 413752
rect 255424 413574 255452 413743
rect 255412 413568 255464 413574
rect 255412 413510 255464 413516
rect 255410 411088 255466 411097
rect 255410 411023 255466 411032
rect 255424 409902 255452 411023
rect 255412 409896 255464 409902
rect 255412 409838 255464 409844
rect 255410 409728 255466 409737
rect 255410 409663 255466 409672
rect 255424 408542 255452 409663
rect 255412 408536 255464 408542
rect 255412 408478 255464 408484
rect 255318 408368 255374 408377
rect 255318 408303 255374 408312
rect 254584 407108 254636 407114
rect 254584 407050 254636 407056
rect 254214 405376 254270 405385
rect 254214 405311 254270 405320
rect 254122 390552 254178 390561
rect 254122 390487 254178 390496
rect 254032 389836 254084 389842
rect 254032 389778 254084 389784
rect 254228 389230 254256 405311
rect 255332 398154 255360 408303
rect 255410 407008 255466 407017
rect 255410 406943 255466 406952
rect 255424 406298 255452 406943
rect 255412 406292 255464 406298
rect 255412 406234 255464 406240
rect 255410 401296 255466 401305
rect 255410 401231 255466 401240
rect 255424 400246 255452 401231
rect 255412 400240 255464 400246
rect 255412 400182 255464 400188
rect 255410 399936 255466 399945
rect 255410 399871 255466 399880
rect 255424 399498 255452 399871
rect 255412 399492 255464 399498
rect 255412 399434 255464 399440
rect 255332 398126 255452 398154
rect 255318 396944 255374 396953
rect 255318 396879 255374 396888
rect 254216 389224 254268 389230
rect 254216 389166 254268 389172
rect 255332 383654 255360 396879
rect 255320 383648 255372 383654
rect 255320 383590 255372 383596
rect 255424 370530 255452 398126
rect 255502 395584 255558 395593
rect 255502 395519 255558 395528
rect 255412 370524 255464 370530
rect 255412 370466 255464 370472
rect 254584 367804 254636 367810
rect 254584 367746 254636 367752
rect 254596 367713 254624 367746
rect 254582 367704 254638 367713
rect 254582 367639 254638 367648
rect 253938 347032 253994 347041
rect 253938 346967 253994 346976
rect 253938 330440 253994 330449
rect 253938 330375 253994 330384
rect 253848 327820 253900 327826
rect 253848 327762 253900 327768
rect 253204 306604 253256 306610
rect 253204 306546 253256 306552
rect 253294 305688 253350 305697
rect 253294 305623 253350 305632
rect 253204 304292 253256 304298
rect 253204 304234 253256 304240
rect 253216 301594 253244 304234
rect 252664 301580 253244 301594
rect 252664 301566 253230 301580
rect 252664 111178 252692 301566
rect 252928 301504 252980 301510
rect 252928 301446 252980 301452
rect 252834 300248 252890 300257
rect 252834 300183 252890 300192
rect 252848 299849 252876 300183
rect 252834 299840 252890 299849
rect 252834 299775 252890 299784
rect 252834 292496 252890 292505
rect 252834 292431 252890 292440
rect 252848 277394 252876 292431
rect 252940 292097 252968 301446
rect 253308 298081 253336 305623
rect 253294 298072 253350 298081
rect 253294 298007 253350 298016
rect 253308 296750 253336 298007
rect 253296 296744 253348 296750
rect 253296 296686 253348 296692
rect 253848 293956 253900 293962
rect 253848 293898 253900 293904
rect 253860 292641 253888 293898
rect 253846 292632 253902 292641
rect 253846 292567 253902 292576
rect 252926 292088 252982 292097
rect 252926 292023 252982 292032
rect 253846 291816 253902 291825
rect 253846 291751 253848 291760
rect 253900 291751 253902 291760
rect 253848 291722 253900 291728
rect 252756 277366 252876 277394
rect 252756 232558 252784 277366
rect 253952 246401 253980 330375
rect 254124 302932 254176 302938
rect 254124 302874 254176 302880
rect 254030 301472 254086 301481
rect 254030 301407 254086 301416
rect 254044 295497 254072 301407
rect 254136 298625 254164 302874
rect 254596 301617 254624 367639
rect 255516 363798 255544 395519
rect 255594 392864 255650 392873
rect 255594 392799 255650 392808
rect 255608 380798 255636 392799
rect 255596 380792 255648 380798
rect 255596 380734 255648 380740
rect 255504 363792 255556 363798
rect 255504 363734 255556 363740
rect 254766 328400 254822 328409
rect 254766 328335 254822 328344
rect 254780 327321 254808 328335
rect 254766 327312 254822 327321
rect 254766 327247 254822 327256
rect 254676 316736 254728 316742
rect 254676 316678 254728 316684
rect 254582 301608 254638 301617
rect 254582 301543 254638 301552
rect 254122 298616 254178 298625
rect 254122 298551 254178 298560
rect 254030 295488 254086 295497
rect 254030 295423 254086 295432
rect 254124 253088 254176 253094
rect 254124 253030 254176 253036
rect 254136 252793 254164 253030
rect 254122 252784 254178 252793
rect 254122 252719 254178 252728
rect 253938 246392 253994 246401
rect 253938 246327 253994 246336
rect 253952 246090 253980 246327
rect 253940 246084 253992 246090
rect 253940 246026 253992 246032
rect 252926 245848 252982 245857
rect 252926 245783 252982 245792
rect 252834 245032 252890 245041
rect 252834 244967 252890 244976
rect 252848 244497 252876 244967
rect 252834 244488 252890 244497
rect 252834 244423 252890 244432
rect 252848 242962 252876 244423
rect 252836 242956 252888 242962
rect 252836 242898 252888 242904
rect 252834 242448 252890 242457
rect 252834 242383 252890 242392
rect 252848 242350 252876 242383
rect 252836 242344 252888 242350
rect 252836 242286 252888 242292
rect 252940 238754 252968 245783
rect 254030 245576 254086 245585
rect 254030 245511 254086 245520
rect 253938 242992 253994 243001
rect 253938 242927 253994 242936
rect 253952 240145 253980 242927
rect 253938 240136 253994 240145
rect 253938 240071 253994 240080
rect 252848 238726 252968 238754
rect 252744 232552 252796 232558
rect 252744 232494 252796 232500
rect 252848 222154 252876 238726
rect 252836 222148 252888 222154
rect 252836 222090 252888 222096
rect 252848 219434 252876 222090
rect 252848 219406 253244 219434
rect 253216 172582 253244 219406
rect 254044 217297 254072 245511
rect 254030 217288 254086 217297
rect 254030 217223 254086 217232
rect 254136 211857 254164 252719
rect 254688 251569 254716 316678
rect 254780 313449 254808 327247
rect 254766 313440 254822 313449
rect 254766 313375 254822 313384
rect 255502 313440 255558 313449
rect 255502 313375 255558 313384
rect 255410 301200 255466 301209
rect 255410 301135 255466 301144
rect 255424 300898 255452 301135
rect 255412 300892 255464 300898
rect 255412 300834 255464 300840
rect 255318 300792 255374 300801
rect 255318 300727 255374 300736
rect 255332 299577 255360 300727
rect 255410 299976 255466 299985
rect 255410 299911 255466 299920
rect 255318 299568 255374 299577
rect 255424 299538 255452 299911
rect 255318 299503 255374 299512
rect 255412 299532 255464 299538
rect 255412 299474 255464 299480
rect 255318 298616 255374 298625
rect 255318 298551 255374 298560
rect 255332 292574 255360 298551
rect 255410 298208 255466 298217
rect 255410 298143 255412 298152
rect 255464 298143 255466 298152
rect 255412 298114 255464 298120
rect 255412 297764 255464 297770
rect 255412 297706 255464 297712
rect 255424 297401 255452 297706
rect 255410 297392 255466 297401
rect 255410 297327 255466 297336
rect 255516 296138 255544 313375
rect 255608 300393 255636 380734
rect 255686 376000 255742 376009
rect 255686 375935 255742 375944
rect 255700 374678 255728 375935
rect 255688 374672 255740 374678
rect 255688 374614 255740 374620
rect 256712 316169 256740 451318
rect 256804 425746 256832 459614
rect 258184 442066 258212 480218
rect 258264 467900 258316 467906
rect 258264 467842 258316 467848
rect 258172 442060 258224 442066
rect 258172 442002 258224 442008
rect 258276 438190 258304 467842
rect 259642 465216 259698 465225
rect 259552 465180 259604 465186
rect 259642 465151 259698 465160
rect 259552 465122 259604 465128
rect 258356 459604 258408 459610
rect 258356 459546 258408 459552
rect 258264 438184 258316 438190
rect 258264 438126 258316 438132
rect 256792 425740 256844 425746
rect 256792 425682 256844 425688
rect 258172 413568 258224 413574
rect 258172 413510 258224 413516
rect 256790 404016 256846 404025
rect 256790 403951 256846 403960
rect 256804 374678 256832 403951
rect 256882 394224 256938 394233
rect 256882 394159 256938 394168
rect 256896 393378 256924 394159
rect 256884 393372 256936 393378
rect 256884 393314 256936 393320
rect 256896 386374 256924 393314
rect 256884 386368 256936 386374
rect 256884 386310 256936 386316
rect 258184 384946 258212 413510
rect 258264 399492 258316 399498
rect 258264 399434 258316 399440
rect 258172 384940 258224 384946
rect 258172 384882 258224 384888
rect 258276 377369 258304 399434
rect 258262 377360 258318 377369
rect 258262 377295 258318 377304
rect 256792 374672 256844 374678
rect 256792 374614 256844 374620
rect 256792 328500 256844 328506
rect 256792 328442 256844 328448
rect 256698 316160 256754 316169
rect 256698 316095 256754 316104
rect 255964 308440 256016 308446
rect 255964 308382 256016 308388
rect 255686 307048 255742 307057
rect 255686 306983 255742 306992
rect 255594 300384 255650 300393
rect 255594 300319 255650 300328
rect 255504 296132 255556 296138
rect 255504 296074 255556 296080
rect 255504 295996 255556 296002
rect 255504 295938 255556 295944
rect 255410 295216 255466 295225
rect 255410 295151 255466 295160
rect 255424 294642 255452 295151
rect 255412 294636 255464 294642
rect 255412 294578 255464 294584
rect 255516 294409 255544 295938
rect 255502 294400 255558 294409
rect 255502 294335 255558 294344
rect 255412 294024 255464 294030
rect 255410 293992 255412 294001
rect 255464 293992 255466 294001
rect 255410 293927 255466 293936
rect 255504 293276 255556 293282
rect 255504 293218 255556 293224
rect 255516 293185 255544 293218
rect 255502 293176 255558 293185
rect 255502 293111 255558 293120
rect 255332 292546 255452 292574
rect 255320 281512 255372 281518
rect 255320 281454 255372 281460
rect 255332 280265 255360 281454
rect 255318 280256 255374 280265
rect 255318 280191 255374 280200
rect 255318 279440 255374 279449
rect 255318 279375 255374 279384
rect 255332 278798 255360 279375
rect 255320 278792 255372 278798
rect 255320 278734 255372 278740
rect 255320 277364 255372 277370
rect 255320 277306 255372 277312
rect 255332 276457 255360 277306
rect 255318 276448 255374 276457
rect 255318 276383 255374 276392
rect 255320 276004 255372 276010
rect 255320 275946 255372 275952
rect 255332 275097 255360 275946
rect 255318 275088 255374 275097
rect 255318 275023 255374 275032
rect 255320 274644 255372 274650
rect 255320 274586 255372 274592
rect 255332 273873 255360 274586
rect 255318 273864 255374 273873
rect 255318 273799 255374 273808
rect 255318 273184 255374 273193
rect 255318 273119 255374 273128
rect 255332 272105 255360 273119
rect 255318 272096 255374 272105
rect 255318 272031 255374 272040
rect 255320 270496 255372 270502
rect 255320 270438 255372 270444
rect 255332 269929 255360 270438
rect 255318 269920 255374 269929
rect 255318 269855 255374 269864
rect 255318 266928 255374 266937
rect 255318 266863 255374 266872
rect 255332 266422 255360 266863
rect 255320 266416 255372 266422
rect 255320 266358 255372 266364
rect 255318 264888 255374 264897
rect 255318 264823 255374 264832
rect 255332 263702 255360 264823
rect 255320 263696 255372 263702
rect 255320 263638 255372 263644
rect 254674 251560 254730 251569
rect 254674 251495 254730 251504
rect 254674 249792 254730 249801
rect 254674 249727 254730 249736
rect 254688 248402 254716 249727
rect 254676 248396 254728 248402
rect 254676 248338 254728 248344
rect 254688 244274 254716 248338
rect 255318 244760 255374 244769
rect 255318 244695 255374 244704
rect 254596 244246 254716 244274
rect 254596 227050 254624 244246
rect 255332 243574 255360 244695
rect 255320 243568 255372 243574
rect 255320 243510 255372 243516
rect 255424 232529 255452 292546
rect 255502 282432 255558 282441
rect 255502 282367 255558 282376
rect 255516 282198 255544 282367
rect 255504 282192 255556 282198
rect 255504 282134 255556 282140
rect 255504 281444 255556 281450
rect 255504 281386 255556 281392
rect 255516 281081 255544 281386
rect 255502 281072 255558 281081
rect 255502 281007 255558 281016
rect 255504 280152 255556 280158
rect 255504 280094 255556 280100
rect 255516 279041 255544 280094
rect 255502 279032 255558 279041
rect 255502 278967 255558 278976
rect 255502 278488 255558 278497
rect 255502 278423 255558 278432
rect 255516 278118 255544 278423
rect 255504 278112 255556 278118
rect 255504 278054 255556 278060
rect 255504 277296 255556 277302
rect 255502 277264 255504 277273
rect 255556 277264 255558 277273
rect 255502 277199 255558 277208
rect 255504 275528 255556 275534
rect 255502 275496 255504 275505
rect 255556 275496 255558 275505
rect 255502 275431 255558 275440
rect 255504 274304 255556 274310
rect 255502 274272 255504 274281
rect 255556 274272 255558 274281
rect 255502 274207 255558 274216
rect 255504 272944 255556 272950
rect 255504 272886 255556 272892
rect 255516 272513 255544 272886
rect 255502 272504 255558 272513
rect 255502 272439 255558 272448
rect 255502 271280 255558 271289
rect 255502 271215 255558 271224
rect 255516 270978 255544 271215
rect 255504 270972 255556 270978
rect 255504 270914 255556 270920
rect 255502 270872 255558 270881
rect 255502 270807 255558 270816
rect 255516 270570 255544 270807
rect 255504 270564 255556 270570
rect 255504 270506 255556 270512
rect 255502 270464 255558 270473
rect 255502 270399 255504 270408
rect 255556 270399 255558 270408
rect 255504 270370 255556 270376
rect 255502 267880 255558 267889
rect 255502 267815 255504 267824
rect 255556 267815 255558 267824
rect 255504 267786 255556 267792
rect 255504 266348 255556 266354
rect 255504 266290 255556 266296
rect 255516 266121 255544 266290
rect 255502 266112 255558 266121
rect 255502 266047 255558 266056
rect 255502 265704 255558 265713
rect 255502 265639 255558 265648
rect 255516 264994 255544 265639
rect 255504 264988 255556 264994
rect 255504 264930 255556 264936
rect 255502 263936 255558 263945
rect 255502 263871 255558 263880
rect 255516 263634 255544 263871
rect 255504 263628 255556 263634
rect 255504 263570 255556 263576
rect 255502 243400 255558 243409
rect 255502 243335 255558 243344
rect 255516 242457 255544 243335
rect 255502 242448 255558 242457
rect 255502 242383 255558 242392
rect 255502 242176 255558 242185
rect 255502 242111 255558 242120
rect 255516 241534 255544 242111
rect 255504 241528 255556 241534
rect 255504 241470 255556 241476
rect 255410 232520 255466 232529
rect 255410 232455 255466 232464
rect 255608 229770 255636 300319
rect 255700 299169 255728 306983
rect 255778 299704 255834 299713
rect 255778 299639 255834 299648
rect 255792 299606 255820 299639
rect 255780 299600 255832 299606
rect 255780 299542 255832 299548
rect 255686 299160 255742 299169
rect 255686 299095 255742 299104
rect 255976 297129 256004 308382
rect 256698 301472 256754 301481
rect 256698 301407 256754 301416
rect 255962 297120 256018 297129
rect 255962 297055 256018 297064
rect 255976 296714 256004 297055
rect 255884 296686 256004 296714
rect 255884 296177 255912 296686
rect 256606 296576 256662 296585
rect 256712 296562 256740 301407
rect 256662 296534 256740 296562
rect 256606 296511 256662 296520
rect 255870 296168 255926 296177
rect 255688 296132 255740 296138
rect 255870 296103 255926 296112
rect 255688 296074 255740 296080
rect 255700 293593 255728 296074
rect 255686 293584 255742 293593
rect 255686 293519 255742 293528
rect 256146 292088 256202 292097
rect 256146 292023 256202 292032
rect 256160 291281 256188 292023
rect 256424 291848 256476 291854
rect 256424 291790 256476 291796
rect 256436 291417 256464 291790
rect 256608 291780 256660 291786
rect 256608 291722 256660 291728
rect 256620 291417 256648 291722
rect 256422 291408 256478 291417
rect 256422 291343 256478 291352
rect 256606 291408 256662 291417
rect 256606 291343 256662 291352
rect 256146 291272 256202 291281
rect 256146 291207 256202 291216
rect 256516 291100 256568 291106
rect 256516 291042 256568 291048
rect 256528 290057 256556 291042
rect 256514 290048 256570 290057
rect 256514 289983 256570 289992
rect 255964 288924 256016 288930
rect 255964 288866 256016 288872
rect 255976 288833 256004 288866
rect 255962 288824 256018 288833
rect 255962 288759 256018 288768
rect 256606 288416 256662 288425
rect 255872 288380 255924 288386
rect 256606 288351 256662 288360
rect 255872 288322 255924 288328
rect 255780 288312 255832 288318
rect 255780 288254 255832 288260
rect 255792 287609 255820 288254
rect 255884 288017 255912 288322
rect 255870 288008 255926 288017
rect 255870 287943 255926 287952
rect 255778 287600 255834 287609
rect 255778 287535 255834 287544
rect 256620 287337 256648 288351
rect 256606 287328 256662 287337
rect 256606 287263 256662 287272
rect 256514 286920 256570 286929
rect 256514 286855 256570 286864
rect 256422 286240 256478 286249
rect 256422 286175 256478 286184
rect 256436 285734 256464 286175
rect 256424 285728 256476 285734
rect 256424 285670 256476 285676
rect 256332 284232 256384 284238
rect 256332 284174 256384 284180
rect 256344 283257 256372 284174
rect 256330 283248 256386 283257
rect 256330 283183 256386 283192
rect 256528 280106 256556 286855
rect 256608 286680 256660 286686
rect 256606 286648 256608 286657
rect 256660 286648 256662 286657
rect 256606 286583 256662 286592
rect 256608 285660 256660 285666
rect 256608 285602 256660 285608
rect 256620 285433 256648 285602
rect 256606 285424 256662 285433
rect 256606 285359 256662 285368
rect 256608 284300 256660 284306
rect 256608 284242 256660 284248
rect 256620 284073 256648 284242
rect 256606 284064 256662 284073
rect 256606 283999 256662 284008
rect 256804 282914 256832 328442
rect 256882 324456 256938 324465
rect 256882 324391 256938 324400
rect 256896 291009 256924 324391
rect 258080 322244 258132 322250
rect 258080 322186 258132 322192
rect 257434 316160 257490 316169
rect 257434 316095 257490 316104
rect 257344 316056 257396 316062
rect 257344 315998 257396 316004
rect 257356 298246 257384 315998
rect 257448 302938 257476 316095
rect 257436 302932 257488 302938
rect 257436 302874 257488 302880
rect 257344 298240 257396 298246
rect 257344 298182 257396 298188
rect 256882 291000 256938 291009
rect 256882 290935 256938 290944
rect 258092 288318 258120 322186
rect 258368 319433 258396 459546
rect 259460 458244 259512 458250
rect 259460 458186 259512 458192
rect 259472 443426 259500 458186
rect 259460 443420 259512 443426
rect 259460 443362 259512 443368
rect 258724 442060 258776 442066
rect 258724 442002 258776 442008
rect 258736 396681 258764 442002
rect 258722 396672 258778 396681
rect 258722 396607 258778 396616
rect 258722 328672 258778 328681
rect 258722 328607 258778 328616
rect 258354 319424 258410 319433
rect 258354 319359 258410 319368
rect 258264 306604 258316 306610
rect 258264 306546 258316 306552
rect 258172 298240 258224 298246
rect 258172 298182 258224 298188
rect 258080 288312 258132 288318
rect 258080 288254 258132 288260
rect 258184 283665 258212 298182
rect 258276 294642 258304 306546
rect 258448 302184 258500 302190
rect 258448 302126 258500 302132
rect 258264 294636 258316 294642
rect 258264 294578 258316 294584
rect 258460 293282 258488 302126
rect 258736 300966 258764 328607
rect 259472 323678 259500 443362
rect 259564 429554 259592 465122
rect 259656 435402 259684 465151
rect 262220 463752 262272 463758
rect 262220 463694 262272 463700
rect 260840 462392 260892 462398
rect 260840 462334 260892 462340
rect 259644 435396 259696 435402
rect 259644 435338 259696 435344
rect 259552 429548 259604 429554
rect 259552 429490 259604 429496
rect 260852 427786 260880 462334
rect 261484 455524 261536 455530
rect 261484 455466 261536 455472
rect 260840 427780 260892 427786
rect 260840 427722 260892 427728
rect 260840 419552 260892 419558
rect 260840 419494 260892 419500
rect 259552 407108 259604 407114
rect 259552 407050 259604 407056
rect 259460 323672 259512 323678
rect 259458 323640 259460 323649
rect 259512 323640 259514 323649
rect 259458 323575 259514 323584
rect 258814 321600 258870 321609
rect 258814 321535 258870 321544
rect 258828 302841 258856 321535
rect 259366 319424 259422 319433
rect 259366 319359 259368 319368
rect 259420 319359 259422 319368
rect 259368 319330 259420 319336
rect 259564 309262 259592 407050
rect 259644 406292 259696 406298
rect 259644 406234 259696 406240
rect 259656 371210 259684 406234
rect 260852 380905 260880 419494
rect 260838 380896 260894 380905
rect 260838 380831 260894 380840
rect 259644 371204 259696 371210
rect 259644 371146 259696 371152
rect 260748 371204 260800 371210
rect 260748 371146 260800 371152
rect 260760 370530 260788 371146
rect 260838 370560 260894 370569
rect 260748 370524 260800 370530
rect 260838 370495 260894 370504
rect 260748 370466 260800 370472
rect 259828 326392 259880 326398
rect 259828 326334 259880 326340
rect 259736 324352 259788 324358
rect 259736 324294 259788 324300
rect 259552 309256 259604 309262
rect 259552 309198 259604 309204
rect 258814 302832 258870 302841
rect 258814 302767 258870 302776
rect 258724 300960 258776 300966
rect 258724 300902 258776 300908
rect 259460 300960 259512 300966
rect 259460 300902 259512 300908
rect 259368 299600 259420 299606
rect 259368 299542 259420 299548
rect 259380 298790 259408 299542
rect 259368 298784 259420 298790
rect 259368 298726 259420 298732
rect 259472 297770 259500 300902
rect 259460 297764 259512 297770
rect 259460 297706 259512 297712
rect 258538 294808 258594 294817
rect 258538 294743 258594 294752
rect 258448 293276 258500 293282
rect 258448 293218 258500 293224
rect 258552 293185 258580 294743
rect 258538 293176 258594 293185
rect 258538 293111 258594 293120
rect 258354 289776 258410 289785
rect 258354 289711 258410 289720
rect 258368 285025 258396 289711
rect 259368 288448 259420 288454
rect 259368 288390 259420 288396
rect 258354 285016 258410 285025
rect 258354 284951 258410 284960
rect 258170 283656 258226 283665
rect 258170 283591 258226 283600
rect 259274 283520 259330 283529
rect 259274 283455 259330 283464
rect 256712 282886 256832 282914
rect 256606 282024 256662 282033
rect 256712 282010 256740 282886
rect 256662 281982 256740 282010
rect 256606 281959 256662 281968
rect 259288 281489 259316 283455
rect 259274 281480 259330 281489
rect 259274 281415 259330 281424
rect 256528 280078 256740 280106
rect 255686 279848 255742 279857
rect 255686 279783 255742 279792
rect 255700 278225 255728 279783
rect 255686 278216 255742 278225
rect 255686 278151 255742 278160
rect 256712 277394 256740 280078
rect 258080 278044 258132 278050
rect 258080 277986 258132 277992
rect 256712 277366 257016 277394
rect 256606 269104 256662 269113
rect 256662 269062 256740 269090
rect 256606 269039 256662 269048
rect 256712 267734 256740 269062
rect 256712 267706 256832 267734
rect 256422 263528 256478 263537
rect 256422 263463 256478 263472
rect 256436 262342 256464 263463
rect 256424 262336 256476 262342
rect 256424 262278 256476 262284
rect 256608 261520 256660 261526
rect 256608 261462 256660 261468
rect 256620 261361 256648 261462
rect 256606 261352 256662 261361
rect 256606 261287 256662 261296
rect 256608 260160 256660 260166
rect 256606 260128 256608 260137
rect 256660 260128 256662 260137
rect 256606 260063 256662 260072
rect 255962 259312 256018 259321
rect 255962 259247 256018 259256
rect 255976 258806 256004 259247
rect 256606 258904 256662 258913
rect 256606 258839 256662 258848
rect 255964 258800 256016 258806
rect 255964 258742 256016 258748
rect 256620 258738 256648 258839
rect 256608 258732 256660 258738
rect 256608 258674 256660 258680
rect 256332 258052 256384 258058
rect 256332 257994 256384 258000
rect 256344 257145 256372 257994
rect 256608 257440 256660 257446
rect 256608 257382 256660 257388
rect 256330 257136 256386 257145
rect 256330 257071 256386 257080
rect 256620 256737 256648 257382
rect 256606 256728 256662 256737
rect 256606 256663 256662 256672
rect 256606 256320 256662 256329
rect 256606 256255 256662 256264
rect 256620 256018 256648 256255
rect 256608 256012 256660 256018
rect 256608 255954 256660 255960
rect 256606 255368 256662 255377
rect 256606 255303 256608 255312
rect 256660 255303 256662 255312
rect 256608 255274 256660 255280
rect 256608 254652 256660 254658
rect 256608 254594 256660 254600
rect 256620 254561 256648 254594
rect 256606 254552 256662 254561
rect 256606 254487 256662 254496
rect 255778 253328 255834 253337
rect 255778 253263 255834 253272
rect 255792 252618 255820 253263
rect 255780 252612 255832 252618
rect 255780 252554 255832 252560
rect 256422 252376 256478 252385
rect 256422 252311 256478 252320
rect 256436 251326 256464 252311
rect 256606 251560 256662 251569
rect 256606 251495 256662 251504
rect 256424 251320 256476 251326
rect 256424 251262 256476 251268
rect 256620 251258 256648 251495
rect 256608 251252 256660 251258
rect 256608 251194 256660 251200
rect 256606 250744 256662 250753
rect 256606 250679 256662 250688
rect 256620 250510 256648 250679
rect 256608 250504 256660 250510
rect 256608 250446 256660 250452
rect 256712 250374 256740 250405
rect 256700 250368 256752 250374
rect 256606 250336 256662 250345
rect 256662 250316 256700 250322
rect 256662 250310 256752 250316
rect 256662 250294 256740 250310
rect 256606 250271 256662 250280
rect 256238 249384 256294 249393
rect 256238 249319 256294 249328
rect 256252 248470 256280 249319
rect 256606 248976 256662 248985
rect 256606 248911 256662 248920
rect 256620 248538 256648 248911
rect 256608 248532 256660 248538
rect 256608 248474 256660 248480
rect 256240 248464 256292 248470
rect 256240 248406 256292 248412
rect 256514 247208 256570 247217
rect 256514 247143 256570 247152
rect 256528 246265 256556 247143
rect 256608 247036 256660 247042
rect 256608 246978 256660 246984
rect 256620 246809 256648 246978
rect 256606 246800 256662 246809
rect 256606 246735 256662 246744
rect 256514 246256 256570 246265
rect 256514 246191 256570 246200
rect 255686 244216 255742 244225
rect 255686 244151 255742 244160
rect 255700 242962 255728 244151
rect 255778 243808 255834 243817
rect 255778 243743 255834 243752
rect 255688 242956 255740 242962
rect 255688 242898 255740 242904
rect 255792 241505 255820 243743
rect 255778 241496 255834 241505
rect 255778 241431 255834 241440
rect 256712 240854 256740 250294
rect 256700 240848 256752 240854
rect 256700 240790 256752 240796
rect 256804 234598 256832 267706
rect 256882 263120 256938 263129
rect 256882 263055 256938 263064
rect 256896 240825 256924 263055
rect 256882 240816 256938 240825
rect 256882 240751 256938 240760
rect 256792 234592 256844 234598
rect 256792 234534 256844 234540
rect 255596 229764 255648 229770
rect 255596 229706 255648 229712
rect 254584 227044 254636 227050
rect 254584 226986 254636 226992
rect 255320 222896 255372 222902
rect 255320 222838 255372 222844
rect 255332 221474 255360 222838
rect 255320 221468 255372 221474
rect 255320 221410 255372 221416
rect 256608 217320 256660 217326
rect 256608 217262 256660 217268
rect 254122 211848 254178 211857
rect 254122 211783 254178 211792
rect 253848 211200 253900 211206
rect 253848 211142 253900 211148
rect 253860 209001 253888 211142
rect 253846 208992 253902 209001
rect 253846 208927 253902 208936
rect 254136 200114 254164 211783
rect 255962 204912 256018 204921
rect 255962 204847 256018 204856
rect 253952 200086 254164 200114
rect 253204 172576 253256 172582
rect 253204 172518 253256 172524
rect 253216 166433 253244 172518
rect 253202 166424 253258 166433
rect 253202 166359 253258 166368
rect 252744 117360 252796 117366
rect 252744 117302 252796 117308
rect 252652 111172 252704 111178
rect 252652 111114 252704 111120
rect 252558 92576 252614 92585
rect 252558 92511 252614 92520
rect 252756 82754 252784 117302
rect 253952 89593 253980 200086
rect 255318 175808 255374 175817
rect 255318 175743 255374 175752
rect 255332 175409 255360 175743
rect 255318 175400 255374 175409
rect 255318 175335 255374 175344
rect 253938 89584 253994 89593
rect 253938 89519 253994 89528
rect 252744 82748 252796 82754
rect 252744 82690 252796 82696
rect 252756 81462 252784 82690
rect 252744 81456 252796 81462
rect 252744 81398 252796 81404
rect 253204 81456 253256 81462
rect 253204 81398 253256 81404
rect 251284 16546 252416 16574
rect 250536 7676 250588 7682
rect 250536 7618 250588 7624
rect 251180 3324 251232 3330
rect 251180 3266 251232 3272
rect 251192 480 251220 3266
rect 252388 480 252416 16546
rect 253216 15230 253244 81398
rect 255332 16574 255360 175335
rect 255976 158982 256004 204847
rect 256056 199436 256108 199442
rect 256056 199378 256108 199384
rect 256068 175817 256096 199378
rect 256054 175808 256110 175817
rect 256054 175743 256110 175752
rect 255412 158976 255464 158982
rect 255412 158918 255464 158924
rect 255964 158976 256016 158982
rect 255964 158918 256016 158924
rect 255424 158846 255452 158918
rect 255412 158840 255464 158846
rect 255412 158782 255464 158788
rect 255424 126954 255452 158782
rect 256620 141001 256648 217262
rect 256988 156058 257016 277366
rect 258092 275534 258120 277986
rect 259380 277394 259408 288390
rect 259458 278080 259514 278089
rect 259458 278015 259514 278024
rect 259288 277366 259408 277394
rect 258080 275528 258132 275534
rect 258080 275470 258132 275476
rect 259288 274310 259316 277366
rect 259368 275324 259420 275330
rect 259368 275266 259420 275272
rect 259276 274304 259328 274310
rect 259276 274246 259328 274252
rect 259380 272950 259408 275266
rect 259368 272944 259420 272950
rect 259368 272886 259420 272892
rect 258078 272776 258134 272785
rect 258078 272711 258134 272720
rect 257344 267028 257396 267034
rect 257344 266970 257396 266976
rect 257356 250374 257384 266970
rect 257344 250368 257396 250374
rect 257344 250310 257396 250316
rect 257342 240272 257398 240281
rect 257342 240207 257398 240216
rect 257356 225690 257384 240207
rect 257988 233912 258040 233918
rect 257988 233854 258040 233860
rect 257344 225684 257396 225690
rect 257344 225626 257396 225632
rect 256976 156052 257028 156058
rect 256976 155994 257028 156000
rect 256988 142154 257016 155994
rect 258000 146946 258028 233854
rect 258092 204338 258120 272711
rect 258724 270972 258776 270978
rect 258724 270914 258776 270920
rect 258736 261594 258764 270914
rect 258724 261588 258776 261594
rect 258724 261530 258776 261536
rect 258724 259480 258776 259486
rect 258724 259422 258776 259428
rect 258736 258058 258764 259422
rect 258724 258052 258776 258058
rect 258724 257994 258776 258000
rect 258262 257544 258318 257553
rect 258262 257479 258318 257488
rect 258172 257372 258224 257378
rect 258172 257314 258224 257320
rect 258184 255785 258212 257314
rect 258170 255776 258226 255785
rect 258170 255711 258226 255720
rect 258172 246084 258224 246090
rect 258172 246026 258224 246032
rect 258184 211206 258212 246026
rect 258276 222873 258304 257479
rect 259368 254584 259420 254590
rect 259368 254526 259420 254532
rect 259380 253094 259408 254526
rect 259368 253088 259420 253094
rect 259368 253030 259420 253036
rect 258356 252612 258408 252618
rect 258356 252554 258408 252560
rect 258368 237969 258396 252554
rect 258354 237960 258410 237969
rect 258354 237895 258410 237904
rect 258724 232552 258776 232558
rect 258724 232494 258776 232500
rect 258262 222864 258318 222873
rect 258262 222799 258318 222808
rect 258172 211200 258224 211206
rect 258172 211142 258224 211148
rect 258080 204332 258132 204338
rect 258080 204274 258132 204280
rect 257988 146940 258040 146946
rect 257988 146882 258040 146888
rect 256712 142126 257016 142154
rect 256606 140992 256662 141001
rect 256606 140927 256662 140936
rect 256712 131034 256740 142126
rect 256700 131028 256752 131034
rect 256700 130970 256752 130976
rect 255412 126948 255464 126954
rect 255412 126890 255464 126896
rect 258092 109750 258120 204274
rect 258736 144226 258764 232494
rect 259368 211812 259420 211818
rect 259368 211754 259420 211760
rect 259380 211206 259408 211754
rect 259368 211200 259420 211206
rect 259368 211142 259420 211148
rect 259472 150657 259500 278015
rect 259564 276865 259592 309198
rect 259642 298072 259698 298081
rect 259642 298007 259698 298016
rect 259550 276856 259606 276865
rect 259550 276791 259606 276800
rect 259552 274304 259604 274310
rect 259552 274246 259604 274252
rect 259564 167686 259592 274246
rect 259656 242214 259684 298007
rect 259748 288930 259776 324294
rect 259736 288924 259788 288930
rect 259736 288866 259788 288872
rect 259840 282198 259868 326334
rect 260852 284889 260880 370495
rect 260930 333296 260986 333305
rect 260930 333231 260986 333240
rect 260838 284880 260894 284889
rect 260838 284815 260894 284824
rect 259828 282192 259880 282198
rect 259828 282134 259880 282140
rect 260944 272785 260972 333231
rect 261496 326398 261524 455466
rect 262232 434722 262260 463694
rect 267004 454096 267056 454102
rect 267004 454038 267056 454044
rect 263598 452976 263654 452985
rect 263598 452911 263654 452920
rect 263416 437436 263468 437442
rect 263416 437378 263468 437384
rect 263428 436937 263456 437378
rect 262310 436928 262366 436937
rect 262310 436863 262366 436872
rect 263414 436928 263470 436937
rect 263414 436863 263470 436872
rect 262324 436762 262352 436863
rect 262312 436756 262364 436762
rect 262312 436698 262364 436704
rect 262220 434716 262272 434722
rect 262220 434658 262272 434664
rect 262220 431996 262272 432002
rect 262220 431938 262272 431944
rect 262128 427780 262180 427786
rect 262128 427722 262180 427728
rect 262140 427106 262168 427722
rect 262128 427100 262180 427106
rect 262128 427042 262180 427048
rect 261666 380896 261722 380905
rect 261666 380831 261722 380840
rect 261680 379273 261708 380831
rect 261666 379264 261722 379273
rect 261666 379199 261722 379208
rect 262232 367878 262260 431938
rect 262864 421592 262916 421598
rect 262864 421534 262916 421540
rect 262220 367872 262272 367878
rect 262220 367814 262272 367820
rect 262220 356720 262272 356726
rect 262220 356662 262272 356668
rect 261484 326392 261536 326398
rect 261484 326334 261536 326340
rect 261024 317484 261076 317490
rect 261024 317426 261076 317432
rect 261036 286686 261064 317426
rect 261116 302932 261168 302938
rect 261116 302874 261168 302880
rect 261128 288454 261156 302874
rect 261116 288448 261168 288454
rect 261116 288390 261168 288396
rect 261024 286680 261076 286686
rect 261024 286622 261076 286628
rect 262232 277545 262260 356662
rect 262404 320952 262456 320958
rect 262404 320894 262456 320900
rect 262312 307080 262364 307086
rect 262312 307022 262364 307028
rect 262324 281450 262352 307022
rect 262312 281444 262364 281450
rect 262312 281386 262364 281392
rect 262312 279472 262364 279478
rect 262312 279414 262364 279420
rect 262324 278798 262352 279414
rect 262312 278792 262364 278798
rect 262312 278734 262364 278740
rect 262218 277536 262274 277545
rect 262218 277471 262274 277480
rect 260930 272776 260986 272785
rect 260930 272711 260986 272720
rect 262218 271824 262274 271833
rect 262218 271759 262274 271768
rect 262232 271561 262260 271759
rect 262218 271552 262274 271561
rect 262218 271487 262274 271496
rect 261022 266520 261078 266529
rect 261022 266455 261078 266464
rect 260838 264480 260894 264489
rect 260838 264415 260894 264424
rect 260852 263702 260880 264415
rect 260840 263696 260892 263702
rect 260840 263638 260892 263644
rect 259734 254144 259790 254153
rect 259734 254079 259790 254088
rect 259644 242208 259696 242214
rect 259644 242150 259696 242156
rect 259748 224942 259776 254079
rect 259736 224936 259788 224942
rect 259736 224878 259788 224884
rect 260852 195294 260880 263638
rect 260930 253736 260986 253745
rect 260930 253671 260986 253680
rect 260944 243681 260972 253671
rect 260930 243672 260986 243681
rect 260930 243607 260986 243616
rect 261036 238066 261064 266455
rect 261206 246256 261262 246265
rect 261206 246191 261262 246200
rect 261114 242312 261170 242321
rect 261114 242247 261170 242256
rect 261128 241534 261156 242247
rect 261116 241528 261168 241534
rect 261116 241470 261168 241476
rect 261024 238060 261076 238066
rect 261024 238002 261076 238008
rect 261128 234025 261156 241470
rect 261114 234016 261170 234025
rect 261114 233951 261170 233960
rect 261220 217977 261248 246191
rect 262232 230450 262260 271487
rect 262220 230444 262272 230450
rect 262220 230386 262272 230392
rect 261206 217968 261262 217977
rect 261206 217903 261262 217912
rect 262126 217288 262182 217297
rect 262126 217223 262182 217232
rect 260840 195288 260892 195294
rect 260840 195230 260892 195236
rect 259552 167680 259604 167686
rect 259552 167622 259604 167628
rect 259458 150648 259514 150657
rect 259458 150583 259514 150592
rect 258816 146940 258868 146946
rect 258816 146882 258868 146888
rect 258724 144220 258776 144226
rect 258724 144162 258776 144168
rect 258080 109744 258132 109750
rect 258080 109686 258132 109692
rect 258828 93158 258856 146882
rect 259472 125594 259500 150583
rect 260102 140992 260158 141001
rect 260102 140927 260158 140936
rect 259460 125588 259512 125594
rect 259460 125530 259512 125536
rect 258816 93152 258868 93158
rect 258816 93094 258868 93100
rect 258724 91792 258776 91798
rect 258724 91734 258776 91740
rect 255332 16546 255912 16574
rect 253480 15904 253532 15910
rect 253480 15846 253532 15852
rect 253204 15224 253256 15230
rect 253204 15166 253256 15172
rect 253492 480 253520 15846
rect 254676 6180 254728 6186
rect 254676 6122 254728 6128
rect 254688 480 254716 6122
rect 255884 480 255912 16546
rect 256700 15224 256752 15230
rect 256700 15166 256752 15172
rect 256712 490 256740 15166
rect 258264 8968 258316 8974
rect 258264 8910 258316 8916
rect 256896 598 257108 626
rect 256896 490 256924 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 256712 462 256924 490
rect 257080 480 257108 598
rect 258276 480 258304 8910
rect 258736 7614 258764 91734
rect 259366 87544 259422 87553
rect 259366 87479 259422 87488
rect 259380 86970 259408 87479
rect 259368 86964 259420 86970
rect 259368 86906 259420 86912
rect 259550 83464 259606 83473
rect 259550 83399 259606 83408
rect 258816 38004 258868 38010
rect 258816 37946 258868 37952
rect 258724 7608 258776 7614
rect 258724 7550 258776 7556
rect 258828 3534 258856 37946
rect 259564 6914 259592 83399
rect 259472 6886 259592 6914
rect 258816 3528 258868 3534
rect 258816 3470 258868 3476
rect 259472 480 259500 6886
rect 260116 3466 260144 140927
rect 262140 80102 262168 217223
rect 262232 116686 262260 230386
rect 262324 208350 262352 278734
rect 262416 270434 262444 320894
rect 262876 317665 262904 421534
rect 263612 341562 263640 452911
rect 263784 444440 263836 444446
rect 263784 444382 263836 444388
rect 263692 434716 263744 434722
rect 263692 434658 263744 434664
rect 263704 347857 263732 434658
rect 263796 360874 263824 444382
rect 266360 438184 266412 438190
rect 266360 438126 266412 438132
rect 265256 417512 265308 417518
rect 265256 417454 265308 417460
rect 265268 416906 265296 417454
rect 265072 416900 265124 416906
rect 265072 416842 265124 416848
rect 265256 416900 265308 416906
rect 265256 416842 265308 416848
rect 264980 381540 265032 381546
rect 264980 381482 265032 381488
rect 263784 360868 263836 360874
rect 263784 360810 263836 360816
rect 263690 347848 263746 347857
rect 263690 347783 263746 347792
rect 263600 341556 263652 341562
rect 263600 341498 263652 341504
rect 263600 320884 263652 320890
rect 263600 320826 263652 320832
rect 262862 317656 262918 317665
rect 262862 317591 262918 317600
rect 262496 311976 262548 311982
rect 262496 311918 262548 311924
rect 262508 285734 262536 311918
rect 263506 292496 263562 292505
rect 263506 292431 263562 292440
rect 262496 285728 262548 285734
rect 262496 285670 262548 285676
rect 263520 282985 263548 292431
rect 263612 285666 263640 320826
rect 263704 286929 263732 347783
rect 263874 325000 263930 325009
rect 263874 324935 263930 324944
rect 263784 319388 263836 319394
rect 263784 319330 263836 319336
rect 263690 286920 263746 286929
rect 263690 286855 263746 286864
rect 263600 285660 263652 285666
rect 263600 285602 263652 285608
rect 263506 282976 263562 282985
rect 263506 282911 263562 282920
rect 263692 282192 263744 282198
rect 263692 282134 263744 282140
rect 262404 270428 262456 270434
rect 262404 270370 262456 270376
rect 262680 270428 262732 270434
rect 262680 270370 262732 270376
rect 262692 269142 262720 270370
rect 262680 269136 262732 269142
rect 262680 269078 262732 269084
rect 262404 266416 262456 266422
rect 262404 266358 262456 266364
rect 262416 237289 262444 266358
rect 263232 260160 263284 260166
rect 263230 260128 263232 260137
rect 263284 260128 263286 260137
rect 263230 260063 263286 260072
rect 262496 255332 262548 255338
rect 262496 255274 262548 255280
rect 262402 237280 262458 237289
rect 262402 237215 262458 237224
rect 262508 230489 262536 255274
rect 262494 230480 262550 230489
rect 262494 230415 262550 230424
rect 262312 208344 262364 208350
rect 262312 208286 262364 208292
rect 262220 116680 262272 116686
rect 262220 116622 262272 116628
rect 262324 96626 262352 208286
rect 263704 207058 263732 282134
rect 263796 273601 263824 319330
rect 263888 291106 263916 324935
rect 264992 291854 265020 381482
rect 265084 378049 265112 416842
rect 265070 378040 265126 378049
rect 265070 377975 265126 377984
rect 265256 327820 265308 327826
rect 265256 327762 265308 327768
rect 265072 315308 265124 315314
rect 265072 315250 265124 315256
rect 264980 291848 265032 291854
rect 264980 291790 265032 291796
rect 263876 291100 263928 291106
rect 263876 291042 263928 291048
rect 263968 285728 264020 285734
rect 263968 285670 264020 285676
rect 263782 273592 263838 273601
rect 263782 273527 263838 273536
rect 263782 262848 263838 262857
rect 263782 262783 263838 262792
rect 263796 260953 263824 262783
rect 263874 262712 263930 262721
rect 263874 262647 263930 262656
rect 263782 260944 263838 260953
rect 263782 260879 263838 260888
rect 263692 207052 263744 207058
rect 263692 206994 263744 207000
rect 262312 96620 262364 96626
rect 262312 96562 262364 96568
rect 263704 85542 263732 206994
rect 263796 188358 263824 260879
rect 263888 236609 263916 262647
rect 263874 236600 263930 236609
rect 263874 236535 263930 236544
rect 263784 188352 263836 188358
rect 263784 188294 263836 188300
rect 263980 151094 264008 285670
rect 263968 151088 264020 151094
rect 263968 151030 264020 151036
rect 264992 93226 265020 291790
rect 265084 266354 265112 315250
rect 265164 303680 265216 303686
rect 265164 303622 265216 303628
rect 265072 266348 265124 266354
rect 265072 266290 265124 266296
rect 265070 259448 265126 259457
rect 265070 259383 265126 259392
rect 265084 258806 265112 259383
rect 265072 258800 265124 258806
rect 265072 258742 265124 258748
rect 265072 258664 265124 258670
rect 265072 258606 265124 258612
rect 265084 189786 265112 258606
rect 265176 233918 265204 303622
rect 265268 296002 265296 327762
rect 266372 320249 266400 438126
rect 266452 409896 266504 409902
rect 266452 409838 266504 409844
rect 266464 382265 266492 409838
rect 267016 391270 267044 454038
rect 268384 452804 268436 452810
rect 268384 452746 268436 452752
rect 267740 450016 267792 450022
rect 267740 449958 267792 449964
rect 267004 391264 267056 391270
rect 267004 391206 267056 391212
rect 266544 384328 266596 384334
rect 266544 384270 266596 384276
rect 266450 382256 266506 382265
rect 266450 382191 266506 382200
rect 266358 320240 266414 320249
rect 266358 320175 266414 320184
rect 265256 295996 265308 296002
rect 265256 295938 265308 295944
rect 266372 285977 266400 320175
rect 266358 285968 266414 285977
rect 266358 285903 266414 285912
rect 266358 284472 266414 284481
rect 266358 284407 266414 284416
rect 265254 269784 265310 269793
rect 265254 269719 265310 269728
rect 265268 269385 265296 269719
rect 265254 269376 265310 269385
rect 265254 269311 265310 269320
rect 265268 238649 265296 269311
rect 265806 263392 265862 263401
rect 265806 263327 265862 263336
rect 265820 262342 265848 263327
rect 265348 262336 265400 262342
rect 265348 262278 265400 262284
rect 265808 262336 265860 262342
rect 265808 262278 265860 262284
rect 265360 258670 265388 262278
rect 265348 258664 265400 258670
rect 265348 258606 265400 258612
rect 265254 238640 265310 238649
rect 265254 238575 265310 238584
rect 265164 233912 265216 233918
rect 265164 233854 265216 233860
rect 266372 213246 266400 284407
rect 266464 271833 266492 382191
rect 266556 278118 266584 384270
rect 267752 310622 267780 449958
rect 267832 382968 267884 382974
rect 267832 382910 267884 382916
rect 267740 310616 267792 310622
rect 267740 310558 267792 310564
rect 266636 298172 266688 298178
rect 266636 298114 266688 298120
rect 266648 295225 266676 298114
rect 266634 295216 266690 295225
rect 266634 295151 266690 295160
rect 267002 295216 267058 295225
rect 267002 295151 267058 295160
rect 266636 284844 266688 284850
rect 266636 284786 266688 284792
rect 266648 284481 266676 284786
rect 266634 284472 266690 284481
rect 266634 284407 266690 284416
rect 266544 278112 266596 278118
rect 266544 278054 266596 278060
rect 266450 271824 266506 271833
rect 266450 271759 266506 271768
rect 266452 264988 266504 264994
rect 266452 264930 266504 264936
rect 266464 231810 266492 264930
rect 266452 231804 266504 231810
rect 266452 231746 266504 231752
rect 266360 213240 266412 213246
rect 266360 213182 266412 213188
rect 265072 189780 265124 189786
rect 265072 189722 265124 189728
rect 266372 102134 266400 213182
rect 266556 204950 266584 278054
rect 266728 265668 266780 265674
rect 266728 265610 266780 265616
rect 266740 264994 266768 265610
rect 266728 264988 266780 264994
rect 266728 264930 266780 264936
rect 267016 239426 267044 295151
rect 267752 277302 267780 310558
rect 267844 284850 267872 382910
rect 268396 320890 268424 452746
rect 269120 449200 269172 449206
rect 269120 449142 269172 449148
rect 268384 320884 268436 320890
rect 268384 320826 268436 320832
rect 267922 305008 267978 305017
rect 267922 304943 267978 304952
rect 267832 284844 267884 284850
rect 267832 284786 267884 284792
rect 267740 277296 267792 277302
rect 267740 277238 267792 277244
rect 267832 269068 267884 269074
rect 267832 269010 267884 269016
rect 267844 267850 267872 269010
rect 267832 267844 267884 267850
rect 267832 267786 267884 267792
rect 267740 258052 267792 258058
rect 267740 257994 267792 258000
rect 267752 257446 267780 257994
rect 267740 257440 267792 257446
rect 267738 257408 267740 257417
rect 267792 257408 267794 257417
rect 267738 257343 267794 257352
rect 267004 239420 267056 239426
rect 267004 239362 267056 239368
rect 266544 204944 266596 204950
rect 266544 204886 266596 204892
rect 267004 203652 267056 203658
rect 267004 203594 267056 203600
rect 267016 105602 267044 203594
rect 267844 153105 267872 267786
rect 267936 199442 267964 304943
rect 269132 293962 269160 449142
rect 270592 428460 270644 428466
rect 270592 428402 270644 428408
rect 269212 425740 269264 425746
rect 269212 425682 269264 425688
rect 269224 325694 269252 425682
rect 270408 417444 270460 417450
rect 270408 417386 270460 417392
rect 270420 416838 270448 417386
rect 269304 416832 269356 416838
rect 269304 416774 269356 416780
rect 270408 416832 270460 416838
rect 270408 416774 270460 416780
rect 269316 387569 269344 416774
rect 269302 387560 269358 387569
rect 269302 387495 269358 387504
rect 270500 386436 270552 386442
rect 270500 386378 270552 386384
rect 269224 325666 269344 325694
rect 269316 312225 269344 325666
rect 269396 313948 269448 313954
rect 269396 313890 269448 313896
rect 269302 312216 269358 312225
rect 269302 312151 269358 312160
rect 269120 293956 269172 293962
rect 269120 293898 269172 293904
rect 269210 291272 269266 291281
rect 269210 291207 269266 291216
rect 269118 288416 269174 288425
rect 269118 288351 269174 288360
rect 269132 287337 269160 288351
rect 269118 287328 269174 287337
rect 269118 287263 269174 287272
rect 268014 285696 268070 285705
rect 268014 285631 268070 285640
rect 267924 199436 267976 199442
rect 267924 199378 267976 199384
rect 267830 153096 267886 153105
rect 267830 153031 267886 153040
rect 268028 133890 268056 285631
rect 268290 242448 268346 242457
rect 268290 242383 268346 242392
rect 268304 241466 268332 242383
rect 268292 241460 268344 241466
rect 268292 241402 268344 241408
rect 268304 238754 268332 241402
rect 268304 238726 268424 238754
rect 268396 222193 268424 238726
rect 268382 222184 268438 222193
rect 268382 222119 268438 222128
rect 269132 171086 269160 287263
rect 269224 235278 269252 291207
rect 269316 278089 269344 312151
rect 269408 283529 269436 313890
rect 269394 283520 269450 283529
rect 269394 283455 269450 283464
rect 269302 278080 269358 278089
rect 269302 278015 269358 278024
rect 270512 276010 270540 386378
rect 270604 349858 270632 428402
rect 271156 417518 271184 702918
rect 271236 449268 271288 449274
rect 271236 449210 271288 449216
rect 271144 417512 271196 417518
rect 271144 417454 271196 417460
rect 271248 395350 271276 449210
rect 271880 435396 271932 435402
rect 271880 435338 271932 435344
rect 271236 395344 271288 395350
rect 271236 395286 271288 395292
rect 270592 349852 270644 349858
rect 270592 349794 270644 349800
rect 270592 330540 270644 330546
rect 270592 330482 270644 330488
rect 270604 279478 270632 330482
rect 271892 309194 271920 435338
rect 273352 408536 273404 408542
rect 273352 408478 273404 408484
rect 271972 393372 272024 393378
rect 271972 393314 272024 393320
rect 271880 309188 271932 309194
rect 271880 309130 271932 309136
rect 270774 308408 270830 308417
rect 270774 308343 270830 308352
rect 270684 305040 270736 305046
rect 270684 304982 270736 304988
rect 270592 279472 270644 279478
rect 270592 279414 270644 279420
rect 270500 276004 270552 276010
rect 270500 275946 270552 275952
rect 270498 275224 270554 275233
rect 270498 275159 270554 275168
rect 269304 269136 269356 269142
rect 269304 269078 269356 269084
rect 269212 235272 269264 235278
rect 269212 235214 269264 235220
rect 269210 218104 269266 218113
rect 269210 218039 269266 218048
rect 269120 171080 269172 171086
rect 269120 171022 269172 171028
rect 268016 133884 268068 133890
rect 268016 133826 268068 133832
rect 267832 127696 267884 127702
rect 267832 127638 267884 127644
rect 267004 105596 267056 105602
rect 267004 105538 267056 105544
rect 266360 102128 266412 102134
rect 266360 102070 266412 102076
rect 264980 93220 265032 93226
rect 264980 93162 265032 93168
rect 263692 85536 263744 85542
rect 263692 85478 263744 85484
rect 262128 80096 262180 80102
rect 262128 80038 262180 80044
rect 263600 80096 263652 80102
rect 263600 80038 263652 80044
rect 262218 77888 262274 77897
rect 262218 77823 262274 77832
rect 262232 16574 262260 77823
rect 263612 75886 263640 80038
rect 263600 75880 263652 75886
rect 263600 75822 263652 75828
rect 263612 16574 263640 75822
rect 264980 60036 265032 60042
rect 264980 59978 265032 59984
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 261760 7676 261812 7682
rect 261760 7618 261812 7624
rect 260656 3528 260708 3534
rect 260656 3470 260708 3476
rect 260104 3460 260156 3466
rect 260104 3402 260156 3408
rect 260668 480 260696 3470
rect 261772 480 261800 7618
rect 262508 490 262536 16546
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 264992 490 265020 59978
rect 266544 11756 266596 11762
rect 266544 11698 266596 11704
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 11698
rect 267016 7682 267044 105538
rect 267844 16574 267872 127638
rect 269224 108322 269252 218039
rect 269316 206990 269344 269078
rect 270408 251864 270460 251870
rect 270408 251806 270460 251812
rect 270420 251326 270448 251806
rect 269396 251320 269448 251326
rect 269396 251262 269448 251268
rect 270408 251320 270460 251326
rect 270408 251262 270460 251268
rect 269408 233889 269436 251262
rect 269394 233880 269450 233889
rect 269394 233815 269450 233824
rect 269764 233708 269816 233714
rect 269764 233650 269816 233656
rect 269304 206984 269356 206990
rect 269304 206926 269356 206932
rect 269212 108316 269264 108322
rect 269212 108258 269264 108264
rect 269118 82104 269174 82113
rect 269118 82039 269174 82048
rect 269132 16574 269160 82039
rect 269776 74526 269804 233650
rect 270512 209817 270540 275159
rect 270590 273864 270646 273873
rect 270590 273799 270646 273808
rect 270498 209808 270554 209817
rect 270498 209743 270554 209752
rect 270512 94761 270540 209743
rect 270604 159390 270632 273799
rect 270696 232558 270724 304982
rect 270788 269074 270816 308343
rect 271892 276049 271920 309130
rect 271984 277370 272012 393314
rect 273364 383489 273392 408478
rect 273444 391264 273496 391270
rect 273444 391206 273496 391212
rect 273350 383480 273406 383489
rect 273350 383415 273406 383424
rect 272064 337408 272116 337414
rect 272064 337350 272116 337356
rect 271972 277364 272024 277370
rect 271972 277306 272024 277312
rect 271878 276040 271934 276049
rect 271878 275975 271934 275984
rect 271972 271856 272024 271862
rect 271972 271798 272024 271804
rect 271984 270570 272012 271798
rect 271972 270564 272024 270570
rect 271972 270506 272024 270512
rect 270776 269068 270828 269074
rect 270776 269010 270828 269016
rect 270774 266792 270830 266801
rect 270774 266727 270830 266736
rect 270788 232665 270816 266727
rect 271878 259448 271934 259457
rect 271878 259383 271934 259392
rect 271892 258738 271920 259383
rect 271880 258732 271932 258738
rect 271880 258674 271932 258680
rect 271880 251252 271932 251258
rect 271880 251194 271932 251200
rect 270774 232656 270830 232665
rect 270774 232591 270830 232600
rect 270684 232552 270736 232558
rect 270684 232494 270736 232500
rect 270592 159384 270644 159390
rect 270592 159326 270644 159332
rect 271892 149734 271920 251194
rect 271984 213897 272012 270506
rect 272076 240106 272104 337350
rect 273260 312588 273312 312594
rect 273260 312530 273312 312536
rect 272154 302832 272210 302841
rect 272154 302767 272210 302776
rect 272168 288425 272196 302767
rect 272154 288416 272210 288425
rect 272154 288351 272210 288360
rect 273272 284238 273300 312530
rect 273260 284232 273312 284238
rect 273260 284174 273312 284180
rect 272154 281480 272210 281489
rect 272154 281415 272210 281424
rect 272168 280401 272196 281415
rect 272154 280392 272210 280401
rect 272154 280327 272210 280336
rect 272064 240100 272116 240106
rect 272064 240042 272116 240048
rect 272168 224913 272196 280327
rect 273258 276040 273314 276049
rect 273258 275975 273314 275984
rect 272154 224904 272210 224913
rect 272154 224839 272210 224848
rect 271970 213888 272026 213897
rect 271970 213823 272026 213832
rect 271880 149728 271932 149734
rect 271880 149670 271932 149676
rect 273272 131102 273300 275975
rect 273364 268161 273392 383415
rect 273456 303793 273484 391206
rect 273916 388929 273944 703054
rect 280804 702772 280856 702778
rect 280804 702714 280856 702720
rect 280158 460184 280214 460193
rect 280158 460119 280214 460128
rect 274640 452668 274692 452674
rect 274640 452610 274692 452616
rect 273902 388920 273958 388929
rect 273902 388855 273958 388864
rect 273536 323604 273588 323610
rect 273536 323546 273588 323552
rect 273442 303784 273498 303793
rect 273442 303719 273498 303728
rect 273350 268152 273406 268161
rect 273350 268087 273406 268096
rect 273350 265160 273406 265169
rect 273350 265095 273406 265104
rect 273364 262886 273392 265095
rect 273352 262880 273404 262886
rect 273352 262822 273404 262828
rect 273352 252612 273404 252618
rect 273352 252554 273404 252560
rect 273364 250510 273392 252554
rect 273352 250504 273404 250510
rect 273352 250446 273404 250452
rect 273364 229090 273392 250446
rect 273352 229084 273404 229090
rect 273352 229026 273404 229032
rect 273456 217326 273484 303719
rect 273548 288697 273576 323546
rect 274652 305017 274680 452610
rect 277398 450392 277454 450401
rect 277398 450327 277454 450336
rect 276112 422340 276164 422346
rect 276112 422282 276164 422288
rect 276020 380928 276072 380934
rect 276020 380870 276072 380876
rect 274732 380860 274784 380866
rect 274732 380802 274784 380808
rect 274744 380225 274772 380802
rect 274730 380216 274786 380225
rect 274730 380151 274786 380160
rect 274732 334620 274784 334626
rect 274732 334562 274784 334568
rect 274638 305008 274694 305017
rect 274638 304943 274694 304952
rect 273534 288688 273590 288697
rect 273534 288623 273590 288632
rect 273534 284880 273590 284889
rect 273534 284815 273590 284824
rect 273444 217320 273496 217326
rect 273444 217262 273496 217268
rect 273548 209774 273576 284815
rect 274744 281489 274772 334562
rect 275006 306504 275062 306513
rect 275006 306439 275062 306448
rect 274822 296984 274878 296993
rect 274822 296919 274878 296928
rect 274730 281480 274786 281489
rect 274730 281415 274786 281424
rect 274732 258732 274784 258738
rect 274732 258674 274784 258680
rect 274744 254658 274772 258674
rect 274732 254652 274784 254658
rect 274732 254594 274784 254600
rect 273364 209746 273576 209774
rect 273364 208418 273392 209746
rect 273352 208412 273404 208418
rect 273352 208354 273404 208360
rect 273260 131096 273312 131102
rect 273260 131038 273312 131044
rect 273364 95946 273392 208354
rect 274744 177342 274772 254594
rect 274836 233714 274864 296919
rect 274914 250200 274970 250209
rect 274914 250135 274970 250144
rect 274824 233708 274876 233714
rect 274824 233650 274876 233656
rect 274928 216617 274956 250135
rect 274914 216608 274970 216617
rect 274914 216543 274970 216552
rect 274732 177336 274784 177342
rect 274732 177278 274784 177284
rect 273352 95940 273404 95946
rect 273352 95882 273404 95888
rect 270498 94752 270554 94761
rect 270498 94687 270554 94696
rect 271144 90364 271196 90370
rect 271144 90306 271196 90312
rect 269764 74520 269816 74526
rect 269764 74462 269816 74468
rect 270500 69692 270552 69698
rect 270500 69634 270552 69640
rect 270512 16574 270540 69634
rect 267844 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 267004 7676 267056 7682
rect 267004 7618 267056 7624
rect 267740 3460 267792 3466
rect 267740 3402 267792 3408
rect 267752 480 267780 3402
rect 268396 490 268424 16546
rect 269120 7608 269172 7614
rect 269120 7550 269172 7556
rect 269132 3534 269160 7550
rect 269120 3528 269172 3534
rect 269120 3470 269172 3476
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 16546
rect 270788 490 270816 16546
rect 271156 6186 271184 90306
rect 273258 86184 273314 86193
rect 273258 86119 273314 86128
rect 271144 6180 271196 6186
rect 271144 6122 271196 6128
rect 272432 3528 272484 3534
rect 272432 3470 272484 3476
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3470
rect 273272 490 273300 86119
rect 275020 84114 275048 306439
rect 275284 298852 275336 298858
rect 275284 298794 275336 298800
rect 275296 252618 275324 298794
rect 276032 271862 276060 380870
rect 276124 322930 276152 422282
rect 276112 322924 276164 322930
rect 276112 322866 276164 322872
rect 276124 288386 276152 322866
rect 276204 319456 276256 319462
rect 276204 319398 276256 319404
rect 276112 288380 276164 288386
rect 276112 288322 276164 288328
rect 276216 281761 276244 319398
rect 277412 313313 277440 450327
rect 277492 400240 277544 400246
rect 277492 400182 277544 400188
rect 277504 376038 277532 400182
rect 279424 384328 279476 384334
rect 279424 384270 279476 384276
rect 277492 376032 277544 376038
rect 277492 375974 277544 375980
rect 277398 313304 277454 313313
rect 277398 313239 277454 313248
rect 276294 302288 276350 302297
rect 276294 302223 276350 302232
rect 276202 281752 276258 281761
rect 276202 281687 276258 281696
rect 276020 271856 276072 271862
rect 276020 271798 276072 271804
rect 276020 263628 276072 263634
rect 276020 263570 276072 263576
rect 275284 252612 275336 252618
rect 275284 252554 275336 252560
rect 276032 163538 276060 263570
rect 276308 217297 276336 302223
rect 276756 287088 276808 287094
rect 276756 287030 276808 287036
rect 276388 256012 276440 256018
rect 276388 255954 276440 255960
rect 276400 255377 276428 255954
rect 276386 255368 276442 255377
rect 276386 255303 276442 255312
rect 276388 244248 276440 244254
rect 276388 244190 276440 244196
rect 276400 242962 276428 244190
rect 276388 242956 276440 242962
rect 276388 242898 276440 242904
rect 276664 242956 276716 242962
rect 276664 242898 276716 242904
rect 276294 217288 276350 217297
rect 276294 217223 276350 217232
rect 276020 163532 276072 163538
rect 276020 163474 276072 163480
rect 276018 131744 276074 131753
rect 276018 131679 276074 131688
rect 275008 84108 275060 84114
rect 275008 84050 275060 84056
rect 275020 83502 275048 84050
rect 275008 83496 275060 83502
rect 275008 83438 275060 83444
rect 276032 16574 276060 131679
rect 276676 86970 276704 242898
rect 276768 240786 276796 287030
rect 277412 273193 277440 313239
rect 277398 273184 277454 273193
rect 277398 273119 277454 273128
rect 277504 270502 277532 375974
rect 279436 375329 279464 384270
rect 279422 375320 279478 375329
rect 279422 375255 279478 375264
rect 279436 373994 279464 375255
rect 278976 373966 279464 373994
rect 278872 371884 278924 371890
rect 278872 371826 278924 371832
rect 278780 305108 278832 305114
rect 278780 305050 278832 305056
rect 278044 300892 278096 300898
rect 278044 300834 278096 300840
rect 277584 294024 277636 294030
rect 277584 293966 277636 293972
rect 277492 270496 277544 270502
rect 277492 270438 277544 270444
rect 277398 268152 277454 268161
rect 277398 268087 277454 268096
rect 276940 264240 276992 264246
rect 276940 264182 276992 264188
rect 276952 263634 276980 264182
rect 276940 263628 276992 263634
rect 276940 263570 276992 263576
rect 276756 240780 276808 240786
rect 276756 240722 276808 240728
rect 277412 227730 277440 268087
rect 277490 240272 277546 240281
rect 277490 240207 277546 240216
rect 277400 227724 277452 227730
rect 277400 227666 277452 227672
rect 277412 115258 277440 227666
rect 277400 115252 277452 115258
rect 277400 115194 277452 115200
rect 277400 98660 277452 98666
rect 277400 98602 277452 98608
rect 276664 86964 276716 86970
rect 276664 86906 276716 86912
rect 277412 16574 277440 98602
rect 277504 89690 277532 240207
rect 277596 200802 277624 293966
rect 278056 255882 278084 300834
rect 278686 273184 278742 273193
rect 278686 273119 278742 273128
rect 278700 273018 278728 273119
rect 278688 273012 278740 273018
rect 278688 272954 278740 272960
rect 278044 255876 278096 255882
rect 278044 255818 278096 255824
rect 278044 248532 278096 248538
rect 278044 248474 278096 248480
rect 278056 233238 278084 248474
rect 278044 233232 278096 233238
rect 278044 233174 278096 233180
rect 277584 200796 277636 200802
rect 277584 200738 277636 200744
rect 278792 102814 278820 305050
rect 278884 244254 278912 371826
rect 278976 256018 279004 373966
rect 279056 313336 279108 313342
rect 279056 313278 279108 313284
rect 279068 287094 279096 313278
rect 279056 287088 279108 287094
rect 279056 287030 279108 287036
rect 280172 265674 280200 460119
rect 280252 336048 280304 336054
rect 280252 335990 280304 335996
rect 280264 298858 280292 335990
rect 280816 311137 280844 702714
rect 282840 389065 282868 703326
rect 300136 703050 300164 703520
rect 332520 703254 332548 703520
rect 348804 703390 348832 703520
rect 348792 703384 348844 703390
rect 348792 703326 348844 703332
rect 364996 703322 365024 703520
rect 364984 703316 365036 703322
rect 364984 703258 365036 703264
rect 332508 703248 332560 703254
rect 332508 703190 332560 703196
rect 300124 703044 300176 703050
rect 300124 702986 300176 702992
rect 397472 702846 397500 703520
rect 413664 703186 413692 703520
rect 413652 703180 413704 703186
rect 413652 703122 413704 703128
rect 429856 702914 429884 703520
rect 462332 703118 462360 703520
rect 462320 703112 462372 703118
rect 462320 703054 462372 703060
rect 478524 702982 478552 703520
rect 478512 702976 478564 702982
rect 478512 702918 478564 702924
rect 429844 702908 429896 702914
rect 429844 702850 429896 702856
rect 397460 702840 397512 702846
rect 397460 702782 397512 702788
rect 494808 702506 494836 703520
rect 527192 702658 527220 703520
rect 543476 702778 543504 703520
rect 543464 702772 543516 702778
rect 543464 702714 543516 702720
rect 559668 702710 559696 703520
rect 527100 702642 527220 702658
rect 559656 702704 559708 702710
rect 559656 702646 559708 702652
rect 527088 702636 527220 702642
rect 527140 702630 527220 702636
rect 527088 702578 527140 702584
rect 580908 702568 580960 702574
rect 580908 702510 580960 702516
rect 494796 702500 494848 702506
rect 494796 702442 494848 702448
rect 580920 697241 580948 702510
rect 580906 697232 580962 697241
rect 580906 697167 580962 697176
rect 582470 683904 582526 683913
rect 582470 683839 582526 683848
rect 582378 630864 582434 630873
rect 582378 630799 582434 630808
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 295340 472116 295392 472122
rect 295340 472058 295392 472064
rect 286324 461644 286376 461650
rect 286324 461586 286376 461592
rect 286336 460970 286364 461586
rect 286324 460964 286376 460970
rect 286324 460906 286376 460912
rect 284298 458280 284354 458289
rect 284298 458215 284354 458224
rect 283012 420980 283064 420986
rect 283012 420922 283064 420928
rect 282826 389056 282882 389065
rect 282826 388991 282882 389000
rect 281724 378820 281776 378826
rect 281724 378762 281776 378768
rect 280802 311128 280858 311137
rect 280802 311063 280858 311072
rect 281540 302252 281592 302258
rect 281540 302194 281592 302200
rect 280526 299568 280582 299577
rect 280526 299503 280582 299512
rect 280252 298852 280304 298858
rect 280252 298794 280304 298800
rect 280344 294636 280396 294642
rect 280344 294578 280396 294584
rect 280160 265668 280212 265674
rect 280160 265610 280212 265616
rect 280250 262168 280306 262177
rect 280250 262103 280306 262112
rect 279056 261588 279108 261594
rect 279056 261530 279108 261536
rect 278964 256012 279016 256018
rect 278964 255954 279016 255960
rect 278872 244248 278924 244254
rect 278872 244190 278924 244196
rect 278872 233232 278924 233238
rect 278872 233174 278924 233180
rect 278884 231878 278912 233174
rect 279068 233170 279096 261530
rect 280264 261526 280292 262103
rect 280252 261520 280304 261526
rect 280252 261462 280304 261468
rect 279056 233164 279108 233170
rect 279056 233106 279108 233112
rect 278872 231872 278924 231878
rect 278872 231814 278924 231820
rect 278884 216646 278912 231814
rect 278872 216640 278924 216646
rect 278872 216582 278924 216588
rect 280160 205692 280212 205698
rect 280160 205634 280212 205640
rect 278780 102808 278832 102814
rect 278780 102750 278832 102756
rect 280172 97481 280200 205634
rect 280356 202162 280384 294578
rect 280434 291408 280490 291417
rect 280434 291343 280490 291352
rect 280448 205698 280476 291343
rect 280436 205692 280488 205698
rect 280436 205634 280488 205640
rect 280344 202156 280396 202162
rect 280344 202098 280396 202104
rect 280540 162178 280568 299503
rect 281356 299464 281408 299470
rect 281356 299406 281408 299412
rect 281368 298858 281396 299406
rect 281356 298852 281408 298858
rect 281356 298794 281408 298800
rect 281264 262880 281316 262886
rect 281264 262822 281316 262828
rect 281276 262206 281304 262822
rect 280804 262200 280856 262206
rect 280804 262142 280856 262148
rect 281264 262200 281316 262206
rect 281264 262142 281316 262148
rect 280816 231130 280844 262142
rect 281448 261520 281500 261526
rect 281448 261462 281500 261468
rect 281460 260914 281488 261462
rect 281448 260908 281500 260914
rect 281448 260850 281500 260856
rect 280804 231124 280856 231130
rect 280804 231066 280856 231072
rect 280528 162172 280580 162178
rect 280528 162114 280580 162120
rect 281446 152008 281502 152017
rect 281446 151943 281502 151952
rect 281460 151774 281488 151943
rect 281448 151768 281500 151774
rect 281448 151710 281500 151716
rect 280158 97472 280214 97481
rect 280158 97407 280214 97416
rect 277492 89684 277544 89690
rect 277492 89626 277544 89632
rect 278688 89684 278740 89690
rect 278688 89626 278740 89632
rect 278700 89010 278728 89626
rect 278688 89004 278740 89010
rect 278688 88946 278740 88952
rect 278780 25560 278832 25566
rect 278780 25502 278832 25508
rect 278792 16574 278820 25502
rect 276032 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 276020 7676 276072 7682
rect 276020 7618 276072 7624
rect 274824 4820 274876 4826
rect 274824 4762 274876 4768
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 4762
rect 276032 480 276060 7618
rect 276676 490 276704 16546
rect 276952 598 277164 626
rect 276952 490 276980 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 462 276980 490
rect 277136 480 277164 598
rect 278332 480 278360 16546
rect 279068 490 279096 16546
rect 281460 3534 281488 151710
rect 281552 116618 281580 302194
rect 281630 301744 281686 301753
rect 281630 301679 281686 301688
rect 281644 174554 281672 301679
rect 281736 274650 281764 378762
rect 281816 370524 281868 370530
rect 281816 370466 281868 370472
rect 281828 281518 281856 370466
rect 282920 307828 282972 307834
rect 282920 307770 282972 307776
rect 281816 281512 281868 281518
rect 281816 281454 281868 281460
rect 281724 274644 281776 274650
rect 281724 274586 281776 274592
rect 281724 273012 281776 273018
rect 281724 272954 281776 272960
rect 281632 174548 281684 174554
rect 281632 174490 281684 174496
rect 281736 153785 281764 272954
rect 281722 153776 281778 153785
rect 281722 153711 281778 153720
rect 282184 120760 282236 120766
rect 282184 120702 282236 120708
rect 281540 116612 281592 116618
rect 281540 116554 281592 116560
rect 281540 68332 281592 68338
rect 281540 68274 281592 68280
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 280712 2100 280764 2106
rect 280712 2042 280764 2048
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 2042
rect 281552 490 281580 68274
rect 282196 2990 282224 120702
rect 282932 107642 282960 307770
rect 283024 247042 283052 420922
rect 283104 326392 283156 326398
rect 283104 326334 283156 326340
rect 283116 248713 283144 326334
rect 284312 318753 284340 458215
rect 285680 427100 285732 427106
rect 285680 427042 285732 427048
rect 285692 426494 285720 427042
rect 285680 426488 285732 426494
rect 285680 426430 285732 426436
rect 285692 422294 285720 426430
rect 285692 422266 285812 422294
rect 284392 373312 284444 373318
rect 284392 373254 284444 373260
rect 284298 318744 284354 318753
rect 284298 318679 284354 318688
rect 284298 293176 284354 293185
rect 284298 293111 284354 293120
rect 283102 248704 283158 248713
rect 283102 248639 283158 248648
rect 283116 248414 283144 248639
rect 283116 248386 283604 248414
rect 283012 247036 283064 247042
rect 283012 246978 283064 246984
rect 283576 234666 283604 248386
rect 283564 234660 283616 234666
rect 283564 234602 283616 234608
rect 283576 218822 283604 234602
rect 283564 218816 283616 218822
rect 283564 218758 283616 218764
rect 282920 107636 282972 107642
rect 282920 107578 282972 107584
rect 282932 106962 282960 107578
rect 282920 106956 282972 106962
rect 282920 106898 282972 106904
rect 284312 78577 284340 293111
rect 284404 242185 284432 373254
rect 284574 318744 284630 318753
rect 284574 318679 284630 318688
rect 284588 317529 284616 318679
rect 284574 317520 284630 317529
rect 284574 317455 284630 317464
rect 284484 295996 284536 296002
rect 284484 295938 284536 295944
rect 284390 242176 284446 242185
rect 284390 242111 284446 242120
rect 284404 81297 284432 242111
rect 284496 218006 284524 295938
rect 284588 264246 284616 317455
rect 284576 264240 284628 264246
rect 284576 264182 284628 264188
rect 285680 260160 285732 260166
rect 285680 260102 285732 260108
rect 285692 259593 285720 260102
rect 285678 259584 285734 259593
rect 285678 259519 285734 259528
rect 285692 259486 285720 259519
rect 285680 259480 285732 259486
rect 285680 259422 285732 259428
rect 285680 255876 285732 255882
rect 285680 255818 285732 255824
rect 284484 218000 284536 218006
rect 284484 217942 284536 217948
rect 284496 203658 284524 217942
rect 284484 203652 284536 203658
rect 284484 203594 284536 203600
rect 284390 81288 284446 81297
rect 284390 81223 284446 81232
rect 284298 78568 284354 78577
rect 284298 78503 284354 78512
rect 282184 2984 282236 2990
rect 282184 2926 282236 2932
rect 283104 2984 283156 2990
rect 283104 2926 283156 2932
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 2926
rect 284312 480 284340 78503
rect 285692 62014 285720 255818
rect 285784 253201 285812 422266
rect 285862 309224 285918 309233
rect 285862 309159 285918 309168
rect 285770 253192 285826 253201
rect 285770 253127 285826 253136
rect 285876 144809 285904 309159
rect 286336 267734 286364 460906
rect 291200 458312 291252 458318
rect 291200 458254 291252 458260
rect 287152 456816 287204 456822
rect 287152 456758 287204 456764
rect 287060 447840 287112 447846
rect 287060 447782 287112 447788
rect 286416 320884 286468 320890
rect 286416 320826 286468 320832
rect 286244 267706 286364 267734
rect 286244 257378 286272 267706
rect 286428 258074 286456 320826
rect 286336 258046 286456 258074
rect 286232 257372 286284 257378
rect 286232 257314 286284 257320
rect 286244 256766 286272 257314
rect 286232 256760 286284 256766
rect 286232 256702 286284 256708
rect 286336 256698 286364 258046
rect 286324 256692 286376 256698
rect 286324 256634 286376 256640
rect 286336 248402 286364 256634
rect 286324 248396 286376 248402
rect 286324 248338 286376 248344
rect 287072 247489 287100 447782
rect 287164 258738 287192 456758
rect 288532 439544 288584 439550
rect 288532 439486 288584 439492
rect 288440 427848 288492 427854
rect 288440 427790 288492 427796
rect 287244 395344 287296 395350
rect 287244 395286 287296 395292
rect 287152 258732 287204 258738
rect 287152 258674 287204 258680
rect 287152 256760 287204 256766
rect 287152 256702 287204 256708
rect 287058 247480 287114 247489
rect 287058 247415 287114 247424
rect 287060 243568 287112 243574
rect 287060 243510 287112 243516
rect 287072 211138 287100 243510
rect 287060 211132 287112 211138
rect 287060 211074 287112 211080
rect 285862 144800 285918 144809
rect 285862 144735 285918 144744
rect 286782 144800 286838 144809
rect 286782 144735 286838 144744
rect 286796 144226 286824 144735
rect 286784 144220 286836 144226
rect 286784 144162 286836 144168
rect 287072 88233 287100 211074
rect 287164 193866 287192 256702
rect 287256 237386 287284 395286
rect 287334 389056 287390 389065
rect 287334 388991 287390 389000
rect 287348 262206 287376 388991
rect 287336 262200 287388 262206
rect 287336 262142 287388 262148
rect 287334 247480 287390 247489
rect 287334 247415 287390 247424
rect 287244 237380 287296 237386
rect 287244 237322 287296 237328
rect 287348 222902 287376 247415
rect 288452 235958 288480 427790
rect 288544 260166 288572 439486
rect 289728 418804 289780 418810
rect 289728 418746 289780 418752
rect 289740 418198 289768 418746
rect 288624 418192 288676 418198
rect 288624 418134 288676 418140
rect 289728 418192 289780 418198
rect 289728 418134 289780 418140
rect 288636 387705 288664 418134
rect 288622 387696 288678 387705
rect 288622 387631 288678 387640
rect 288532 260160 288584 260166
rect 288532 260102 288584 260108
rect 288636 258058 288664 387631
rect 289910 385112 289966 385121
rect 289910 385047 289912 385056
rect 289964 385047 289966 385056
rect 289912 385018 289964 385024
rect 289818 307864 289874 307873
rect 289818 307799 289874 307808
rect 288716 299532 288768 299538
rect 288716 299474 288768 299480
rect 288624 258052 288676 258058
rect 288624 257994 288676 258000
rect 288532 247036 288584 247042
rect 288532 246978 288584 246984
rect 288440 235952 288492 235958
rect 288440 235894 288492 235900
rect 287336 222896 287388 222902
rect 287336 222838 287388 222844
rect 287152 193860 287204 193866
rect 287152 193802 287204 193808
rect 287704 140072 287756 140078
rect 287704 140014 287756 140020
rect 287058 88224 287114 88233
rect 287058 88159 287114 88168
rect 285680 62008 285732 62014
rect 285680 61950 285732 61956
rect 286600 62008 286652 62014
rect 286600 61950 286652 61956
rect 286612 61402 286640 61950
rect 286600 61396 286652 61402
rect 286600 61338 286652 61344
rect 286324 53100 286376 53106
rect 286324 53042 286376 53048
rect 284392 20052 284444 20058
rect 284392 19994 284444 20000
rect 284404 16574 284432 19994
rect 284404 16546 284984 16574
rect 284956 490 284984 16546
rect 286336 3369 286364 53042
rect 287060 28280 287112 28286
rect 287060 28222 287112 28228
rect 287072 16574 287100 28222
rect 287072 16546 287376 16574
rect 286600 3528 286652 3534
rect 286600 3470 286652 3476
rect 286322 3360 286378 3369
rect 286322 3295 286378 3304
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 3470
rect 287348 490 287376 16546
rect 287716 3398 287744 140014
rect 288544 124166 288572 246978
rect 288728 171902 288756 299474
rect 288716 171896 288768 171902
rect 288716 171838 288768 171844
rect 289084 140820 289136 140826
rect 289084 140762 289136 140768
rect 288532 124160 288584 124166
rect 288532 124102 288584 124108
rect 288440 44872 288492 44878
rect 288440 44814 288492 44820
rect 288452 16574 288480 44814
rect 288452 16546 289032 16574
rect 287704 3392 287756 3398
rect 287704 3334 287756 3340
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 16546
rect 289096 3262 289124 140762
rect 289832 59362 289860 307799
rect 289924 254590 289952 385018
rect 291212 295225 291240 458254
rect 291292 374672 291344 374678
rect 291292 374614 291344 374620
rect 291198 295216 291254 295225
rect 291198 295151 291254 295160
rect 290004 293276 290056 293282
rect 290004 293218 290056 293224
rect 289912 254584 289964 254590
rect 289912 254526 289964 254532
rect 290016 225622 290044 293218
rect 291304 267714 291332 374614
rect 294052 347812 294104 347818
rect 294052 347754 294104 347760
rect 292580 345092 292632 345098
rect 292580 345034 292632 345040
rect 291384 343732 291436 343738
rect 291384 343674 291436 343680
rect 291396 280158 291424 343674
rect 291474 295352 291530 295361
rect 291474 295287 291530 295296
rect 291384 280152 291436 280158
rect 291384 280094 291436 280100
rect 291292 267708 291344 267714
rect 291292 267650 291344 267656
rect 291304 267034 291332 267650
rect 291292 267028 291344 267034
rect 291292 266970 291344 266976
rect 291292 248464 291344 248470
rect 291292 248406 291344 248412
rect 290004 225616 290056 225622
rect 290004 225558 290056 225564
rect 291304 198694 291332 248406
rect 291292 198688 291344 198694
rect 291292 198630 291344 198636
rect 291488 151774 291516 295287
rect 292592 275330 292620 345034
rect 293960 298784 294012 298790
rect 293960 298726 294012 298732
rect 292580 275324 292632 275330
rect 292580 275266 292632 275272
rect 292578 268560 292634 268569
rect 292578 268495 292634 268504
rect 292592 186318 292620 268495
rect 292580 186312 292632 186318
rect 292580 186254 292632 186260
rect 291476 151768 291528 151774
rect 291476 151710 291528 151716
rect 291842 142488 291898 142497
rect 291842 142423 291898 142432
rect 289820 59356 289872 59362
rect 289820 59298 289872 59304
rect 291856 29646 291884 142423
rect 293972 67590 294000 298726
rect 294064 284306 294092 347754
rect 294052 284300 294104 284306
rect 294052 284242 294104 284248
rect 295352 269793 295380 472058
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 298098 451888 298154 451897
rect 298098 451823 298154 451832
rect 295524 339516 295576 339522
rect 295524 339458 295576 339464
rect 295430 296848 295486 296857
rect 295430 296783 295486 296792
rect 295338 269784 295394 269793
rect 295338 269719 295394 269728
rect 295340 260908 295392 260914
rect 295340 260850 295392 260856
rect 295352 182850 295380 260850
rect 295340 182844 295392 182850
rect 295340 182786 295392 182792
rect 295340 144220 295392 144226
rect 295340 144162 295392 144168
rect 293960 67584 294012 67590
rect 293960 67526 294012 67532
rect 291936 46232 291988 46238
rect 291936 46174 291988 46180
rect 291200 29640 291252 29646
rect 291200 29582 291252 29588
rect 291844 29640 291896 29646
rect 291844 29582 291896 29588
rect 291212 16574 291240 29582
rect 291212 16546 291424 16574
rect 290188 3392 290240 3398
rect 290188 3334 290240 3340
rect 289084 3256 289136 3262
rect 289084 3198 289136 3204
rect 290200 480 290228 3334
rect 291396 480 291424 16546
rect 291948 3534 291976 46174
rect 295352 16574 295380 144162
rect 295444 63510 295472 296783
rect 295536 278050 295564 339458
rect 296720 296744 296772 296750
rect 296720 296686 296772 296692
rect 295524 278044 295576 278050
rect 295524 277986 295576 277992
rect 296732 91050 296760 296686
rect 298112 241466 298140 451823
rect 582392 380866 582420 630799
rect 582484 437442 582512 683839
rect 582654 670712 582710 670721
rect 582654 670647 582710 670656
rect 582562 644056 582618 644065
rect 582562 643991 582618 644000
rect 582472 437436 582524 437442
rect 582472 437378 582524 437384
rect 582470 431624 582526 431633
rect 582470 431559 582526 431568
rect 582380 380860 582432 380866
rect 582380 380802 582432 380808
rect 582484 367062 582512 431559
rect 582576 398041 582604 643991
rect 582668 456113 582696 670647
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582760 585818 582788 617471
rect 582838 591016 582894 591025
rect 582838 590951 582894 590960
rect 582748 585812 582800 585818
rect 582748 585754 582800 585760
rect 582746 577688 582802 577697
rect 582746 577623 582802 577632
rect 582654 456104 582710 456113
rect 582654 456039 582710 456048
rect 582656 426488 582708 426494
rect 582656 426430 582708 426436
rect 582562 398032 582618 398041
rect 582562 397967 582618 397976
rect 582564 385076 582616 385082
rect 582564 385018 582616 385024
rect 582576 378457 582604 385018
rect 582562 378448 582618 378457
rect 582562 378383 582618 378392
rect 582472 367056 582524 367062
rect 582472 366998 582524 367004
rect 582470 365120 582526 365129
rect 582470 365055 582526 365064
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579632 316742 579660 325207
rect 579620 316736 579672 316742
rect 579620 316678 579672 316684
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 580276 267714 580304 272167
rect 580264 267708 580316 267714
rect 580264 267650 580316 267656
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 580920 256698 580948 258839
rect 580908 256692 580960 256698
rect 580908 256634 580960 256640
rect 582484 251870 582512 365055
rect 582668 351937 582696 426430
rect 582760 367810 582788 577623
rect 582852 399498 582880 590951
rect 583022 564360 583078 564369
rect 583022 564295 583078 564304
rect 582930 524512 582986 524521
rect 582930 524447 582986 524456
rect 582840 399492 582892 399498
rect 582840 399434 582892 399440
rect 582944 384334 582972 524447
rect 583036 439550 583064 564295
rect 583114 537840 583170 537849
rect 583114 537775 583170 537784
rect 583024 439544 583076 439550
rect 583024 439486 583076 439492
rect 583128 418810 583156 537775
rect 583298 511320 583354 511329
rect 583298 511255 583354 511264
rect 583206 471472 583262 471481
rect 583206 471407 583262 471416
rect 583116 418804 583168 418810
rect 583116 418746 583168 418752
rect 583022 418296 583078 418305
rect 583022 418231 583078 418240
rect 582932 384328 582984 384334
rect 582932 384270 582984 384276
rect 583036 379409 583064 418231
rect 583220 417450 583248 471407
rect 583312 461650 583340 511255
rect 583300 461644 583352 461650
rect 583300 461586 583352 461592
rect 583300 451308 583352 451314
rect 583300 451250 583352 451256
rect 583208 417444 583260 417450
rect 583208 417386 583260 417392
rect 583312 404977 583340 451250
rect 583298 404968 583354 404977
rect 583298 404903 583354 404912
rect 583022 379400 583078 379409
rect 583022 379335 583078 379344
rect 582748 367804 582800 367810
rect 582748 367746 582800 367752
rect 582654 351928 582710 351937
rect 582654 351863 582710 351872
rect 582654 312080 582710 312089
rect 582654 312015 582710 312024
rect 582562 289912 582618 289921
rect 582562 289847 582618 289856
rect 582472 251864 582524 251870
rect 582472 251806 582524 251812
rect 582380 248464 582432 248470
rect 582380 248406 582432 248412
rect 582392 245585 582420 248406
rect 582378 245576 582434 245585
rect 582378 245511 582434 245520
rect 298100 241460 298152 241466
rect 298100 241402 298152 241408
rect 580264 234660 580316 234666
rect 580264 234602 580316 234608
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 580276 219065 580304 234602
rect 580356 222896 580408 222902
rect 580356 222838 580408 222844
rect 580262 219056 580318 219065
rect 580262 218991 580318 219000
rect 580368 205737 580396 222838
rect 580354 205728 580410 205737
rect 580354 205663 580410 205672
rect 582472 203584 582524 203590
rect 582472 203526 582524 203532
rect 580170 192536 580226 192545
rect 580170 192471 580172 192480
rect 580224 192471 580226 192480
rect 580172 192442 580224 192448
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178702 580212 179143
rect 580172 178696 580224 178702
rect 580172 178638 580224 178644
rect 306380 174548 306432 174554
rect 306380 174490 306432 174496
rect 300124 168428 300176 168434
rect 300124 168370 300176 168376
rect 298744 134564 298796 134570
rect 298744 134506 298796 134512
rect 296720 91044 296772 91050
rect 296720 90986 296772 90992
rect 298098 72448 298154 72457
rect 298098 72383 298154 72392
rect 295432 63504 295484 63510
rect 295432 63446 295484 63452
rect 295352 16546 295656 16574
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 294880 3528 294932 3534
rect 294880 3470 294932 3476
rect 293682 3360 293738 3369
rect 293682 3295 293738 3304
rect 292580 3256 292632 3262
rect 292580 3198 292632 3204
rect 292592 480 292620 3198
rect 293696 480 293724 3295
rect 294892 480 294920 3470
rect 295628 490 295656 16546
rect 297272 6180 297324 6186
rect 297272 6122 297324 6128
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 6122
rect 298112 490 298140 72383
rect 298756 3330 298784 134506
rect 299480 128376 299532 128382
rect 299480 128318 299532 128324
rect 298744 3324 298796 3330
rect 298744 3266 298796 3272
rect 299492 2242 299520 128318
rect 300136 3641 300164 168370
rect 302240 160132 302292 160138
rect 302240 160074 302292 160080
rect 301504 35216 301556 35222
rect 301504 35158 301556 35164
rect 300122 3632 300178 3641
rect 300122 3567 300178 3576
rect 301516 3534 301544 35158
rect 301504 3528 301556 3534
rect 301504 3470 301556 3476
rect 301964 3324 302016 3330
rect 301964 3266 302016 3272
rect 299664 3120 299716 3126
rect 299664 3062 299716 3068
rect 299480 2236 299532 2242
rect 299480 2178 299532 2184
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3062
rect 300768 2236 300820 2242
rect 300768 2178 300820 2184
rect 300780 480 300808 2178
rect 301976 480 302004 3266
rect 302252 3126 302280 160074
rect 304264 135924 304316 135930
rect 304264 135866 304316 135872
rect 302884 13116 302936 13122
rect 302884 13058 302936 13064
rect 302896 3505 302924 13058
rect 303160 3528 303212 3534
rect 302882 3496 302938 3505
rect 303160 3470 303212 3476
rect 302882 3431 302938 3440
rect 302240 3120 302292 3126
rect 302240 3062 302292 3068
rect 303172 480 303200 3470
rect 304276 3466 304304 135866
rect 304356 116612 304408 116618
rect 304356 116554 304408 116560
rect 304368 3806 304396 116554
rect 305644 104168 305696 104174
rect 305644 104110 305696 104116
rect 305656 42090 305684 104110
rect 305736 43444 305788 43450
rect 305736 43386 305788 43392
rect 305644 42084 305696 42090
rect 305644 42026 305696 42032
rect 305748 5574 305776 43386
rect 305736 5568 305788 5574
rect 305736 5510 305788 5516
rect 304356 3800 304408 3806
rect 304356 3742 304408 3748
rect 304354 3632 304410 3641
rect 304354 3567 304410 3576
rect 304264 3460 304316 3466
rect 304264 3402 304316 3408
rect 304368 480 304396 3567
rect 305550 3496 305606 3505
rect 305550 3431 305606 3440
rect 305564 480 305592 3431
rect 306392 490 306420 174490
rect 340144 162172 340196 162178
rect 340144 162114 340196 162120
rect 333980 153264 334032 153270
rect 333980 153206 334032 153212
rect 317418 148336 317474 148345
rect 317418 148271 317474 148280
rect 313278 137320 313334 137329
rect 313278 137255 313334 137264
rect 309784 122120 309836 122126
rect 309784 122062 309836 122068
rect 309048 5568 309100 5574
rect 309048 5510 309100 5516
rect 307944 3800 307996 3806
rect 307944 3742 307996 3748
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3742
rect 309060 480 309088 5510
rect 309796 3058 309824 122062
rect 310520 49020 310572 49026
rect 310520 48962 310572 48968
rect 310532 16574 310560 48962
rect 311900 31068 311952 31074
rect 311900 31010 311952 31016
rect 311912 16574 311940 31010
rect 313292 16574 313320 137255
rect 316040 93152 316092 93158
rect 316040 93094 316092 93100
rect 316052 16574 316080 93094
rect 317432 16574 317460 148271
rect 331864 127628 331916 127634
rect 331864 127570 331916 127576
rect 324320 111852 324372 111858
rect 324320 111794 324372 111800
rect 321652 102808 321704 102814
rect 321652 102750 321704 102756
rect 320824 99408 320876 99414
rect 320824 99350 320876 99356
rect 320180 54528 320232 54534
rect 320180 54470 320232 54476
rect 318798 32464 318854 32473
rect 318798 32399 318854 32408
rect 318812 16574 318840 32399
rect 320192 16574 320220 54470
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 310244 3460 310296 3466
rect 310244 3402 310296 3408
rect 309784 3052 309836 3058
rect 309784 2994 309836 3000
rect 310256 480 310284 3402
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 16546
rect 315028 3052 315080 3058
rect 315028 2994 315080 3000
rect 315040 480 315068 2994
rect 316236 480 316264 16546
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 317340 480 317368 3266
rect 318076 490 318104 16546
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 16546
rect 320468 490 320496 16546
rect 320836 8974 320864 99350
rect 321560 10328 321612 10334
rect 321560 10270 321612 10276
rect 320824 8968 320876 8974
rect 320824 8910 320876 8916
rect 321572 3210 321600 10270
rect 321664 3330 321692 102750
rect 322940 83496 322992 83502
rect 322940 83438 322992 83444
rect 321652 3324 321704 3330
rect 321652 3266 321704 3272
rect 321572 3182 322152 3210
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 3182
rect 322952 490 322980 83438
rect 324332 3534 324360 111794
rect 327722 84824 327778 84833
rect 327722 84759 327778 84768
rect 327080 36576 327132 36582
rect 327080 36518 327132 36524
rect 325700 29640 325752 29646
rect 325700 29582 325752 29588
rect 324412 21412 324464 21418
rect 324412 21354 324464 21360
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 21354
rect 325712 16574 325740 29582
rect 325712 16546 326384 16574
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326356 490 326384 16546
rect 327092 3534 327120 36518
rect 327080 3528 327132 3534
rect 327080 3470 327132 3476
rect 327736 3466 327764 84759
rect 329840 42084 329892 42090
rect 329840 42026 329892 42032
rect 329852 16574 329880 42026
rect 331220 17264 331272 17270
rect 331220 17206 331272 17212
rect 329852 16546 330432 16574
rect 328000 3528 328052 3534
rect 328000 3470 328052 3476
rect 327724 3460 327776 3466
rect 327724 3402 327776 3408
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 3470
rect 329196 3460 329248 3466
rect 329196 3402 329248 3408
rect 329208 480 329236 3402
rect 330404 480 330432 16546
rect 331232 490 331260 17206
rect 331876 4554 331904 127570
rect 332692 8968 332744 8974
rect 332692 8910 332744 8916
rect 331864 4548 331916 4554
rect 331864 4490 331916 4496
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 8910
rect 333992 3482 334020 153206
rect 338120 145580 338172 145586
rect 338120 145522 338172 145528
rect 335360 50380 335412 50386
rect 335360 50322 335412 50328
rect 334072 22772 334124 22778
rect 334072 22714 334124 22720
rect 334084 16574 334112 22714
rect 335372 16574 335400 50322
rect 338132 16574 338160 145522
rect 339500 18624 339552 18630
rect 339500 18566 339552 18572
rect 334084 16546 334664 16574
rect 335372 16546 336320 16574
rect 338132 16546 338712 16574
rect 333900 3454 334020 3482
rect 333900 480 333928 3454
rect 334636 490 334664 16546
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 16546
rect 337476 4548 337528 4554
rect 337476 4490 337528 4496
rect 337488 480 337516 4490
rect 338684 480 338712 16546
rect 339512 490 339540 18566
rect 340156 3534 340184 162114
rect 582380 155984 582432 155990
rect 582380 155926 582432 155932
rect 341524 146328 341576 146334
rect 341524 146270 341576 146276
rect 340972 33788 341024 33794
rect 340972 33730 341024 33736
rect 340144 3528 340196 3534
rect 340144 3470 340196 3476
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 33730
rect 341536 3466 341564 146270
rect 582392 126041 582420 155926
rect 582378 126032 582434 126041
rect 582378 125967 582434 125976
rect 353300 117972 353352 117978
rect 353300 117914 353352 117920
rect 342904 106956 342956 106962
rect 342904 106898 342956 106904
rect 342260 55888 342312 55894
rect 342260 55830 342312 55836
rect 342272 6914 342300 55830
rect 342916 16574 342944 106898
rect 351920 71052 351972 71058
rect 351920 70994 351972 71000
rect 345020 61396 345072 61402
rect 345020 61338 345072 61344
rect 345032 16574 345060 61338
rect 349804 40724 349856 40730
rect 349804 40666 349856 40672
rect 342916 16546 343036 16574
rect 345032 16546 345336 16574
rect 342272 6886 342944 6914
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 341524 3460 341576 3466
rect 341524 3402 341576 3408
rect 342180 480 342208 3470
rect 342916 490 342944 6886
rect 343008 4146 343036 16546
rect 344560 14476 344612 14482
rect 344560 14418 344612 14424
rect 342996 4140 343048 4146
rect 342996 4082 343048 4088
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 14418
rect 345308 490 345336 16546
rect 349816 5574 349844 40666
rect 349804 5568 349856 5574
rect 349804 5510 349856 5516
rect 351644 5568 351696 5574
rect 351644 5510 351696 5516
rect 346952 4140 347004 4146
rect 346952 4082 347004 4088
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 4082
rect 350448 3460 350500 3466
rect 350448 3402 350500 3408
rect 349252 3188 349304 3194
rect 349252 3130 349304 3136
rect 348056 3052 348108 3058
rect 348056 2994 348108 3000
rect 348068 480 348096 2994
rect 349264 480 349292 3130
rect 350460 480 350488 3402
rect 351656 480 351684 5510
rect 351932 3194 351960 70994
rect 351920 3188 351972 3194
rect 351920 3130 351972 3136
rect 353312 3058 353340 117914
rect 582380 89004 582432 89010
rect 582380 88946 582432 88952
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 582392 73001 582420 88946
rect 582378 72992 582434 73001
rect 582378 72927 582434 72936
rect 580172 51740 580224 51746
rect 580172 51682 580224 51688
rect 580184 46345 580212 51682
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 353300 3052 353352 3058
rect 353300 2994 353352 3000
rect 581000 3052 581052 3058
rect 581000 2994 581052 3000
rect 581012 480 581040 2994
rect 582208 480 582236 3470
rect 582484 2938 582512 203526
rect 582576 3058 582604 289847
rect 582668 250481 582696 312015
rect 583114 303920 583170 303929
rect 583114 303855 583170 303864
rect 582654 250472 582710 250481
rect 582654 250407 582710 250416
rect 582656 211812 582708 211818
rect 582656 211754 582708 211760
rect 582668 152697 582696 211754
rect 583024 172576 583076 172582
rect 583024 172518 583076 172524
rect 582930 165880 582986 165889
rect 582930 165815 582986 165824
rect 582748 157412 582800 157418
rect 582748 157354 582800 157360
rect 582654 152688 582710 152697
rect 582654 152623 582710 152632
rect 582654 138680 582710 138689
rect 582654 138615 582710 138624
rect 582668 19825 582696 138615
rect 582760 59673 582788 157354
rect 582838 154592 582894 154601
rect 582838 154527 582894 154536
rect 582852 112849 582880 154527
rect 582944 124166 582972 165815
rect 583036 139369 583064 172518
rect 583022 139360 583078 139369
rect 583022 139295 583078 139304
rect 582932 124160 582984 124166
rect 582932 124102 582984 124108
rect 582838 112840 582894 112849
rect 582838 112775 582894 112784
rect 582838 99512 582894 99521
rect 582838 99447 582894 99456
rect 582852 88233 582880 99447
rect 582838 88224 582894 88233
rect 582838 88159 582894 88168
rect 582838 80744 582894 80753
rect 582838 80679 582894 80688
rect 582746 59664 582802 59673
rect 582746 59599 582802 59608
rect 582654 19816 582710 19825
rect 582654 19751 582710 19760
rect 582852 6633 582880 80679
rect 582930 79384 582986 79393
rect 582930 79319 582986 79328
rect 582944 33153 582972 79319
rect 582930 33144 582986 33153
rect 582930 33079 582986 33088
rect 582838 6624 582894 6633
rect 582838 6559 582894 6568
rect 583128 3534 583156 303855
rect 583116 3528 583168 3534
rect 583116 3470 583168 3476
rect 582564 3052 582616 3058
rect 582564 2994 582616 3000
rect 582484 2910 583432 2938
rect 583404 480 583432 2910
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 3146 579944 3202 580000
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 566888 3478 566944
rect 2778 553852 2834 553888
rect 2778 553832 2780 553852
rect 2780 553832 2832 553852
rect 2832 553832 2834 553852
rect 41326 582528 41382 582584
rect 3514 527856 3570 527912
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3422 501744 3478 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3238 449520 3294 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397432 3478 397488
rect 3514 371320 3570 371376
rect 7654 389272 7710 389328
rect 21362 441496 21418 441552
rect 2778 358436 2780 358456
rect 2780 358436 2832 358456
rect 2832 358436 2834 358456
rect 2778 358400 2834 358436
rect 3330 345344 3386 345400
rect 4066 319232 4122 319288
rect 3422 306176 3478 306232
rect 4066 297336 4122 297392
rect 3514 293120 3570 293176
rect 3514 267144 3570 267200
rect 2778 254088 2834 254144
rect 3422 241068 3424 241088
rect 3424 241068 3476 241088
rect 3476 241068 3478 241088
rect 3422 241032 3478 241068
rect 3422 214956 3424 214976
rect 3424 214956 3476 214976
rect 3476 214956 3478 214976
rect 3422 214920 3478 214956
rect 3238 201864 3294 201920
rect 3422 188844 3424 188864
rect 3424 188844 3476 188864
rect 3476 188844 3478 188864
rect 3422 188808 3478 188844
rect 3422 162832 3478 162888
rect 3146 149776 3202 149832
rect 3146 145696 3202 145752
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 3146 71576 3202 71632
rect 3054 58520 3110 58576
rect 3330 45464 3386 45520
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 5446 221448 5502 221504
rect 6826 203496 6882 203552
rect 13726 332560 13782 332616
rect 11702 288360 11758 288416
rect 10966 156576 11022 156632
rect 41326 417424 41382 417480
rect 31666 335416 31722 335472
rect 22006 329840 22062 329896
rect 17866 307808 17922 307864
rect 14462 241304 14518 241360
rect 15106 236544 15162 236600
rect 20626 218592 20682 218648
rect 25502 322904 25558 322960
rect 23386 311888 23442 311944
rect 24766 186904 24822 186960
rect 30286 310528 30342 310584
rect 26146 299512 26202 299568
rect 28906 235184 28962 235240
rect 35806 334056 35862 334112
rect 34426 331200 34482 331256
rect 32402 312024 32458 312080
rect 34334 251776 34390 251832
rect 33046 217232 33102 217288
rect 37094 44784 37150 44840
rect 38566 325760 38622 325816
rect 39946 233824 40002 233880
rect 41326 313384 41382 313440
rect 43442 301280 43498 301336
rect 45466 298696 45522 298752
rect 48134 377984 48190 378040
rect 47582 340856 47638 340912
rect 46754 90752 46810 90808
rect 48226 339496 48282 339552
rect 50986 442176 51042 442232
rect 50802 379344 50858 379400
rect 49606 266464 49662 266520
rect 51446 388320 51502 388376
rect 52182 311072 52238 311128
rect 52182 285912 52238 285968
rect 50986 284280 51042 284336
rect 52366 311072 52422 311128
rect 52182 138624 52238 138680
rect 51722 136720 51778 136776
rect 53286 139440 53342 139496
rect 54758 270680 54814 270736
rect 54850 265004 54852 265024
rect 54852 265004 54904 265024
rect 54904 265004 54906 265024
rect 54850 264968 54906 265004
rect 55126 382064 55182 382120
rect 55126 226888 55182 226944
rect 54942 160656 54998 160712
rect 53654 139440 53710 139496
rect 56506 239400 56562 239456
rect 57518 238312 57574 238368
rect 58898 430616 58954 430672
rect 57886 399472 57942 399528
rect 59082 385600 59138 385656
rect 57610 138760 57666 138816
rect 61842 534656 61898 534712
rect 61658 429256 61714 429312
rect 60554 283328 60610 283384
rect 60462 258168 60518 258224
rect 59174 143656 59230 143712
rect 60462 233144 60518 233200
rect 61750 414296 61806 414352
rect 65982 579944 66038 580000
rect 61934 436192 61990 436248
rect 61750 290400 61806 290456
rect 61014 260888 61070 260944
rect 65890 567568 65946 567624
rect 65890 538736 65946 538792
rect 67178 578584 67234 578640
rect 66718 573144 66774 573200
rect 66810 571784 66866 571840
rect 66902 570152 66958 570208
rect 66534 568928 66590 568984
rect 66902 564712 66958 564768
rect 66902 563352 66958 563408
rect 66166 561992 66222 562048
rect 66074 544040 66130 544096
rect 63130 289040 63186 289096
rect 61842 196560 61898 196616
rect 63038 252728 63094 252784
rect 66074 439592 66130 439648
rect 66074 430344 66130 430400
rect 65982 425176 66038 425232
rect 65890 399472 65946 399528
rect 65890 398792 65946 398848
rect 65890 373904 65946 373960
rect 65706 273128 65762 273184
rect 64694 252728 64750 252784
rect 63222 139576 63278 139632
rect 61382 79872 61438 79928
rect 64510 151000 64566 151056
rect 65982 287544 66038 287600
rect 65982 286184 66038 286240
rect 66810 560632 66866 560688
rect 66810 559272 66866 559328
rect 66810 557912 66866 557968
rect 66902 553560 66958 553616
rect 66718 549480 66774 549536
rect 66810 546760 66866 546816
rect 66810 545400 66866 545456
rect 66626 541320 66682 541376
rect 66810 433336 66866 433392
rect 67086 428168 67142 428224
rect 66994 427352 67050 427408
rect 66626 424088 66682 424144
rect 66810 423272 66866 423328
rect 67086 422184 67142 422240
rect 66626 421096 66682 421152
rect 66810 420008 66866 420064
rect 66810 418920 66866 418976
rect 67086 418124 67142 418160
rect 67086 418104 67088 418124
rect 67088 418104 67140 418124
rect 67140 418104 67142 418124
rect 66258 415928 66314 415984
rect 66810 414840 66866 414896
rect 66258 414296 66314 414352
rect 66902 414024 66958 414080
rect 66258 412936 66314 412992
rect 66258 411848 66314 411904
rect 66626 410760 66682 410816
rect 66810 408856 66866 408912
rect 66902 407768 66958 407824
rect 66810 406680 66866 406736
rect 66810 404504 66866 404560
rect 66810 403688 66866 403744
rect 67454 577224 67510 577280
rect 67362 555192 67418 555248
rect 67270 552200 67326 552256
rect 67546 575320 67602 575376
rect 71778 596264 71834 596320
rect 74262 581168 74318 581224
rect 75366 581032 75422 581088
rect 80702 582392 80758 582448
rect 83002 582528 83058 582584
rect 85486 583888 85542 583944
rect 71502 580760 71558 580816
rect 72422 580760 72478 580816
rect 79874 580760 79930 580816
rect 88246 582528 88302 582584
rect 92110 583752 92166 583808
rect 88706 580760 88762 580816
rect 92386 580760 92442 580816
rect 67730 575864 67786 575920
rect 67638 566616 67694 566672
rect 95238 574776 95294 574832
rect 94686 563624 94742 563680
rect 67822 556552 67878 556608
rect 68650 548256 68706 548312
rect 68650 543496 68706 543552
rect 68374 543292 68430 543348
rect 70306 539708 70362 539744
rect 70306 539688 70308 539708
rect 70308 539688 70360 539708
rect 70360 539688 70362 539708
rect 67730 479440 67786 479496
rect 67270 427352 67326 427408
rect 67270 426264 67326 426320
rect 67546 432520 67602 432576
rect 67546 426264 67602 426320
rect 67454 418104 67510 418160
rect 67362 405592 67418 405648
rect 67178 402600 67234 402656
rect 67178 401648 67234 401704
rect 66718 401512 66774 401568
rect 66810 399608 66866 399664
rect 67178 397468 67180 397488
rect 67180 397468 67232 397488
rect 67232 397468 67234 397488
rect 67178 397432 67234 397468
rect 67178 395256 67234 395312
rect 66810 392264 66866 392320
rect 67362 387232 67418 387288
rect 67638 417016 67694 417072
rect 67546 400424 67602 400480
rect 69662 466520 69718 466576
rect 69754 445576 69810 445632
rect 70306 445576 70362 445632
rect 68006 434696 68062 434752
rect 67822 396344 67878 396400
rect 67638 393388 67640 393408
rect 67640 393388 67692 393408
rect 67692 393388 67694 393408
rect 67638 393352 67694 393388
rect 66166 287544 66222 287600
rect 66166 287136 66222 287192
rect 66074 273128 66130 273184
rect 66258 282940 66314 282976
rect 66258 282920 66260 282940
rect 66260 282920 66312 282940
rect 66312 282920 66314 282940
rect 67362 279656 67418 279712
rect 66810 278840 66866 278896
rect 66810 278024 66866 278080
rect 66810 276392 66866 276448
rect 66810 275576 66866 275632
rect 66718 274760 66774 274816
rect 66810 273944 66866 274000
rect 66810 272312 66866 272368
rect 66810 270680 66866 270736
rect 66626 269864 66682 269920
rect 66166 269048 66222 269104
rect 66810 268232 66866 268288
rect 66810 266600 66866 266656
rect 66534 264988 66590 265024
rect 66534 264968 66536 264988
rect 66536 264968 66588 264988
rect 66588 264968 66590 264988
rect 66810 264152 66866 264208
rect 67546 289176 67602 289232
rect 67638 282784 67694 282840
rect 67546 282104 67602 282160
rect 67086 263336 67142 263392
rect 67454 263336 67510 263392
rect 66534 262520 66590 262576
rect 66258 260888 66314 260944
rect 66534 260072 66590 260128
rect 66442 257624 66498 257680
rect 66534 256672 66590 256728
rect 66258 255312 66314 255368
rect 66810 255212 66812 255232
rect 66812 255212 66864 255232
rect 66864 255212 66866 255232
rect 66810 255176 66866 255212
rect 66810 254360 66866 254416
rect 66994 253544 67050 253600
rect 66626 251912 66682 251968
rect 64602 88168 64658 88224
rect 65890 130600 65946 130656
rect 66534 251776 66590 251832
rect 66810 250280 66866 250336
rect 66810 248648 66866 248704
rect 66534 247832 66590 247888
rect 66810 245384 66866 245440
rect 66902 243752 66958 243808
rect 66718 242936 66774 242992
rect 66810 242120 66866 242176
rect 67454 246200 67510 246256
rect 67362 238176 67418 238232
rect 66166 140800 66222 140856
rect 65982 122168 66038 122224
rect 65982 108568 66038 108624
rect 64786 94424 64842 94480
rect 65890 84088 65946 84144
rect 66074 102584 66130 102640
rect 65982 77016 66038 77072
rect 66902 131960 66958 132016
rect 66350 131144 66406 131200
rect 66902 127608 66958 127664
rect 66810 126792 66866 126848
rect 66718 125976 66774 126032
rect 66258 123800 66314 123856
rect 66626 122984 66682 123040
rect 66810 121372 66866 121408
rect 66810 121352 66812 121372
rect 66812 121352 66864 121372
rect 66864 121352 66866 121372
rect 66902 120536 66958 120592
rect 66810 120012 66866 120048
rect 66810 119992 66812 120012
rect 66812 119992 66864 120012
rect 66864 119992 66866 120012
rect 66902 119176 66958 119232
rect 66718 117544 66774 117600
rect 66810 117000 66866 117056
rect 66258 116184 66314 116240
rect 66902 115368 66958 115424
rect 66810 114552 66866 114608
rect 66810 113736 66866 113792
rect 66902 113192 66958 113248
rect 66810 111560 66866 111616
rect 66810 110744 66866 110800
rect 66810 110200 66866 110256
rect 66810 107752 66866 107808
rect 66810 106936 66866 106992
rect 66534 105596 66590 105632
rect 66534 105576 66536 105596
rect 66536 105576 66588 105596
rect 66588 105576 66590 105596
rect 66810 104796 66812 104816
rect 66812 104796 66864 104816
rect 66864 104796 66866 104816
rect 66810 104760 66866 104796
rect 67362 103944 67418 104000
rect 66810 103128 66866 103184
rect 66626 101768 66682 101824
rect 67362 100136 67418 100192
rect 66810 99592 66866 99648
rect 66810 98776 66866 98832
rect 66442 96328 66498 96384
rect 66810 94968 66866 95024
rect 66994 93336 67050 93392
rect 62026 72392 62082 72448
rect 67638 277208 67694 277264
rect 67914 395256 67970 395312
rect 67914 372544 67970 372600
rect 67822 371184 67878 371240
rect 71042 453056 71098 453112
rect 69202 434288 69258 434344
rect 71226 434832 71282 434888
rect 71226 434560 71282 434616
rect 71870 436056 71926 436112
rect 72698 436056 72754 436112
rect 72606 435240 72662 435296
rect 75918 459584 75974 459640
rect 76746 539552 76802 539608
rect 76562 458768 76618 458824
rect 73802 434696 73858 434752
rect 74170 434696 74226 434752
rect 75826 435376 75882 435432
rect 76378 434288 76434 434344
rect 81438 472504 81494 472560
rect 77390 454008 77446 454064
rect 77114 433744 77170 433800
rect 80978 436192 81034 436248
rect 80334 436056 80390 436112
rect 81346 436056 81402 436112
rect 81898 434288 81954 434344
rect 82818 439592 82874 439648
rect 83094 436056 83150 436112
rect 83094 434288 83150 434344
rect 83830 434016 83886 434072
rect 84658 434288 84714 434344
rect 86222 449928 86278 449984
rect 88430 534792 88486 534848
rect 90362 536696 90418 536752
rect 88338 461488 88394 461544
rect 90914 476720 90970 476776
rect 86958 446392 87014 446448
rect 88522 449928 88578 449984
rect 85854 434288 85910 434344
rect 94318 539688 94374 539744
rect 93950 538872 94006 538928
rect 94686 520920 94742 520976
rect 95330 567160 95386 567216
rect 97170 578856 97226 578912
rect 96710 565800 96766 565856
rect 96802 562264 96858 562320
rect 96802 560904 96858 560960
rect 96986 573416 97042 573472
rect 101402 583888 101458 583944
rect 97906 577496 97962 577552
rect 97906 576716 97908 576736
rect 97908 576716 97960 576736
rect 97960 576716 97962 576736
rect 97906 576680 97962 576716
rect 97538 572056 97594 572112
rect 97906 570016 97962 570072
rect 97262 569200 97318 569256
rect 97078 559544 97134 559600
rect 96894 558728 96950 558784
rect 97906 558728 97962 558784
rect 96618 556824 96674 556880
rect 95422 552472 95478 552528
rect 96710 555464 96766 555520
rect 96894 554104 96950 554160
rect 96986 552744 97042 552800
rect 97078 552472 97134 552528
rect 96710 545672 96766 545728
rect 96618 541592 96674 541648
rect 95330 523640 95386 523696
rect 96710 468424 96766 468480
rect 95330 442176 95386 442232
rect 97446 549364 97502 549400
rect 97446 549344 97448 549364
rect 97448 549344 97500 549364
rect 97500 549344 97502 549364
rect 97078 544312 97134 544368
rect 97078 542952 97134 543008
rect 95606 436736 95662 436792
rect 96894 436056 96950 436112
rect 96250 434288 96306 434344
rect 99378 569200 99434 569256
rect 104162 582528 104218 582584
rect 100758 448568 100814 448624
rect 100022 442176 100078 442232
rect 98642 438096 98698 438152
rect 101218 436192 101274 436248
rect 100390 434288 100446 434344
rect 92846 434152 92902 434208
rect 85854 434016 85910 434072
rect 104254 441496 104310 441552
rect 104898 434560 104954 434616
rect 106922 437280 106978 437336
rect 109682 463528 109738 463584
rect 110326 463528 110382 463584
rect 110326 462304 110382 462360
rect 110326 442312 110382 442368
rect 119342 583752 119398 583808
rect 110786 437008 110842 437064
rect 97722 433880 97778 433936
rect 101126 433880 101182 433936
rect 105358 433880 105414 433936
rect 110142 433880 110198 433936
rect 75458 433608 75514 433664
rect 77482 433608 77538 433664
rect 87234 433608 87290 433664
rect 87970 433608 88026 433664
rect 89626 433608 89682 433664
rect 90086 433608 90142 433664
rect 91282 433608 91338 433664
rect 91558 433608 91614 433664
rect 92938 433608 92994 433664
rect 97722 433608 97778 433664
rect 98366 433608 98422 433664
rect 99194 433608 99250 433664
rect 100666 433608 100722 433664
rect 101126 433608 101182 433664
rect 105358 433608 105414 433664
rect 106738 433608 106794 433664
rect 109038 433608 109094 433664
rect 110142 433608 110198 433664
rect 68650 433064 68706 433120
rect 68374 431840 68430 431896
rect 112718 429800 112774 429856
rect 112718 418376 112774 418432
rect 70398 390904 70454 390960
rect 71686 390904 71742 390960
rect 73986 390904 74042 390960
rect 69110 390088 69166 390144
rect 69110 389136 69166 389192
rect 70076 390088 70132 390144
rect 68834 303592 68890 303648
rect 68006 282920 68062 282976
rect 68558 275984 68614 276040
rect 68190 258712 68246 258768
rect 67822 249464 67878 249520
rect 69294 316104 69350 316160
rect 69202 284280 69258 284336
rect 69110 283192 69166 283248
rect 72422 389000 72478 389056
rect 73066 389000 73122 389056
rect 73066 383560 73122 383616
rect 72514 380840 72570 380896
rect 111982 390904 112038 390960
rect 91282 390768 91338 390824
rect 74446 388728 74502 388784
rect 72422 373224 72478 373280
rect 70858 285776 70914 285832
rect 70398 285640 70454 285696
rect 70306 284824 70362 284880
rect 69294 283464 69350 283520
rect 75826 386144 75882 386200
rect 78586 389408 78642 389464
rect 79138 389000 79194 389056
rect 77206 386280 77262 386336
rect 75182 317328 75238 317384
rect 71962 283600 72018 283656
rect 72422 282920 72478 282976
rect 73802 286184 73858 286240
rect 73710 285640 73766 285696
rect 74906 285912 74962 285968
rect 75182 285912 75238 285968
rect 75918 320048 75974 320104
rect 77298 292712 77354 292768
rect 76010 292576 76066 292632
rect 79874 389000 79930 389056
rect 80058 389000 80114 389056
rect 79322 386960 79378 387016
rect 78586 322768 78642 322824
rect 79966 388320 80022 388376
rect 79874 382200 79930 382256
rect 79966 318008 80022 318064
rect 107934 390632 107990 390688
rect 80978 389000 81034 389056
rect 80426 385600 80482 385656
rect 83002 388320 83058 388376
rect 81346 309848 81402 309904
rect 81806 297472 81862 297528
rect 79322 285640 79378 285696
rect 72698 283056 72754 283112
rect 73710 283056 73766 283112
rect 81530 286048 81586 286104
rect 80978 285912 81034 285968
rect 83462 384240 83518 384296
rect 82910 313248 82966 313304
rect 83094 291760 83150 291816
rect 82082 286048 82138 286104
rect 83186 286048 83242 286104
rect 85026 378664 85082 378720
rect 86866 387368 86922 387424
rect 84106 293256 84162 293312
rect 84106 286048 84162 286104
rect 86866 319368 86922 319424
rect 86774 309712 86830 309768
rect 86682 283736 86738 283792
rect 88982 382880 89038 382936
rect 89626 385600 89682 385656
rect 88154 318008 88210 318064
rect 87050 317328 87106 317384
rect 88430 304136 88486 304192
rect 89534 293120 89590 293176
rect 89534 283464 89590 283520
rect 91098 387776 91154 387832
rect 91006 383696 91062 383752
rect 89718 289720 89774 289776
rect 90270 286048 90326 286104
rect 90086 283464 90142 283520
rect 90822 285640 90878 285696
rect 91006 286048 91062 286104
rect 96986 390496 97042 390552
rect 93766 329024 93822 329080
rect 91282 291080 91338 291136
rect 95146 319368 95202 319424
rect 94502 316104 94558 316160
rect 93858 285640 93914 285696
rect 93858 284960 93914 285016
rect 94042 283464 94098 283520
rect 97446 389000 97502 389056
rect 96894 388864 96950 388920
rect 97906 389000 97962 389056
rect 99654 390360 99710 390416
rect 101034 390496 101090 390552
rect 98918 387504 98974 387560
rect 100850 385736 100906 385792
rect 96526 309712 96582 309768
rect 95238 288496 95294 288552
rect 97262 324944 97318 325000
rect 96618 289856 96674 289912
rect 96434 285640 96490 285696
rect 97262 287680 97318 287736
rect 97262 286320 97318 286376
rect 83462 283192 83518 283248
rect 88154 283192 88210 283248
rect 92386 283192 92442 283248
rect 73526 282920 73582 282976
rect 97906 282920 97962 282976
rect 100022 297472 100078 297528
rect 98734 284824 98790 284880
rect 68834 281152 68890 281208
rect 70950 241712 71006 241768
rect 83830 241712 83886 241768
rect 86590 241712 86646 241768
rect 90362 241712 90418 241768
rect 91558 241712 91614 241768
rect 68926 241440 68982 241496
rect 68650 240760 68706 240816
rect 68558 240080 68614 240136
rect 67546 129784 67602 129840
rect 67546 128832 67602 128888
rect 67546 125160 67602 125216
rect 67546 109384 67602 109440
rect 67454 97144 67510 97200
rect 67454 91976 67510 92032
rect 71410 240080 71466 240136
rect 71870 240080 71926 240136
rect 70306 239128 70362 239184
rect 68926 231104 68982 231160
rect 67730 165552 67786 165608
rect 67730 164328 67786 164384
rect 67822 137944 67878 138000
rect 67730 132776 67786 132832
rect 67730 128968 67786 129024
rect 70306 215192 70362 215248
rect 69662 214784 69718 214840
rect 70306 214784 70362 214840
rect 69294 140800 69350 140856
rect 69846 137400 69902 137456
rect 70490 153040 70546 153096
rect 70306 134952 70362 135008
rect 71778 146920 71834 146976
rect 70582 143384 70638 143440
rect 71134 140800 71190 140856
rect 72238 239944 72294 240000
rect 72974 240080 73030 240136
rect 72882 239400 72938 239456
rect 72790 239264 72846 239320
rect 73526 239808 73582 239864
rect 74354 240080 74410 240136
rect 72330 138624 72386 138680
rect 73342 147736 73398 147792
rect 75918 238448 75974 238504
rect 76562 239128 76618 239184
rect 74814 220088 74870 220144
rect 74538 162016 74594 162072
rect 74814 145560 74870 145616
rect 75918 140936 75974 140992
rect 75366 136720 75422 136776
rect 76102 137944 76158 138000
rect 77942 240760 77998 240816
rect 77574 238312 77630 238368
rect 82266 239944 82322 240000
rect 78678 175208 78734 175264
rect 79322 175208 79378 175264
rect 78126 138624 78182 138680
rect 78862 167592 78918 167648
rect 79966 157392 80022 157448
rect 79322 137264 79378 137320
rect 80242 151816 80298 151872
rect 81438 153720 81494 153776
rect 80702 137400 80758 137456
rect 84106 238720 84162 238776
rect 85854 241576 85910 241632
rect 86866 239400 86922 239456
rect 84290 234504 84346 234560
rect 86866 226344 86922 226400
rect 86222 171128 86278 171184
rect 83462 168952 83518 169008
rect 83002 143520 83058 143576
rect 83462 142432 83518 142488
rect 83002 138760 83058 138816
rect 84658 138760 84714 138816
rect 84750 137944 84806 138000
rect 86314 168408 86370 168464
rect 87602 239808 87658 239864
rect 88246 220904 88302 220960
rect 90914 240080 90970 240136
rect 90822 227024 90878 227080
rect 89074 175344 89130 175400
rect 88338 154536 88394 154592
rect 92340 241440 92396 241496
rect 93122 241304 93178 241360
rect 93444 241304 93500 241360
rect 92478 232464 92534 232520
rect 91006 167728 91062 167784
rect 89718 136720 89774 136776
rect 92662 166232 92718 166288
rect 89994 139576 90050 139632
rect 89994 136584 90050 136640
rect 91098 140800 91154 140856
rect 91098 137808 91154 137864
rect 92570 136720 92626 136776
rect 93674 140800 93730 140856
rect 93950 237360 94006 237416
rect 94134 236680 94190 236736
rect 94226 139984 94282 140040
rect 67914 128152 67970 128208
rect 67822 112376 67878 112432
rect 67822 100952 67878 101008
rect 67914 93880 67970 93936
rect 69708 92656 69764 92712
rect 71180 92656 71236 92712
rect 68282 81232 68338 81288
rect 71778 91024 71834 91080
rect 70306 82048 70362 82104
rect 71778 86808 71834 86864
rect 73342 92384 73398 92440
rect 74262 90752 74318 90808
rect 76286 90888 76342 90944
rect 78034 89528 78090 89584
rect 78402 85312 78458 85368
rect 80978 87896 81034 87952
rect 77298 81096 77354 81152
rect 83002 89664 83058 89720
rect 84658 92248 84714 92304
rect 84106 86536 84162 86592
rect 86682 92112 86738 92168
rect 85670 83952 85726 84008
rect 86866 77832 86922 77888
rect 87234 88032 87290 88088
rect 93260 92656 93316 92712
rect 91834 92384 91890 92440
rect 92754 86672 92810 86728
rect 91282 85176 91338 85232
rect 95882 241712 95938 241768
rect 96526 238720 96582 238776
rect 95146 103536 95202 103592
rect 95330 120264 95386 120320
rect 93122 83408 93178 83464
rect 89994 82728 90050 82784
rect 89902 80008 89958 80064
rect 97538 240080 97594 240136
rect 96710 233960 96766 234016
rect 97814 233960 97870 234016
rect 96710 145696 96766 145752
rect 96066 134000 96122 134056
rect 96618 133048 96674 133104
rect 96618 132232 96674 132288
rect 96618 130872 96674 130928
rect 96618 130056 96674 130112
rect 96066 120300 96068 120320
rect 96068 120300 96120 120320
rect 96120 120300 96122 120320
rect 96066 120264 96122 120300
rect 95974 105032 96030 105088
rect 96526 103400 96582 103456
rect 95882 92928 95938 92984
rect 96802 133864 96858 133920
rect 96710 127608 96766 127664
rect 97078 124616 97134 124672
rect 97170 123256 97226 123312
rect 97354 131416 97410 131472
rect 97538 127064 97594 127120
rect 97814 126248 97870 126304
rect 97814 124108 97816 124128
rect 97816 124108 97868 124128
rect 97868 124108 97870 124128
rect 97814 124072 97870 124108
rect 97262 122440 97318 122496
rect 97538 121624 97594 121680
rect 96986 120808 97042 120864
rect 97354 117000 97410 117056
rect 97906 119448 97962 119504
rect 97906 118652 97962 118688
rect 97906 118632 97908 118652
rect 97908 118632 97960 118652
rect 97960 118632 97962 118652
rect 97906 116456 97962 116512
rect 97906 115640 97962 115696
rect 97814 114824 97870 114880
rect 97814 114028 97870 114064
rect 97814 114008 97816 114028
rect 97816 114008 97868 114028
rect 97868 114008 97870 114028
rect 97906 113464 97962 113520
rect 97078 111868 97080 111888
rect 97080 111868 97132 111888
rect 97132 111868 97134 111888
rect 97078 111832 97134 111868
rect 96710 111016 96766 111072
rect 97906 110200 97962 110256
rect 97814 109656 97870 109712
rect 96710 107208 96766 107264
rect 97906 108024 97962 108080
rect 96802 104216 96858 104272
rect 97906 102856 97962 102912
rect 99378 280200 99434 280256
rect 98182 261296 98238 261352
rect 99286 258032 99342 258088
rect 98274 248784 98330 248840
rect 98734 242528 98790 242584
rect 99102 242392 99158 242448
rect 98734 241712 98790 241768
rect 98274 239944 98330 240000
rect 98734 239944 98790 240000
rect 98458 125432 98514 125488
rect 98090 108840 98146 108896
rect 97906 102076 97908 102096
rect 97908 102076 97960 102096
rect 97960 102076 97962 102096
rect 97906 102040 97962 102076
rect 97538 100408 97594 100464
rect 97906 99592 97962 99648
rect 97814 99048 97870 99104
rect 97906 98232 97962 98288
rect 98826 146376 98882 146432
rect 100114 282920 100170 282976
rect 100022 258984 100078 259040
rect 100850 283328 100906 283384
rect 100758 282648 100814 282704
rect 100758 278604 100760 278624
rect 100760 278604 100812 278624
rect 100812 278604 100814 278624
rect 100758 278568 100814 278604
rect 100758 276120 100814 276176
rect 100758 274488 100814 274544
rect 100850 273672 100906 273728
rect 100758 272856 100814 272912
rect 100758 270444 100760 270464
rect 100760 270444 100812 270464
rect 100812 270444 100814 270464
rect 100758 270408 100814 270444
rect 101678 281016 101734 281072
rect 105266 390360 105322 390416
rect 105542 388864 105598 388920
rect 103702 382064 103758 382120
rect 104254 382064 104310 382120
rect 101402 272040 101458 272096
rect 101126 271224 101182 271280
rect 100942 268776 100998 268832
rect 100758 267996 100760 268016
rect 100760 267996 100812 268016
rect 100812 267996 100814 268016
rect 100758 267960 100814 267996
rect 100758 266364 100760 266384
rect 100760 266364 100812 266384
rect 100812 266364 100814 266384
rect 100758 266328 100814 266364
rect 100758 265512 100814 265568
rect 100850 264696 100906 264752
rect 100758 263064 100814 263120
rect 100666 262248 100722 262304
rect 100942 262248 100998 262304
rect 100574 254904 100630 254960
rect 100114 247560 100170 247616
rect 96710 96600 96766 96656
rect 97078 95276 97080 95296
rect 97080 95276 97132 95296
rect 97132 95276 97134 95296
rect 97078 95240 97134 95276
rect 97906 96056 97962 96112
rect 97814 94424 97870 94480
rect 97906 93608 97962 93664
rect 96710 90364 96766 90400
rect 96710 90344 96712 90364
rect 96712 90344 96764 90364
rect 96764 90344 96766 90364
rect 96618 83408 96674 83464
rect 95146 75112 95202 75168
rect 98642 85448 98698 85504
rect 98642 85176 98698 85232
rect 100850 260616 100906 260672
rect 100758 259800 100814 259856
rect 100758 258168 100814 258224
rect 102046 257388 102048 257408
rect 102048 257388 102100 257408
rect 102100 257388 102102 257408
rect 102046 257352 102102 257388
rect 100758 256536 100814 256592
rect 100850 255720 100906 255776
rect 100758 254924 100814 254960
rect 100758 254904 100760 254924
rect 100760 254904 100812 254924
rect 100812 254904 100814 254924
rect 100758 254088 100814 254144
rect 100758 253272 100814 253328
rect 100850 252492 100852 252512
rect 100852 252492 100904 252512
rect 100904 252492 100906 252512
rect 100850 252456 100906 252492
rect 100758 251640 100814 251696
rect 100758 250824 100814 250880
rect 100850 250008 100906 250064
rect 100942 248376 100998 248432
rect 100942 246744 100998 246800
rect 101402 246200 101458 246256
rect 100942 245112 100998 245168
rect 101034 244296 101090 244352
rect 99470 101224 99526 101280
rect 98734 74432 98790 74488
rect 100298 100000 100354 100056
rect 100298 92248 100354 92304
rect 100114 92112 100170 92168
rect 102230 261432 102286 261488
rect 103426 281424 103482 281480
rect 103426 280200 103482 280256
rect 102230 242664 102286 242720
rect 104254 363568 104310 363624
rect 104438 304136 104494 304192
rect 103426 239944 103482 240000
rect 103426 238040 103482 238096
rect 102874 162832 102930 162888
rect 102966 144880 103022 144936
rect 102782 90344 102838 90400
rect 101678 88168 101734 88224
rect 101586 86536 101642 86592
rect 101494 77152 101550 77208
rect 97446 3440 97502 3496
rect 104438 244840 104494 244896
rect 104346 241848 104402 241904
rect 104254 225528 104310 225584
rect 104254 182824 104310 182880
rect 104162 83952 104218 84008
rect 106738 390360 106794 390416
rect 107750 390360 107806 390416
rect 107842 389272 107898 389328
rect 109682 384920 109738 384976
rect 107014 260752 107070 260808
rect 104806 150456 104862 150512
rect 104806 145696 104862 145752
rect 104346 139440 104402 139496
rect 104254 75112 104310 75168
rect 105450 90480 105506 90536
rect 106370 210296 106426 210352
rect 106370 209752 106426 209808
rect 105634 90480 105690 90536
rect 105450 89528 105506 89584
rect 106186 81368 106242 81424
rect 107474 108976 107530 109032
rect 110602 389408 110658 389464
rect 109682 260752 109738 260808
rect 115202 537376 115258 537432
rect 114742 442176 114798 442232
rect 113270 436872 113326 436928
rect 114558 430072 114614 430128
rect 113362 425992 113418 426048
rect 113270 416744 113326 416800
rect 113178 413752 113234 413808
rect 110602 238448 110658 238504
rect 108486 146956 108488 146976
rect 108488 146956 108540 146976
rect 108540 146956 108542 146976
rect 108486 146920 108542 146956
rect 108394 143656 108450 143712
rect 108302 90616 108358 90672
rect 107658 85312 107714 85368
rect 108118 85312 108174 85368
rect 108302 81096 108358 81152
rect 109682 87896 109738 87952
rect 112810 278160 112866 278216
rect 112442 242528 112498 242584
rect 111246 232464 111302 232520
rect 111154 219272 111210 219328
rect 113546 420008 113602 420064
rect 113454 402364 113456 402384
rect 113456 402364 113508 402384
rect 113508 402364 113510 402384
rect 113454 402328 113510 402364
rect 113362 384240 113418 384296
rect 113914 416744 113970 416800
rect 114650 417832 114706 417888
rect 115018 424088 115074 424144
rect 115018 423000 115074 423056
rect 115202 421912 115258 421968
rect 115754 433336 115810 433392
rect 115846 432248 115902 432304
rect 115846 431196 115848 431216
rect 115848 431196 115900 431216
rect 115900 431196 115902 431216
rect 115846 431160 115902 431196
rect 115846 428168 115902 428224
rect 115386 425992 115442 426048
rect 115386 424940 115388 424960
rect 115388 424940 115440 424960
rect 115440 424940 115442 424960
rect 115386 424904 115442 424940
rect 115754 420824 115810 420880
rect 116582 456864 116638 456920
rect 116582 437008 116638 437064
rect 116582 434696 116638 434752
rect 118698 461488 118754 461544
rect 118698 460944 118754 461000
rect 117962 448432 118018 448488
rect 117502 442312 117558 442368
rect 115846 415656 115902 415712
rect 115846 414840 115902 414896
rect 115294 412664 115350 412720
rect 114742 410488 114798 410544
rect 115846 411576 115902 411632
rect 115846 408584 115902 408640
rect 115386 407496 115442 407552
rect 115202 406408 115258 406464
rect 114926 405456 114982 405512
rect 114926 404368 114982 404424
rect 114742 400424 114798 400480
rect 115754 405612 115810 405648
rect 115754 405592 115756 405612
rect 115756 405592 115808 405612
rect 115808 405592 115810 405612
rect 115846 404504 115902 404560
rect 115846 403416 115902 403472
rect 115570 401240 115626 401296
rect 115846 399336 115902 399392
rect 115386 398248 115442 398304
rect 115202 397296 115258 397352
rect 115754 397296 115810 397352
rect 115294 397180 115350 397216
rect 115294 397160 115296 397180
rect 115296 397160 115348 397180
rect 115348 397160 115350 397180
rect 114926 396344 114982 396400
rect 115754 396208 115810 396264
rect 115846 395256 115902 395312
rect 115754 394168 115810 394224
rect 115570 393080 115626 393136
rect 115754 392012 115810 392048
rect 115754 391992 115756 392012
rect 115756 391992 115808 392012
rect 115808 391992 115810 392012
rect 114834 391176 114890 391232
rect 117226 391040 117282 391096
rect 116674 388048 116730 388104
rect 116674 387368 116730 387424
rect 116674 364928 116730 364984
rect 113914 284960 113970 285016
rect 113270 269320 113326 269376
rect 104530 3304 104586 3360
rect 112534 87896 112590 87952
rect 112994 87896 113050 87952
rect 113822 238176 113878 238232
rect 115202 226208 115258 226264
rect 114558 225528 114614 225584
rect 114466 167728 114522 167784
rect 114558 108976 114614 109032
rect 115294 108976 115350 109032
rect 116582 291216 116638 291272
rect 116490 281424 116546 281480
rect 116582 236680 116638 236736
rect 115938 137944 115994 138000
rect 116490 137944 116546 138000
rect 116490 137264 116546 137320
rect 120722 465160 120778 465216
rect 118882 433744 118938 433800
rect 119434 377304 119490 377360
rect 121458 388048 121514 388104
rect 122102 451288 122158 451344
rect 122838 441632 122894 441688
rect 122102 388456 122158 388512
rect 122102 356632 122158 356688
rect 119986 309168 120042 309224
rect 119342 292576 119398 292632
rect 117318 266600 117374 266656
rect 116766 235864 116822 235920
rect 116674 149640 116730 149696
rect 116674 117272 116730 117328
rect 116582 86672 116638 86728
rect 117962 138760 118018 138816
rect 118790 190984 118846 191040
rect 120814 291760 120870 291816
rect 120722 287136 120778 287192
rect 122194 331336 122250 331392
rect 122746 309304 122802 309360
rect 122102 236680 122158 236736
rect 120078 100000 120134 100056
rect 121458 88032 121514 88088
rect 124126 451832 124182 451888
rect 125598 388456 125654 388512
rect 124218 384920 124274 384976
rect 122838 304136 122894 304192
rect 124126 306856 124182 306912
rect 123482 77016 123538 77072
rect 124862 358672 124918 358728
rect 129738 581032 129794 581088
rect 128358 387776 128414 387832
rect 129002 387776 129058 387832
rect 129738 387640 129794 387696
rect 128358 386280 128414 386336
rect 127622 329976 127678 330032
rect 126334 327120 126390 327176
rect 126242 304952 126298 305008
rect 124954 289176 125010 289232
rect 124862 82728 124918 82784
rect 129002 336776 129058 336832
rect 128358 231104 128414 231160
rect 127806 158752 127862 158808
rect 129646 297472 129702 297528
rect 132498 435240 132554 435296
rect 130474 387640 130530 387696
rect 130382 377984 130438 378040
rect 130382 305088 130438 305144
rect 129186 242392 129242 242448
rect 131854 305224 131910 305280
rect 130658 263608 130714 263664
rect 130658 254496 130714 254552
rect 131854 226888 131910 226944
rect 133142 450064 133198 450120
rect 133142 437416 133198 437472
rect 133142 325896 133198 325952
rect 133326 281560 133382 281616
rect 133326 220768 133382 220824
rect 130382 3440 130438 3496
rect 136638 536696 136694 536752
rect 135994 347792 136050 347848
rect 134614 317600 134670 317656
rect 142158 538736 142214 538792
rect 140134 324400 140190 324456
rect 138754 298968 138810 299024
rect 141422 307944 141478 308000
rect 141514 293120 141570 293176
rect 147586 454144 147642 454200
rect 142802 314880 142858 314936
rect 142894 282104 142950 282160
rect 144274 227568 144330 227624
rect 147034 328480 147090 328536
rect 145654 139984 145710 140040
rect 151082 410080 151138 410136
rect 148414 375944 148470 376000
rect 148414 342216 148470 342272
rect 151082 377984 151138 378040
rect 149794 321680 149850 321736
rect 149702 314744 149758 314800
rect 149058 285640 149114 285696
rect 151082 320184 151138 320240
rect 151174 319368 151230 319424
rect 151174 294480 151230 294536
rect 148506 156032 148562 156088
rect 151082 266328 151138 266384
rect 149794 250416 149850 250472
rect 149794 223488 149850 223544
rect 153934 302504 153990 302560
rect 152738 282104 152794 282160
rect 152554 244840 152610 244896
rect 152554 229744 152610 229800
rect 152554 228248 152610 228304
rect 155222 304000 155278 304056
rect 154486 258712 154542 258768
rect 155314 244840 155370 244896
rect 155406 153176 155462 153232
rect 157982 375264 158038 375320
rect 158074 327664 158130 327720
rect 156694 233144 156750 233200
rect 156602 216552 156658 216608
rect 155866 143384 155922 143440
rect 156694 81232 156750 81288
rect 159362 369688 159418 369744
rect 159362 323040 159418 323096
rect 158074 136584 158130 136640
rect 159546 371184 159602 371240
rect 160742 372544 160798 372600
rect 160190 371320 160246 371376
rect 160742 371320 160798 371376
rect 160742 301552 160798 301608
rect 162766 324944 162822 325000
rect 162306 300056 162362 300112
rect 160742 237360 160798 237416
rect 159546 235864 159602 235920
rect 160006 235864 160062 235920
rect 160926 238584 160982 238640
rect 160926 237360 160982 237416
rect 162214 280064 162270 280120
rect 162398 278840 162454 278896
rect 162214 228248 162270 228304
rect 160742 180784 160798 180840
rect 161294 167592 161350 167648
rect 160742 155216 160798 155272
rect 160834 150592 160890 150648
rect 148322 3304 148378 3360
rect 160926 139984 160982 140040
rect 161478 151000 161534 151056
rect 161386 135904 161442 135960
rect 160926 128424 160982 128480
rect 165526 393352 165582 393408
rect 163686 265512 163742 265568
rect 167734 388728 167790 388784
rect 166262 316240 166318 316296
rect 166354 137808 166410 137864
rect 166446 94424 166502 94480
rect 166906 94424 166962 94480
rect 168378 380180 168434 380216
rect 168378 380160 168380 380180
rect 168380 380160 168432 380180
rect 168432 380160 168434 380180
rect 169206 404368 169262 404424
rect 169114 380160 169170 380216
rect 168378 240080 168434 240136
rect 168378 239264 168434 239320
rect 169206 369688 169262 369744
rect 173806 457000 173862 457056
rect 170494 387776 170550 387832
rect 170494 372000 170550 372056
rect 171046 372000 171102 372056
rect 170494 320320 170550 320376
rect 169206 312160 169262 312216
rect 169666 280880 169722 280936
rect 169114 240080 169170 240136
rect 169574 228928 169630 228984
rect 169574 162016 169630 162072
rect 170494 246200 170550 246256
rect 171782 310664 171838 310720
rect 171782 259528 171838 259584
rect 170954 239944 171010 240000
rect 171138 233960 171194 234016
rect 171046 202136 171102 202192
rect 170586 146512 170642 146568
rect 173070 388320 173126 388376
rect 173162 387504 173218 387560
rect 173070 382200 173126 382256
rect 176658 454280 176714 454336
rect 176658 454008 176714 454064
rect 173254 309440 173310 309496
rect 172426 175208 172482 175264
rect 172426 174528 172482 174584
rect 173346 247560 173402 247616
rect 174542 290400 174598 290456
rect 173714 240760 173770 240816
rect 173254 199280 173310 199336
rect 173254 75792 173310 75848
rect 175278 280744 175334 280800
rect 175186 237224 175242 237280
rect 175186 145560 175242 145616
rect 176014 220088 176070 220144
rect 179234 458360 179290 458416
rect 177946 454280 178002 454336
rect 177302 388320 177358 388376
rect 179234 449792 179290 449848
rect 179234 448568 179290 448624
rect 178038 389000 178094 389056
rect 178774 389000 178830 389056
rect 178682 379344 178738 379400
rect 177302 280880 177358 280936
rect 176014 92112 176070 92168
rect 177394 153720 177450 153776
rect 177394 149096 177450 149152
rect 177394 106256 177450 106312
rect 177394 75656 177450 75712
rect 178958 318824 179014 318880
rect 180154 454416 180210 454472
rect 180062 448568 180118 448624
rect 178958 255312 179014 255368
rect 178958 230424 179014 230480
rect 178774 112104 178830 112160
rect 179234 107616 179290 107672
rect 178774 77016 178830 77072
rect 182086 447888 182142 447944
rect 180246 388184 180302 388240
rect 180154 382200 180210 382256
rect 180154 302368 180210 302424
rect 180062 237904 180118 237960
rect 180062 229744 180118 229800
rect 180062 220088 180118 220144
rect 180062 135904 180118 135960
rect 181350 365744 181406 365800
rect 180798 288496 180854 288552
rect 180338 239944 180394 240000
rect 180706 233144 180762 233200
rect 181626 244840 181682 244896
rect 182086 320048 182142 320104
rect 183466 452920 183522 452976
rect 184202 439456 184258 439512
rect 184202 338680 184258 338736
rect 182270 240760 182326 240816
rect 181626 235320 181682 235376
rect 181534 234504 181590 234560
rect 182270 214648 182326 214704
rect 181442 167728 181498 167784
rect 181258 79872 181314 79928
rect 180154 72392 180210 72448
rect 184386 328616 184442 328672
rect 184202 305224 184258 305280
rect 184202 254496 184258 254552
rect 184202 240760 184258 240816
rect 187606 455504 187662 455560
rect 187514 452784 187570 452840
rect 187146 450200 187202 450256
rect 187054 448432 187110 448488
rect 187146 436736 187202 436792
rect 182086 79872 182142 79928
rect 183466 160792 183522 160848
rect 183098 143656 183154 143712
rect 184202 131144 184258 131200
rect 185490 129784 185546 129840
rect 184754 108160 184810 108216
rect 186134 292304 186190 292360
rect 186134 291216 186190 291272
rect 186042 253952 186098 254008
rect 187054 387640 187110 387696
rect 187146 383424 187202 383480
rect 186962 321544 187018 321600
rect 187698 415948 187754 415984
rect 187698 415928 187700 415948
rect 187700 415928 187752 415948
rect 187752 415928 187754 415948
rect 189722 459584 189778 459640
rect 188526 387232 188582 387288
rect 188434 385736 188490 385792
rect 188526 375264 188582 375320
rect 188894 327664 188950 327720
rect 187606 321544 187662 321600
rect 188342 317464 188398 317520
rect 188342 286320 188398 286376
rect 186410 282920 186466 282976
rect 187054 282920 187110 282976
rect 186962 241576 187018 241632
rect 186134 222808 186190 222864
rect 187146 238040 187202 238096
rect 188342 233824 188398 233880
rect 187054 162016 187110 162072
rect 186962 156576 187018 156632
rect 187054 144064 187110 144120
rect 186962 133864 187018 133920
rect 186318 108160 186374 108216
rect 186318 107752 186374 107808
rect 187514 91976 187570 92032
rect 186318 84088 186374 84144
rect 186318 82864 186374 82920
rect 186962 82864 187018 82920
rect 189078 327256 189134 327312
rect 191102 451424 191158 451480
rect 191010 447752 191066 447808
rect 191654 449112 191710 449168
rect 191654 446392 191710 446448
rect 191654 442040 191710 442096
rect 191654 441632 191710 441688
rect 191378 440680 191434 440736
rect 191378 439320 191434 439376
rect 191562 437960 191618 438016
rect 191562 435240 191618 435296
rect 190642 432248 190698 432304
rect 191102 430888 191158 430944
rect 190642 426808 190698 426864
rect 190642 422456 190698 422512
rect 190366 420960 190422 421016
rect 190642 415384 190698 415440
rect 191010 409944 191066 410000
rect 191010 408584 191066 408640
rect 190826 398520 190882 398576
rect 190826 395800 190882 395856
rect 190826 394440 190882 394496
rect 190458 393352 190514 393408
rect 190458 391720 190514 391776
rect 190366 327256 190422 327312
rect 189906 302232 189962 302288
rect 189814 295296 189870 295352
rect 189814 280744 189870 280800
rect 189722 247016 189778 247072
rect 189906 245656 189962 245712
rect 191010 298696 191066 298752
rect 191194 429528 191250 429584
rect 194598 466520 194654 466576
rect 192666 455640 192722 455696
rect 192482 436600 192538 436656
rect 191746 428168 191802 428224
rect 191746 425448 191802 425504
rect 191746 419736 191802 419792
rect 191746 418376 191802 418432
rect 191746 417016 191802 417072
rect 191746 414044 191802 414080
rect 191746 414024 191748 414044
rect 191748 414024 191800 414044
rect 191800 414024 191802 414044
rect 191746 411304 191802 411360
rect 191746 406952 191802 407008
rect 191746 405592 191802 405648
rect 191746 404232 191802 404288
rect 191654 402328 191710 402384
rect 191746 400152 191802 400208
rect 191746 397160 191802 397216
rect 191562 393080 191618 393136
rect 191470 299648 191526 299704
rect 191194 293256 191250 293312
rect 191286 292168 191342 292224
rect 191102 286728 191158 286784
rect 190458 282376 190514 282432
rect 190550 281288 190606 281344
rect 190458 279112 190514 279168
rect 190458 278044 190514 278080
rect 190458 278024 190460 278044
rect 190460 278024 190512 278044
rect 190512 278024 190514 278044
rect 190458 276936 190514 276992
rect 190458 275848 190514 275904
rect 190550 274780 190606 274816
rect 190550 274760 190552 274780
rect 190552 274760 190604 274780
rect 190604 274760 190606 274780
rect 190458 273672 190514 273728
rect 190826 272584 190882 272640
rect 190826 270408 190882 270464
rect 190826 265004 190828 265024
rect 190828 265004 190880 265024
rect 190880 265004 190882 265024
rect 190826 264968 190882 265004
rect 190458 258068 190460 258088
rect 190460 258068 190512 258088
rect 190512 258068 190514 258088
rect 190458 258032 190514 258068
rect 190642 256264 190698 256320
rect 190642 250824 190698 250880
rect 190826 249736 190882 249792
rect 189998 242936 190054 242992
rect 189998 236544 190054 236600
rect 189906 235184 189962 235240
rect 189814 233008 189870 233064
rect 189722 217232 189778 217288
rect 188434 166368 188490 166424
rect 188618 155216 188674 155272
rect 188526 145016 188582 145072
rect 188434 143520 188490 143576
rect 188618 144200 188674 144256
rect 190366 155216 190422 155272
rect 190274 134136 190330 134192
rect 190274 129784 190330 129840
rect 188066 96872 188122 96928
rect 188066 91976 188122 92032
rect 188342 84088 188398 84144
rect 189078 110744 189134 110800
rect 190182 94424 190238 94480
rect 188986 78512 189042 78568
rect 191562 296520 191618 296576
rect 191746 378936 191802 378992
rect 191746 373224 191802 373280
rect 191746 372816 191802 372872
rect 191746 367648 191802 367704
rect 192666 447888 192722 447944
rect 193126 445032 193182 445088
rect 194690 453056 194746 453112
rect 195794 458260 195796 458280
rect 195796 458260 195848 458280
rect 195848 458260 195850 458280
rect 195794 458224 195850 458260
rect 195978 452920 196034 452976
rect 197910 454144 197966 454200
rect 203154 453056 203210 453112
rect 207570 457000 207626 457056
rect 207110 454280 207166 454336
rect 205914 452784 205970 452840
rect 210422 458360 210478 458416
rect 209778 451424 209834 451480
rect 212446 452648 212502 452704
rect 211618 451832 211674 451888
rect 212722 455640 212778 455696
rect 214562 455504 214618 455560
rect 216862 459584 216918 459640
rect 220082 459584 220138 459640
rect 219806 457000 219862 457056
rect 220818 455504 220874 455560
rect 225050 453192 225106 453248
rect 224130 452648 224186 452704
rect 228086 450336 228142 450392
rect 231214 454144 231270 454200
rect 230478 450200 230534 450256
rect 233238 455640 233294 455696
rect 234894 454008 234950 454064
rect 234434 452648 234490 452704
rect 240138 460128 240194 460184
rect 238758 459584 238814 459640
rect 240138 459584 240194 459640
rect 237378 453192 237434 453248
rect 236734 451832 236790 451888
rect 220818 449928 220874 449984
rect 238482 449928 238538 449984
rect 242162 453872 242218 453928
rect 244002 453872 244058 453928
rect 244002 452920 244058 452976
rect 249246 458224 249302 458280
rect 247866 451288 247922 451344
rect 250626 456864 250682 456920
rect 253938 460944 253994 461000
rect 250626 452648 250682 452704
rect 244554 450064 244610 450120
rect 248510 449928 248566 449984
rect 193494 449656 193550 449712
rect 245750 449656 245806 449712
rect 253938 446120 253994 446176
rect 253938 440408 253994 440464
rect 253570 402056 253626 402112
rect 193494 390904 193550 390960
rect 252558 390904 252614 390960
rect 223486 390768 223542 390824
rect 195426 389136 195482 389192
rect 194506 389000 194562 389056
rect 193126 370504 193182 370560
rect 192574 315016 192630 315072
rect 192666 313928 192722 313984
rect 191746 299784 191802 299840
rect 191746 297608 191802 297664
rect 191746 291080 191802 291136
rect 191654 289992 191710 290048
rect 191654 288904 191710 288960
rect 191838 288360 191894 288416
rect 191746 287816 191802 287872
rect 191746 284552 191802 284608
rect 191746 283464 191802 283520
rect 191746 281288 191802 281344
rect 191470 280200 191526 280256
rect 191654 271496 191710 271552
rect 191562 269320 191618 269376
rect 191654 268232 191710 268288
rect 191654 266056 191710 266112
rect 191654 263880 191710 263936
rect 191654 262792 191710 262848
rect 191654 261704 191710 261760
rect 191654 260616 191710 260672
rect 191654 257352 191710 257408
rect 191654 255176 191710 255232
rect 191562 254088 191618 254144
rect 191654 253000 191710 253056
rect 191654 251912 191710 251968
rect 191746 238040 191802 238096
rect 191010 130056 191066 130112
rect 191194 129240 191250 129296
rect 191194 128444 191250 128480
rect 191194 128424 191196 128444
rect 191196 128424 191248 128444
rect 191248 128424 191250 128444
rect 192574 290944 192630 291000
rect 193218 315016 193274 315072
rect 193310 301044 193312 301064
rect 193312 301044 193364 301064
rect 193364 301044 193366 301064
rect 193310 301008 193366 301044
rect 197358 385056 197414 385112
rect 197358 383560 197414 383616
rect 198738 380704 198794 380760
rect 201130 388456 201186 388512
rect 200210 385736 200266 385792
rect 200210 380840 200266 380896
rect 200118 380160 200174 380216
rect 202142 380704 202198 380760
rect 205546 389272 205602 389328
rect 205546 387776 205602 387832
rect 204350 381520 204406 381576
rect 204258 372000 204314 372056
rect 202142 344256 202198 344312
rect 199382 331200 199438 331256
rect 198830 322904 198886 322960
rect 197358 306720 197414 306776
rect 197358 305224 197414 305280
rect 196622 303592 196678 303648
rect 196806 302232 196862 302288
rect 197910 306448 197966 306504
rect 197910 302776 197966 302832
rect 201682 329840 201738 329896
rect 201590 307808 201646 307864
rect 201038 302504 201094 302560
rect 200394 302368 200450 302424
rect 203062 310528 203118 310584
rect 206834 387776 206890 387832
rect 205546 345616 205602 345672
rect 213458 388320 213514 388376
rect 214562 387776 214618 387832
rect 213826 363568 213882 363624
rect 213826 361528 213882 361584
rect 205638 340856 205694 340912
rect 204350 313928 204406 313984
rect 204718 313384 204774 313440
rect 205730 339496 205786 339552
rect 207110 321680 207166 321736
rect 209042 317736 209098 317792
rect 213182 334056 213238 334112
rect 211802 315288 211858 315344
rect 209778 314880 209834 314936
rect 209042 302912 209098 302968
rect 210238 309440 210294 309496
rect 211434 310664 211490 310720
rect 213274 329976 213330 330032
rect 214562 365608 214618 365664
rect 215206 365608 215262 365664
rect 215206 364928 215262 364984
rect 215206 363568 215262 363624
rect 218242 387776 218298 387832
rect 216034 327120 216090 327176
rect 215942 325896 215998 325952
rect 215850 324400 215906 324456
rect 213642 307944 213698 308000
rect 212998 303864 213054 303920
rect 207938 301416 207994 301472
rect 198370 301280 198426 301336
rect 194230 301144 194286 301200
rect 214838 305088 214894 305144
rect 215390 304952 215446 305008
rect 220726 365744 220782 365800
rect 219438 332560 219494 332616
rect 220082 330384 220138 330440
rect 218702 314744 218758 314800
rect 218518 309304 218574 309360
rect 219622 306720 219678 306776
rect 220910 312024 220966 312080
rect 221002 311888 221058 311944
rect 222290 335416 222346 335472
rect 221554 333240 221610 333296
rect 222934 323040 222990 323096
rect 223670 325760 223726 325816
rect 225142 328480 225198 328536
rect 224222 306992 224278 307048
rect 225050 302912 225106 302968
rect 228362 388320 228418 388376
rect 228362 356632 228418 356688
rect 227718 336776 227774 336832
rect 226982 316240 227038 316296
rect 226522 306584 226578 306640
rect 227074 309712 227130 309768
rect 227442 304000 227498 304056
rect 226798 302776 226854 302832
rect 227718 301552 227774 301608
rect 228454 331336 228510 331392
rect 229926 317600 229982 317656
rect 228454 304136 228510 304192
rect 229190 303728 229246 303784
rect 231122 386280 231178 386336
rect 231122 359352 231178 359408
rect 230478 305632 230534 305688
rect 231214 342216 231270 342272
rect 231214 303592 231270 303648
rect 232778 304136 232834 304192
rect 232502 301688 232558 301744
rect 234250 386280 234306 386336
rect 234618 385600 234674 385656
rect 234618 380160 234674 380216
rect 238022 389816 238078 389872
rect 233882 366288 233938 366344
rect 233330 318824 233386 318880
rect 233974 308080 234030 308136
rect 234618 303592 234674 303648
rect 238114 388320 238170 388376
rect 238666 366424 238722 366480
rect 240046 361664 240102 361720
rect 239402 320320 239458 320376
rect 237378 309168 237434 309224
rect 238206 306856 238262 306912
rect 238850 303864 238906 303920
rect 242254 389000 242310 389056
rect 242162 371864 242218 371920
rect 240598 304952 240654 305008
rect 242898 385600 242954 385656
rect 242990 370504 243046 370560
rect 243542 370504 243598 370560
rect 242254 361528 242310 361584
rect 242806 308352 242862 308408
rect 242438 303728 242494 303784
rect 241794 302232 241850 302288
rect 242162 302232 242218 302288
rect 244922 371320 244978 371376
rect 243082 313928 243138 313984
rect 244922 309168 244978 309224
rect 247038 388864 247094 388920
rect 247590 388864 247646 388920
rect 249062 384920 249118 384976
rect 246394 327664 246450 327720
rect 246302 302776 246358 302832
rect 249522 384920 249578 384976
rect 249062 311208 249118 311264
rect 249614 306448 249670 306504
rect 248970 304544 249026 304600
rect 247866 303592 247922 303648
rect 246394 301688 246450 301744
rect 247222 301688 247278 301744
rect 247866 301688 247922 301744
rect 250810 307808 250866 307864
rect 251362 303592 251418 303648
rect 242070 301028 242126 301064
rect 242070 301008 242072 301028
rect 242072 301008 242124 301028
rect 242124 301008 242126 301028
rect 194690 300872 194746 300928
rect 209134 300872 209190 300928
rect 252466 300772 252468 300792
rect 252468 300772 252520 300792
rect 252520 300772 252522 300792
rect 252466 300736 252522 300772
rect 193494 298968 193550 299024
rect 192574 285640 192630 285696
rect 193126 285640 193182 285696
rect 193126 239808 193182 239864
rect 192574 236544 192630 236600
rect 193678 242800 193734 242856
rect 193770 241984 193826 242040
rect 194506 241984 194562 242040
rect 195794 242020 195796 242040
rect 195796 242020 195848 242040
rect 195848 242020 195850 242040
rect 195242 239672 195298 239728
rect 195794 241984 195850 242020
rect 248510 242020 248512 242040
rect 248512 242020 248564 242040
rect 248564 242020 248566 242040
rect 248510 241984 248566 242020
rect 193218 166232 193274 166288
rect 191930 164328 191986 164384
rect 191654 139848 191710 139904
rect 191654 137400 191710 137456
rect 191746 136312 191802 136368
rect 191746 135496 191802 135552
rect 191746 132776 191802 132832
rect 191746 127608 191802 127664
rect 191562 126520 191618 126576
rect 191470 123800 191526 123856
rect 191010 122984 191066 123040
rect 190550 118632 190606 118688
rect 191010 118632 191066 118688
rect 191746 122168 191802 122224
rect 191746 121388 191748 121408
rect 191748 121388 191800 121408
rect 191800 121388 191802 121408
rect 191746 121352 191802 121388
rect 191746 120264 191802 120320
rect 191746 119448 191802 119504
rect 191654 117544 191710 117600
rect 191010 115912 191066 115968
rect 190826 115096 190882 115152
rect 191102 109656 191158 109712
rect 191194 106120 191250 106176
rect 190550 97996 190552 98016
rect 190552 97996 190604 98016
rect 190604 97996 190606 98016
rect 190550 97960 190606 97996
rect 190458 97144 190514 97200
rect 191378 95376 191434 95432
rect 190458 93608 190514 93664
rect 190366 85448 190422 85504
rect 191562 100680 191618 100736
rect 191378 84768 191434 84824
rect 191746 116728 191802 116784
rect 191838 114008 191894 114064
rect 191746 113212 191802 113248
rect 191746 113192 191748 113212
rect 191748 113192 191800 113212
rect 191800 113192 191802 113212
rect 191746 112412 191748 112432
rect 191748 112412 191800 112432
rect 191800 112412 191802 112432
rect 191746 112376 191802 112412
rect 191746 110492 191802 110528
rect 191746 110472 191748 110492
rect 191748 110472 191800 110492
rect 191800 110472 191802 110492
rect 192022 108296 192078 108352
rect 192022 107616 192078 107672
rect 191746 106936 191802 106992
rect 191746 105032 191802 105088
rect 193034 138216 193090 138272
rect 192942 131960 192998 132016
rect 192482 104216 192538 104272
rect 191746 103400 191802 103456
rect 191746 101496 191802 101552
rect 191746 99864 191802 99920
rect 192850 93744 192906 93800
rect 193310 139984 193366 140040
rect 193402 138660 193404 138680
rect 193404 138660 193456 138680
rect 193456 138660 193458 138680
rect 193402 138624 193458 138660
rect 194690 147872 194746 147928
rect 193586 144200 193642 144256
rect 194690 143384 194746 143440
rect 195886 151952 195942 152008
rect 195242 141072 195298 141128
rect 196070 152088 196126 152144
rect 197358 237904 197414 237960
rect 197266 175888 197322 175944
rect 196622 143520 196678 143576
rect 196162 143384 196218 143440
rect 201406 205672 201462 205728
rect 198002 167592 198058 167648
rect 202878 233824 202934 233880
rect 202234 214512 202290 214568
rect 201406 167592 201462 167648
rect 198002 149776 198058 149832
rect 198830 148416 198886 148472
rect 201590 155216 201646 155272
rect 200302 147736 200358 147792
rect 201406 147736 201462 147792
rect 201590 145560 201646 145616
rect 201314 144064 201370 144120
rect 206282 222808 206338 222864
rect 204994 208936 205050 208992
rect 210422 217232 210478 217288
rect 209042 202272 209098 202328
rect 205638 174528 205694 174584
rect 204994 153720 205050 153776
rect 202878 140936 202934 140992
rect 204350 147600 204406 147656
rect 205454 140936 205510 140992
rect 196806 140392 196862 140448
rect 209042 167728 209098 167784
rect 207110 149776 207166 149832
rect 206558 140528 206614 140584
rect 208398 157392 208454 157448
rect 208582 157392 208638 157448
rect 208490 153720 208546 153776
rect 208490 151816 208546 151872
rect 213826 227568 213882 227624
rect 211802 189080 211858 189136
rect 211802 186904 211858 186960
rect 210422 169088 210478 169144
rect 213182 148416 213238 148472
rect 212354 147736 212410 147792
rect 211802 147600 211858 147656
rect 214562 226888 214618 226944
rect 214562 222128 214618 222184
rect 214010 175344 214066 175400
rect 217966 240760 218022 240816
rect 215298 233144 215354 233200
rect 215206 232464 215262 232520
rect 214562 171128 214618 171184
rect 213826 149640 213882 149696
rect 213274 144744 213330 144800
rect 212354 142432 212410 142488
rect 215206 148280 215262 148336
rect 215206 147736 215262 147792
rect 206558 140392 206614 140448
rect 218702 240760 218758 240816
rect 218150 235184 218206 235240
rect 218058 153040 218114 153096
rect 218702 224712 218758 224768
rect 222106 236580 222108 236600
rect 222108 236580 222160 236600
rect 222160 236580 222162 236600
rect 219530 235184 219586 235240
rect 220818 217368 220874 217424
rect 219530 169768 219586 169824
rect 219438 168952 219494 169008
rect 218242 154536 218298 154592
rect 218242 153040 218298 153096
rect 218242 142432 218298 142488
rect 222106 236544 222162 236580
rect 222842 231784 222898 231840
rect 223486 231784 223542 231840
rect 220266 169768 220322 169824
rect 220358 168952 220414 169008
rect 220266 154536 220322 154592
rect 221002 149096 221058 149152
rect 222198 161472 222254 161528
rect 222014 149096 222070 149152
rect 222014 146240 222070 146296
rect 221922 142160 221978 142216
rect 223670 166232 223726 166288
rect 222290 144608 222346 144664
rect 223026 144608 223082 144664
rect 223026 143656 223082 143712
rect 223578 140800 223634 140856
rect 224498 140392 224554 140448
rect 193126 124888 193182 124944
rect 193034 102584 193090 102640
rect 192942 86128 192998 86184
rect 225050 128968 225106 129024
rect 227718 233960 227774 234016
rect 225326 140120 225382 140176
rect 225418 130872 225474 130928
rect 226154 128424 226210 128480
rect 225234 116728 225290 116784
rect 225050 113736 225106 113792
rect 193218 104080 193274 104136
rect 193218 96328 193274 96384
rect 193218 95376 193274 95432
rect 193218 92248 193274 92304
rect 194506 92656 194562 92712
rect 194506 72392 194562 72448
rect 196530 89528 196586 89584
rect 197082 86808 197138 86864
rect 198370 88168 198426 88224
rect 202234 93336 202290 93392
rect 224774 93336 224830 93392
rect 224498 93200 224554 93256
rect 200302 92792 200358 92848
rect 201038 92792 201094 92848
rect 200762 92112 200818 92168
rect 203706 90616 203762 90672
rect 203522 90344 203578 90400
rect 204442 90480 204498 90536
rect 203706 81232 203762 81288
rect 204442 87488 204498 87544
rect 206098 92384 206154 92440
rect 205546 92112 205602 92168
rect 205638 91976 205694 92032
rect 208398 92792 208454 92848
rect 208674 90208 208730 90264
rect 209686 90208 209742 90264
rect 209226 87896 209282 87952
rect 207662 77152 207718 77208
rect 210422 92928 210478 92984
rect 210330 89800 210386 89856
rect 212170 92656 212226 92712
rect 212170 90888 212226 90944
rect 211618 89664 211674 89720
rect 210054 79872 210110 79928
rect 214562 92384 214618 92440
rect 215298 90208 215354 90264
rect 216402 90208 216458 90264
rect 218794 92520 218850 92576
rect 221922 86672 221978 86728
rect 220082 85448 220138 85504
rect 220174 80008 220230 80064
rect 224038 92792 224094 92848
rect 225142 109656 225198 109712
rect 225234 97144 225290 97200
rect 226246 97144 226302 97200
rect 230386 225528 230442 225584
rect 229098 223488 229154 223544
rect 230386 223488 230442 223544
rect 227810 220768 227866 220824
rect 227810 162832 227866 162888
rect 227718 156032 227774 156088
rect 229098 158752 229154 158808
rect 227994 150456 228050 150512
rect 226798 146512 226854 146568
rect 226522 137128 226578 137184
rect 226522 135496 226578 135552
rect 227626 139032 227682 139088
rect 226798 136312 226854 136368
rect 226706 134680 226762 134736
rect 226982 134680 227038 134736
rect 226706 133592 226762 133648
rect 226890 132776 226946 132832
rect 226706 131960 226762 132016
rect 226614 130056 226670 130112
rect 226614 127336 226670 127392
rect 226890 126520 226946 126576
rect 226430 125704 226486 125760
rect 226614 124616 226670 124672
rect 226522 123836 226524 123856
rect 226524 123836 226576 123856
rect 226576 123836 226578 123856
rect 226522 123800 226578 123836
rect 226706 122984 226762 123040
rect 226522 122168 226578 122224
rect 227166 129276 227168 129296
rect 227168 129276 227220 129296
rect 227220 129276 227222 129296
rect 227166 129240 227222 129276
rect 226706 120264 226762 120320
rect 226706 118360 226762 118416
rect 226614 117544 226670 117600
rect 226706 115948 226708 115968
rect 226708 115948 226760 115968
rect 226760 115948 226762 115968
rect 226706 115912 226762 115948
rect 226706 114824 226762 114880
rect 226614 114008 226670 114064
rect 226706 112104 226762 112160
rect 227810 138624 227866 138680
rect 232502 222808 232558 222864
rect 229190 146376 229246 146432
rect 231766 148416 231822 148472
rect 230478 144880 230534 144936
rect 231122 144880 231178 144936
rect 229282 143520 229338 143576
rect 231766 143520 231822 143576
rect 227718 110744 227774 110800
rect 227074 110472 227130 110528
rect 226430 108568 226486 108624
rect 226706 107752 226762 107808
rect 226798 106936 226854 106992
rect 226706 105848 226762 105904
rect 226430 105032 226486 105088
rect 226338 95104 226394 95160
rect 226338 94424 226394 94480
rect 226706 104216 226762 104272
rect 226614 103400 226670 103456
rect 226706 102312 226762 102368
rect 226522 101496 226578 101552
rect 226706 100680 226762 100736
rect 226614 99592 226670 99648
rect 227350 97960 227406 98016
rect 227718 97960 227774 98016
rect 226706 96056 226762 96112
rect 227534 95104 227590 95160
rect 226890 93608 226946 93664
rect 227810 95784 227866 95840
rect 227810 84088 227866 84144
rect 229098 75792 229154 75848
rect 230570 75656 230626 75712
rect 231950 92248 232006 92304
rect 234618 157936 234674 157992
rect 235998 217912 236054 217968
rect 237286 217912 237342 217968
rect 236734 89664 236790 89720
rect 233238 77016 233294 77072
rect 240138 220088 240194 220144
rect 240138 153176 240194 153232
rect 239402 90888 239458 90944
rect 247038 240080 247094 240136
rect 246302 239400 246358 239456
rect 246302 226208 246358 226264
rect 245658 224984 245714 225040
rect 246302 224984 246358 225040
rect 246302 95784 246358 95840
rect 247682 232600 247738 232656
rect 247682 147872 247738 147928
rect 251914 240080 251970 240136
rect 252282 239944 252338 240000
rect 252466 145560 252522 145616
rect 250442 92112 250498 92168
rect 254030 415112 254086 415168
rect 254122 412392 254178 412448
rect 254674 446120 254730 446176
rect 255502 454416 255558 454472
rect 255962 450064 256018 450120
rect 255502 448840 255558 448896
rect 255410 447480 255466 447536
rect 255410 444760 255466 444816
rect 255410 443420 255466 443456
rect 255410 443400 255412 443420
rect 255412 443400 255464 443420
rect 255464 443400 255466 443420
rect 255410 442060 255466 442096
rect 255410 442040 255412 442060
rect 255412 442040 255464 442060
rect 255464 442040 255466 442060
rect 255318 439048 255374 439104
rect 255410 437688 255466 437744
rect 255410 436328 255466 436384
rect 255410 434968 255466 435024
rect 255410 433608 255466 433664
rect 255410 431996 255466 432032
rect 255410 431976 255412 431996
rect 255412 431976 255464 431996
rect 255464 431976 255466 431996
rect 254674 431160 254730 431216
rect 255410 430616 255466 430672
rect 255502 429256 255558 429312
rect 255410 427896 255466 427952
rect 255502 426536 255558 426592
rect 255870 425176 255926 425232
rect 255502 423544 255558 423600
rect 255502 422184 255558 422240
rect 255502 420824 255558 420880
rect 255410 419464 255466 419520
rect 255502 418104 255558 418160
rect 255410 416744 255466 416800
rect 255410 413752 255466 413808
rect 255410 411032 255466 411088
rect 255410 409672 255466 409728
rect 255318 408312 255374 408368
rect 254214 405320 254270 405376
rect 254122 390496 254178 390552
rect 255410 406952 255466 407008
rect 255410 401240 255466 401296
rect 255410 399880 255466 399936
rect 255318 396888 255374 396944
rect 255502 395528 255558 395584
rect 254582 367648 254638 367704
rect 253938 346976 253994 347032
rect 253938 330384 253994 330440
rect 253294 305632 253350 305688
rect 252834 300192 252890 300248
rect 252834 299784 252890 299840
rect 252834 292440 252890 292496
rect 253294 298016 253350 298072
rect 253846 292576 253902 292632
rect 252926 292032 252982 292088
rect 253846 291780 253902 291816
rect 253846 291760 253848 291780
rect 253848 291760 253900 291780
rect 253900 291760 253902 291780
rect 254030 301416 254086 301472
rect 255594 392808 255650 392864
rect 254766 328344 254822 328400
rect 254766 327256 254822 327312
rect 254582 301552 254638 301608
rect 254122 298560 254178 298616
rect 254030 295432 254086 295488
rect 254122 252728 254178 252784
rect 253938 246336 253994 246392
rect 252926 245792 252982 245848
rect 252834 244976 252890 245032
rect 252834 244432 252890 244488
rect 252834 242392 252890 242448
rect 254030 245520 254086 245576
rect 253938 242936 253994 242992
rect 253938 240080 253994 240136
rect 254030 217232 254086 217288
rect 254766 313384 254822 313440
rect 255502 313384 255558 313440
rect 255410 301144 255466 301200
rect 255318 300736 255374 300792
rect 255410 299920 255466 299976
rect 255318 299512 255374 299568
rect 255318 298560 255374 298616
rect 255410 298172 255466 298208
rect 255410 298152 255412 298172
rect 255412 298152 255464 298172
rect 255464 298152 255466 298172
rect 255410 297336 255466 297392
rect 255686 375944 255742 376000
rect 259642 465160 259698 465216
rect 256790 403960 256846 404016
rect 256882 394168 256938 394224
rect 258262 377304 258318 377360
rect 256698 316104 256754 316160
rect 255686 306992 255742 307048
rect 255594 300328 255650 300384
rect 255410 295160 255466 295216
rect 255502 294344 255558 294400
rect 255410 293972 255412 293992
rect 255412 293972 255464 293992
rect 255464 293972 255466 293992
rect 255410 293936 255466 293972
rect 255502 293120 255558 293176
rect 255318 280200 255374 280256
rect 255318 279384 255374 279440
rect 255318 276392 255374 276448
rect 255318 275032 255374 275088
rect 255318 273808 255374 273864
rect 255318 273128 255374 273184
rect 255318 272040 255374 272096
rect 255318 269864 255374 269920
rect 255318 266872 255374 266928
rect 255318 264832 255374 264888
rect 254674 251504 254730 251560
rect 254674 249736 254730 249792
rect 255318 244704 255374 244760
rect 255502 282376 255558 282432
rect 255502 281016 255558 281072
rect 255502 278976 255558 279032
rect 255502 278432 255558 278488
rect 255502 277244 255504 277264
rect 255504 277244 255556 277264
rect 255556 277244 255558 277264
rect 255502 277208 255558 277244
rect 255502 275476 255504 275496
rect 255504 275476 255556 275496
rect 255556 275476 255558 275496
rect 255502 275440 255558 275476
rect 255502 274252 255504 274272
rect 255504 274252 255556 274272
rect 255556 274252 255558 274272
rect 255502 274216 255558 274252
rect 255502 272448 255558 272504
rect 255502 271224 255558 271280
rect 255502 270816 255558 270872
rect 255502 270428 255558 270464
rect 255502 270408 255504 270428
rect 255504 270408 255556 270428
rect 255556 270408 255558 270428
rect 255502 267844 255558 267880
rect 255502 267824 255504 267844
rect 255504 267824 255556 267844
rect 255556 267824 255558 267844
rect 255502 266056 255558 266112
rect 255502 265648 255558 265704
rect 255502 263880 255558 263936
rect 255502 243344 255558 243400
rect 255502 242392 255558 242448
rect 255502 242120 255558 242176
rect 255410 232464 255466 232520
rect 255778 299648 255834 299704
rect 255686 299104 255742 299160
rect 256698 301416 256754 301472
rect 255962 297064 256018 297120
rect 256606 296520 256662 296576
rect 255870 296112 255926 296168
rect 255686 293528 255742 293584
rect 256146 292032 256202 292088
rect 256422 291352 256478 291408
rect 256606 291352 256662 291408
rect 256146 291216 256202 291272
rect 256514 289992 256570 290048
rect 255962 288768 256018 288824
rect 256606 288360 256662 288416
rect 255870 287952 255926 288008
rect 255778 287544 255834 287600
rect 256606 287272 256662 287328
rect 256514 286864 256570 286920
rect 256422 286184 256478 286240
rect 256330 283192 256386 283248
rect 256606 286628 256608 286648
rect 256608 286628 256660 286648
rect 256660 286628 256662 286648
rect 256606 286592 256662 286628
rect 256606 285368 256662 285424
rect 256606 284008 256662 284064
rect 256882 324400 256938 324456
rect 257434 316104 257490 316160
rect 256882 290944 256938 291000
rect 258722 396616 258778 396672
rect 258722 328616 258778 328672
rect 258354 319368 258410 319424
rect 259458 323620 259460 323640
rect 259460 323620 259512 323640
rect 259512 323620 259514 323640
rect 259458 323584 259514 323620
rect 258814 321544 258870 321600
rect 259366 319388 259422 319424
rect 259366 319368 259368 319388
rect 259368 319368 259420 319388
rect 259420 319368 259422 319388
rect 260838 380840 260894 380896
rect 260838 370504 260894 370560
rect 258814 302776 258870 302832
rect 258538 294752 258594 294808
rect 258538 293120 258594 293176
rect 258354 289720 258410 289776
rect 258354 284960 258410 285016
rect 258170 283600 258226 283656
rect 259274 283464 259330 283520
rect 256606 281968 256662 282024
rect 259274 281424 259330 281480
rect 255686 279792 255742 279848
rect 255686 278160 255742 278216
rect 256606 269048 256662 269104
rect 256422 263472 256478 263528
rect 256606 261296 256662 261352
rect 256606 260108 256608 260128
rect 256608 260108 256660 260128
rect 256660 260108 256662 260128
rect 256606 260072 256662 260108
rect 255962 259256 256018 259312
rect 256606 258848 256662 258904
rect 256330 257080 256386 257136
rect 256606 256672 256662 256728
rect 256606 256264 256662 256320
rect 256606 255332 256662 255368
rect 256606 255312 256608 255332
rect 256608 255312 256660 255332
rect 256660 255312 256662 255332
rect 256606 254496 256662 254552
rect 255778 253272 255834 253328
rect 256422 252320 256478 252376
rect 256606 251504 256662 251560
rect 256606 250688 256662 250744
rect 256606 250280 256662 250336
rect 256238 249328 256294 249384
rect 256606 248920 256662 248976
rect 256514 247152 256570 247208
rect 256606 246744 256662 246800
rect 256514 246200 256570 246256
rect 255686 244160 255742 244216
rect 255778 243752 255834 243808
rect 255778 241440 255834 241496
rect 256882 263064 256938 263120
rect 256882 240760 256938 240816
rect 254122 211792 254178 211848
rect 253846 208936 253902 208992
rect 255962 204856 256018 204912
rect 253202 166368 253258 166424
rect 252558 92520 252614 92576
rect 255318 175752 255374 175808
rect 255318 175344 255374 175400
rect 253938 89528 253994 89584
rect 256054 175752 256110 175808
rect 259458 278024 259514 278080
rect 258078 272720 258134 272776
rect 257342 240216 257398 240272
rect 258262 257488 258318 257544
rect 258170 255720 258226 255776
rect 258354 237904 258410 237960
rect 258262 222808 258318 222864
rect 256606 140936 256662 140992
rect 259642 298016 259698 298072
rect 259550 276800 259606 276856
rect 260930 333240 260986 333296
rect 260838 284824 260894 284880
rect 263598 452920 263654 452976
rect 262310 436872 262366 436928
rect 263414 436872 263470 436928
rect 261666 380840 261722 380896
rect 261666 379208 261722 379264
rect 262218 277480 262274 277536
rect 260930 272720 260986 272776
rect 262218 271768 262274 271824
rect 262218 271496 262274 271552
rect 261022 266464 261078 266520
rect 260838 264424 260894 264480
rect 259734 254088 259790 254144
rect 260930 253680 260986 253736
rect 260930 243616 260986 243672
rect 261206 246200 261262 246256
rect 261114 242256 261170 242312
rect 261114 233960 261170 234016
rect 261206 217912 261262 217968
rect 262126 217232 262182 217288
rect 259458 150592 259514 150648
rect 260102 140936 260158 140992
rect 259366 87488 259422 87544
rect 259550 83408 259606 83464
rect 263690 347792 263746 347848
rect 262862 317600 262918 317656
rect 263506 292440 263562 292496
rect 263874 324944 263930 325000
rect 263690 286864 263746 286920
rect 263506 282920 263562 282976
rect 263230 260108 263232 260128
rect 263232 260108 263284 260128
rect 263284 260108 263286 260128
rect 263230 260072 263286 260108
rect 262402 237224 262458 237280
rect 262494 230424 262550 230480
rect 265070 377984 265126 378040
rect 263782 273536 263838 273592
rect 263782 262792 263838 262848
rect 263874 262656 263930 262712
rect 263782 260888 263838 260944
rect 263874 236544 263930 236600
rect 265070 259392 265126 259448
rect 266450 382200 266506 382256
rect 266358 320184 266414 320240
rect 266358 285912 266414 285968
rect 266358 284416 266414 284472
rect 265254 269728 265310 269784
rect 265254 269320 265310 269376
rect 265806 263336 265862 263392
rect 265254 238584 265310 238640
rect 266634 295160 266690 295216
rect 267002 295160 267058 295216
rect 266634 284416 266690 284472
rect 266450 271768 266506 271824
rect 267922 304952 267978 305008
rect 267738 257388 267740 257408
rect 267740 257388 267792 257408
rect 267792 257388 267794 257408
rect 267738 257352 267794 257388
rect 269302 387504 269358 387560
rect 269302 312160 269358 312216
rect 269210 291216 269266 291272
rect 269118 288360 269174 288416
rect 269118 287272 269174 287328
rect 268014 285640 268070 285696
rect 267830 153040 267886 153096
rect 268290 242392 268346 242448
rect 268382 222128 268438 222184
rect 269394 283464 269450 283520
rect 269302 278024 269358 278080
rect 270774 308352 270830 308408
rect 270498 275168 270554 275224
rect 269210 218048 269266 218104
rect 262218 77832 262274 77888
rect 269394 233824 269450 233880
rect 269118 82048 269174 82104
rect 270590 273808 270646 273864
rect 270498 209752 270554 209808
rect 273350 383424 273406 383480
rect 271878 275984 271934 276040
rect 270774 266736 270830 266792
rect 271878 259392 271934 259448
rect 270774 232600 270830 232656
rect 272154 302776 272210 302832
rect 272154 288360 272210 288416
rect 272154 281424 272210 281480
rect 272154 280336 272210 280392
rect 273258 275984 273314 276040
rect 272154 224848 272210 224904
rect 271970 213832 272026 213888
rect 280158 460128 280214 460184
rect 273902 388864 273958 388920
rect 273442 303728 273498 303784
rect 273350 268096 273406 268152
rect 273350 265104 273406 265160
rect 277398 450336 277454 450392
rect 274730 380160 274786 380216
rect 274638 304952 274694 305008
rect 273534 288632 273590 288688
rect 273534 284824 273590 284880
rect 275006 306448 275062 306504
rect 274822 296928 274878 296984
rect 274730 281424 274786 281480
rect 274914 250144 274970 250200
rect 274914 216552 274970 216608
rect 270498 94696 270554 94752
rect 273258 86128 273314 86184
rect 277398 313248 277454 313304
rect 276294 302232 276350 302288
rect 276202 281696 276258 281752
rect 276386 255312 276442 255368
rect 276294 217232 276350 217288
rect 276018 131688 276074 131744
rect 277398 273128 277454 273184
rect 279422 375264 279478 375320
rect 277398 268096 277454 268152
rect 277490 240216 277546 240272
rect 278686 273128 278742 273184
rect 580906 697176 580962 697232
rect 582470 683848 582526 683904
rect 582378 630808 582434 630864
rect 580170 484608 580226 484664
rect 284298 458224 284354 458280
rect 282826 389000 282882 389056
rect 280802 311072 280858 311128
rect 280526 299512 280582 299568
rect 280250 262112 280306 262168
rect 280434 291352 280490 291408
rect 281446 151952 281502 152008
rect 280158 97416 280214 97472
rect 281630 301688 281686 301744
rect 281722 153720 281778 153776
rect 284298 318688 284354 318744
rect 284298 293120 284354 293176
rect 283102 248648 283158 248704
rect 284574 318688 284630 318744
rect 284574 317464 284630 317520
rect 284390 242120 284446 242176
rect 285678 259528 285734 259584
rect 284390 81232 284446 81288
rect 284298 78512 284354 78568
rect 285862 309168 285918 309224
rect 285770 253136 285826 253192
rect 287058 247424 287114 247480
rect 285862 144744 285918 144800
rect 286782 144744 286838 144800
rect 287334 389000 287390 389056
rect 287334 247424 287390 247480
rect 288622 387640 288678 387696
rect 289910 385076 289966 385112
rect 289910 385056 289912 385076
rect 289912 385056 289964 385076
rect 289964 385056 289966 385076
rect 289818 307808 289874 307864
rect 287058 88168 287114 88224
rect 286322 3304 286378 3360
rect 291198 295160 291254 295216
rect 291474 295296 291530 295352
rect 292578 268504 292634 268560
rect 291842 142432 291898 142488
rect 580170 458088 580226 458144
rect 298098 451832 298154 451888
rect 295430 296792 295486 296848
rect 295338 269728 295394 269784
rect 582654 670656 582710 670712
rect 582562 644000 582618 644056
rect 582470 431568 582526 431624
rect 582746 617480 582802 617536
rect 582838 590960 582894 591016
rect 582746 577632 582802 577688
rect 582654 456048 582710 456104
rect 582562 397976 582618 398032
rect 582562 378392 582618 378448
rect 582470 365064 582526 365120
rect 579618 325216 579674 325272
rect 580170 298696 580226 298752
rect 580262 272176 580318 272232
rect 580906 258848 580962 258904
rect 583022 564304 583078 564360
rect 582930 524456 582986 524512
rect 583114 537784 583170 537840
rect 583298 511264 583354 511320
rect 583206 471416 583262 471472
rect 583022 418240 583078 418296
rect 583298 404912 583354 404968
rect 583022 379344 583078 379400
rect 582654 351872 582710 351928
rect 582654 312024 582710 312080
rect 582562 289856 582618 289912
rect 582378 245520 582434 245576
rect 580170 232328 580226 232384
rect 580262 219000 580318 219056
rect 580354 205672 580410 205728
rect 580170 192500 580226 192536
rect 580170 192480 580172 192500
rect 580172 192480 580224 192500
rect 580224 192480 580226 192500
rect 580170 179152 580226 179208
rect 298098 72392 298154 72448
rect 293682 3304 293738 3360
rect 300122 3576 300178 3632
rect 302882 3440 302938 3496
rect 304354 3576 304410 3632
rect 305550 3440 305606 3496
rect 317418 148280 317474 148336
rect 313278 137264 313334 137320
rect 318798 32408 318854 32464
rect 327722 84768 327778 84824
rect 582378 125976 582434 126032
rect 580170 86128 580226 86184
rect 582378 72936 582434 72992
rect 580170 46280 580226 46336
rect 583114 303864 583170 303920
rect 582654 250416 582710 250472
rect 582930 165824 582986 165880
rect 582654 152632 582710 152688
rect 582654 138624 582710 138680
rect 582838 154536 582894 154592
rect 583022 139304 583078 139360
rect 582838 112784 582894 112840
rect 582838 99456 582894 99512
rect 582838 88168 582894 88224
rect 582838 80688 582894 80744
rect 582746 59608 582802 59664
rect 582654 19760 582710 19816
rect 582930 79328 582986 79384
rect 582930 33088 582986 33144
rect 582838 6568 582894 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580901 697234 580967 697237
rect 583520 697234 584960 697324
rect 580901 697232 584960 697234
rect 580901 697176 580906 697232
rect 580962 697176 584960 697232
rect 580901 697174 584960 697176
rect 580901 697171 580967 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582465 683906 582531 683909
rect 583520 683906 584960 683996
rect 582465 683904 584960 683906
rect 582465 683848 582470 683904
rect 582526 683848 584960 683904
rect 582465 683846 584960 683848
rect 582465 683843 582531 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 582649 670714 582715 670717
rect 583520 670714 584960 670804
rect 582649 670712 584960 670714
rect 582649 670656 582654 670712
rect 582710 670656 584960 670712
rect 582649 670654 584960 670656
rect 582649 670651 582715 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582557 644058 582623 644061
rect 583520 644058 584960 644148
rect 582557 644056 584960 644058
rect 582557 644000 582562 644056
rect 582618 644000 584960 644056
rect 582557 643998 584960 644000
rect 582557 643995 582623 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582373 630866 582439 630869
rect 583520 630866 584960 630956
rect 582373 630864 584960 630866
rect 582373 630808 582378 630864
rect 582434 630808 584960 630864
rect 582373 630806 584960 630808
rect 582373 630803 582439 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect 71773 596322 71839 596325
rect 75862 596322 75868 596324
rect 71773 596320 75868 596322
rect 71773 596264 71778 596320
rect 71834 596264 75868 596320
rect 71773 596262 75868 596264
rect 71773 596259 71839 596262
rect 75862 596260 75868 596262
rect 75932 596260 75938 596324
rect -960 592908 480 593148
rect 582833 591018 582899 591021
rect 583520 591018 584960 591108
rect 582833 591016 584960 591018
rect 582833 590960 582838 591016
rect 582894 590960 584960 591016
rect 582833 590958 584960 590960
rect 582833 590955 582899 590958
rect 583520 590868 584960 590958
rect 85481 583946 85547 583949
rect 101397 583946 101463 583949
rect 85481 583944 101463 583946
rect 85481 583888 85486 583944
rect 85542 583888 101402 583944
rect 101458 583888 101463 583944
rect 85481 583886 101463 583888
rect 85481 583883 85547 583886
rect 101397 583883 101463 583886
rect 92105 583810 92171 583813
rect 119337 583810 119403 583813
rect 92105 583808 119403 583810
rect 92105 583752 92110 583808
rect 92166 583752 119342 583808
rect 119398 583752 119403 583808
rect 92105 583750 119403 583752
rect 92105 583747 92171 583750
rect 119337 583747 119403 583750
rect 41321 582586 41387 582589
rect 82997 582586 83063 582589
rect 41321 582584 83063 582586
rect 41321 582528 41326 582584
rect 41382 582528 83002 582584
rect 83058 582528 83063 582584
rect 41321 582526 83063 582528
rect 41321 582523 41387 582526
rect 82997 582523 83063 582526
rect 88241 582586 88307 582589
rect 104157 582586 104223 582589
rect 88241 582584 104223 582586
rect 88241 582528 88246 582584
rect 88302 582528 104162 582584
rect 104218 582528 104223 582584
rect 88241 582526 104223 582528
rect 88241 582523 88307 582526
rect 104157 582523 104223 582526
rect 80697 582450 80763 582453
rect 83406 582450 83412 582452
rect 80697 582448 83412 582450
rect 80697 582392 80702 582448
rect 80758 582392 83412 582448
rect 80697 582390 83412 582392
rect 80697 582387 80763 582390
rect 83406 582388 83412 582390
rect 83476 582388 83482 582452
rect 74257 581226 74323 581229
rect 74257 581224 84210 581226
rect 74257 581168 74262 581224
rect 74318 581168 84210 581224
rect 74257 581166 84210 581168
rect 74257 581163 74323 581166
rect 75361 581090 75427 581093
rect 75678 581090 75684 581092
rect 75361 581088 75684 581090
rect 75361 581032 75366 581088
rect 75422 581032 75684 581088
rect 75361 581030 75684 581032
rect 75361 581027 75427 581030
rect 75678 581028 75684 581030
rect 75748 581028 75754 581092
rect 84150 581090 84210 581166
rect 129733 581090 129799 581093
rect 84150 581088 129799 581090
rect 84150 581032 129738 581088
rect 129794 581032 129799 581088
rect 84150 581030 129799 581032
rect 129733 581027 129799 581030
rect 71497 580818 71563 580821
rect 71630 580818 71636 580820
rect 71497 580816 71636 580818
rect 71497 580760 71502 580816
rect 71558 580760 71636 580816
rect 71497 580758 71636 580760
rect 71497 580755 71563 580758
rect 71630 580756 71636 580758
rect 71700 580756 71706 580820
rect 72417 580818 72483 580821
rect 79869 580820 79935 580821
rect 72918 580818 72924 580820
rect 72417 580816 72924 580818
rect 72417 580760 72422 580816
rect 72478 580760 72924 580816
rect 72417 580758 72924 580760
rect 72417 580755 72483 580758
rect 72918 580756 72924 580758
rect 72988 580756 72994 580820
rect 79869 580816 79916 580820
rect 79980 580818 79986 580820
rect 79869 580760 79874 580816
rect 79869 580756 79916 580760
rect 79980 580758 80026 580818
rect 79980 580756 79986 580758
rect 88374 580756 88380 580820
rect 88444 580818 88450 580820
rect 88701 580818 88767 580821
rect 88444 580816 88767 580818
rect 88444 580760 88706 580816
rect 88762 580760 88767 580816
rect 88444 580758 88767 580760
rect 88444 580756 88450 580758
rect 79869 580755 79935 580756
rect 88701 580755 88767 580758
rect 91686 580756 91692 580820
rect 91756 580818 91762 580820
rect 92381 580818 92447 580821
rect 91756 580816 92447 580818
rect 91756 580760 92386 580816
rect 92442 580760 92447 580816
rect 91756 580758 92447 580760
rect 91756 580756 91762 580758
rect 92381 580755 92447 580758
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 65977 580002 66043 580005
rect 68878 580002 68938 580584
rect 65977 580000 68938 580002
rect 65977 579944 65982 580000
rect 66038 579944 68938 580000
rect 65977 579942 68938 579944
rect 65977 579939 66043 579942
rect 67173 578642 67239 578645
rect 68878 578642 68938 579224
rect 94638 578914 94698 579496
rect 97165 578914 97231 578917
rect 94638 578912 97231 578914
rect 94638 578856 97170 578912
rect 97226 578856 97231 578912
rect 94638 578854 97231 578856
rect 97165 578851 97231 578854
rect 67173 578640 68938 578642
rect 67173 578584 67178 578640
rect 67234 578584 68938 578640
rect 67173 578582 68938 578584
rect 67173 578579 67239 578582
rect 67449 577282 67515 577285
rect 68878 577282 68938 577864
rect 94638 577554 94698 578136
rect 582741 577690 582807 577693
rect 583520 577690 584960 577780
rect 582741 577688 584960 577690
rect 582741 577632 582746 577688
rect 582802 577632 584960 577688
rect 582741 577630 584960 577632
rect 582741 577627 582807 577630
rect 97901 577554 97967 577557
rect 94638 577552 97967 577554
rect 94638 577496 97906 577552
rect 97962 577496 97967 577552
rect 583520 577540 584960 577630
rect 94638 577494 97967 577496
rect 97901 577491 97967 577494
rect 67449 577280 68938 577282
rect 67449 577224 67454 577280
rect 67510 577224 68938 577280
rect 67449 577222 68938 577224
rect 67449 577219 67515 577222
rect 94638 576738 94698 576776
rect 97901 576738 97967 576741
rect 94638 576736 97967 576738
rect 94638 576680 97906 576736
rect 97962 576680 97967 576736
rect 94638 576678 97967 576680
rect 97901 576675 97967 576678
rect 67725 575922 67791 575925
rect 68878 575922 68938 576504
rect 67725 575920 68938 575922
rect 67725 575864 67730 575920
rect 67786 575864 68938 575920
rect 67725 575862 68938 575864
rect 67725 575859 67791 575862
rect 67541 575378 67607 575381
rect 67541 575376 68938 575378
rect 67541 575320 67546 575376
rect 67602 575320 68938 575376
rect 67541 575318 68938 575320
rect 67541 575315 67607 575318
rect 68878 575144 68938 575318
rect 94638 574834 94698 575416
rect 95233 574834 95299 574837
rect 94638 574832 95299 574834
rect 94638 574776 95238 574832
rect 95294 574776 95299 574832
rect 94638 574774 95299 574776
rect 95233 574771 95299 574774
rect 66713 573202 66779 573205
rect 68878 573202 68938 573784
rect 94638 573474 94698 574056
rect 96981 573474 97047 573477
rect 94638 573472 97047 573474
rect 94638 573416 96986 573472
rect 97042 573416 97047 573472
rect 94638 573414 97047 573416
rect 96981 573411 97047 573414
rect 66713 573200 68938 573202
rect 66713 573144 66718 573200
rect 66774 573144 68938 573200
rect 66713 573142 68938 573144
rect 66713 573139 66779 573142
rect 66805 571842 66871 571845
rect 68878 571842 68938 572424
rect 94638 572114 94698 572696
rect 97533 572114 97599 572117
rect 94638 572112 97599 572114
rect 94638 572056 97538 572112
rect 97594 572056 97599 572112
rect 94638 572054 97599 572056
rect 97533 572051 97599 572054
rect 66805 571840 68938 571842
rect 66805 571784 66810 571840
rect 66866 571784 68938 571840
rect 66805 571782 68938 571784
rect 66805 571779 66871 571782
rect 104934 571434 104940 571436
rect 94638 571374 104940 571434
rect 94638 571336 94698 571374
rect 104934 571372 104940 571374
rect 105004 571372 105010 571436
rect 66897 570210 66963 570213
rect 68878 570210 68938 570792
rect 66897 570208 68938 570210
rect 66897 570152 66902 570208
rect 66958 570152 68938 570208
rect 66897 570150 68938 570152
rect 66897 570147 66963 570150
rect 97901 570074 97967 570077
rect 94638 570072 97967 570074
rect 94638 570016 97906 570072
rect 97962 570016 97967 570072
rect 94638 570014 97967 570016
rect 94638 569976 94698 570014
rect 97901 570011 97967 570014
rect 66529 568986 66595 568989
rect 68878 568986 68938 569432
rect 97257 569258 97323 569261
rect 66529 568984 68938 568986
rect 66529 568928 66534 568984
rect 66590 568928 68938 568984
rect 66529 568926 68938 568928
rect 94638 569256 97323 569258
rect 94638 569200 97262 569256
rect 97318 569200 97323 569256
rect 94638 569198 97323 569200
rect 66529 568923 66595 568926
rect 94638 568616 94698 569198
rect 97257 569195 97323 569198
rect 99373 569258 99439 569261
rect 115054 569258 115060 569260
rect 99373 569256 115060 569258
rect 99373 569200 99378 569256
rect 99434 569200 115060 569256
rect 99373 569198 115060 569200
rect 99373 569195 99439 569198
rect 115054 569196 115060 569198
rect 115124 569196 115130 569260
rect 65885 567626 65951 567629
rect 68878 567626 68938 568072
rect 65885 567624 68938 567626
rect 65885 567568 65890 567624
rect 65946 567568 68938 567624
rect 65885 567566 68938 567568
rect 65885 567563 65951 567566
rect 94638 567218 94698 567256
rect 95325 567218 95391 567221
rect 94638 567216 95391 567218
rect 94638 567160 95330 567216
rect 95386 567160 95391 567216
rect 94638 567158 95391 567160
rect 95325 567155 95391 567158
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67633 566674 67699 566677
rect 68878 566674 68938 566712
rect 67633 566672 68938 566674
rect 67633 566616 67638 566672
rect 67694 566616 68938 566672
rect 67633 566614 68938 566616
rect 67633 566611 67699 566614
rect 94638 565858 94698 565896
rect 96705 565858 96771 565861
rect 94638 565856 96771 565858
rect 94638 565800 96710 565856
rect 96766 565800 96771 565856
rect 94638 565798 96771 565800
rect 96705 565795 96771 565798
rect 66897 564770 66963 564773
rect 68878 564770 68938 565352
rect 66897 564768 68938 564770
rect 66897 564712 66902 564768
rect 66958 564712 68938 564768
rect 66897 564710 68938 564712
rect 66897 564707 66963 564710
rect 583017 564362 583083 564365
rect 583520 564362 584960 564452
rect 583017 564360 584960 564362
rect 583017 564304 583022 564360
rect 583078 564304 584960 564360
rect 583017 564302 584960 564304
rect 583017 564299 583083 564302
rect 66897 563410 66963 563413
rect 68878 563410 68938 563992
rect 94638 563685 94698 564264
rect 583520 564212 584960 564302
rect 94638 563680 94747 563685
rect 94638 563624 94686 563680
rect 94742 563624 94747 563680
rect 94638 563622 94747 563624
rect 94681 563619 94747 563622
rect 66897 563408 68938 563410
rect 66897 563352 66902 563408
rect 66958 563352 68938 563408
rect 66897 563350 68938 563352
rect 66897 563347 66963 563350
rect 66161 562050 66227 562053
rect 68878 562050 68938 562632
rect 94638 562322 94698 562904
rect 96797 562322 96863 562325
rect 94638 562320 96863 562322
rect 94638 562264 96802 562320
rect 96858 562264 96863 562320
rect 94638 562262 96863 562264
rect 96797 562259 96863 562262
rect 66161 562048 68938 562050
rect 66161 561992 66166 562048
rect 66222 561992 68938 562048
rect 66161 561990 68938 561992
rect 66161 561987 66227 561990
rect 66805 560690 66871 560693
rect 68878 560690 68938 561272
rect 94638 560962 94698 561544
rect 96797 560962 96863 560965
rect 94638 560960 96863 560962
rect 94638 560904 96802 560960
rect 96858 560904 96863 560960
rect 94638 560902 96863 560904
rect 96797 560899 96863 560902
rect 66805 560688 68938 560690
rect 66805 560632 66810 560688
rect 66866 560632 68938 560688
rect 66805 560630 68938 560632
rect 66805 560627 66871 560630
rect 66805 559330 66871 559333
rect 68878 559330 68938 559912
rect 94638 559602 94698 560184
rect 97073 559602 97139 559605
rect 94638 559600 97139 559602
rect 94638 559544 97078 559600
rect 97134 559544 97139 559600
rect 94638 559542 97139 559544
rect 97073 559539 97139 559542
rect 66805 559328 68938 559330
rect 66805 559272 66810 559328
rect 66866 559272 68938 559328
rect 66805 559270 68938 559272
rect 66805 559267 66871 559270
rect 94638 558786 94698 558824
rect 96889 558786 96955 558789
rect 97901 558786 97967 558789
rect 94638 558784 97967 558786
rect 94638 558728 96894 558784
rect 96950 558728 97906 558784
rect 97962 558728 97967 558784
rect 94638 558726 97967 558728
rect 96889 558723 96955 558726
rect 97901 558723 97967 558726
rect 66805 557970 66871 557973
rect 68878 557970 68938 558552
rect 66805 557968 68938 557970
rect 66805 557912 66810 557968
rect 66866 557912 68938 557968
rect 66805 557910 68938 557912
rect 66805 557907 66871 557910
rect 67817 556610 67883 556613
rect 68878 556610 68938 557192
rect 94638 556882 94698 557464
rect 96613 556882 96679 556885
rect 94638 556880 96679 556882
rect 94638 556824 96618 556880
rect 96674 556824 96679 556880
rect 94638 556822 96679 556824
rect 96613 556819 96679 556822
rect 67817 556608 68938 556610
rect 67817 556552 67822 556608
rect 67878 556552 68938 556608
rect 67817 556550 68938 556552
rect 67817 556547 67883 556550
rect 67357 555250 67423 555253
rect 68878 555250 68938 555832
rect 94638 555522 94698 556104
rect 96705 555522 96771 555525
rect 94638 555520 96771 555522
rect 94638 555464 96710 555520
rect 96766 555464 96771 555520
rect 94638 555462 96771 555464
rect 96705 555459 96771 555462
rect 67357 555248 68938 555250
rect 67357 555192 67362 555248
rect 67418 555192 68938 555248
rect 67357 555190 68938 555192
rect 67357 555187 67423 555190
rect -960 553890 480 553980
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 66897 553618 66963 553621
rect 68878 553618 68938 554200
rect 94638 554162 94698 554744
rect 96889 554162 96955 554165
rect 94638 554160 96955 554162
rect 94638 554104 96894 554160
rect 96950 554104 96955 554160
rect 94638 554102 96955 554104
rect 96889 554099 96955 554102
rect 66897 553616 68938 553618
rect 66897 553560 66902 553616
rect 66958 553560 68938 553616
rect 66897 553558 68938 553560
rect 66897 553555 66963 553558
rect 67265 552258 67331 552261
rect 68878 552258 68938 552840
rect 94638 552802 94698 553384
rect 96981 552802 97047 552805
rect 94638 552800 97047 552802
rect 94638 552744 96986 552800
rect 97042 552744 97047 552800
rect 94638 552742 97047 552744
rect 96981 552739 97047 552742
rect 95417 552530 95483 552533
rect 97073 552530 97139 552533
rect 67265 552256 68938 552258
rect 67265 552200 67270 552256
rect 67326 552200 68938 552256
rect 67265 552198 68938 552200
rect 94638 552528 97139 552530
rect 94638 552472 95422 552528
rect 95478 552472 97078 552528
rect 97134 552472 97139 552528
rect 94638 552470 97139 552472
rect 67265 552195 67331 552198
rect 94638 552024 94698 552470
rect 95417 552467 95483 552470
rect 97073 552467 97139 552470
rect 69430 550900 69490 551480
rect 583520 551020 584960 551260
rect 69422 550836 69428 550900
rect 69492 550836 69498 550900
rect 115974 550762 115980 550764
rect 94638 550702 115980 550762
rect 94638 550664 94698 550702
rect 115974 550700 115980 550702
rect 116044 550700 116050 550764
rect 66713 549538 66779 549541
rect 68878 549538 68938 550120
rect 66713 549536 68938 549538
rect 66713 549480 66718 549536
rect 66774 549480 68938 549536
rect 66713 549478 68938 549480
rect 66713 549475 66779 549478
rect 97441 549402 97507 549405
rect 94638 549400 97507 549402
rect 94638 549344 97446 549400
rect 97502 549344 97507 549400
rect 94638 549342 97507 549344
rect 94638 549304 94698 549342
rect 97441 549339 97507 549342
rect 68645 548314 68711 548317
rect 68878 548314 68938 548760
rect 68645 548312 68938 548314
rect 68645 548256 68650 548312
rect 68706 548256 68938 548312
rect 68645 548254 68938 548256
rect 68645 548251 68711 548254
rect 66805 546818 66871 546821
rect 68878 546818 68938 547400
rect 94638 547090 94698 547672
rect 96654 547090 96660 547092
rect 94638 547030 96660 547090
rect 96654 547028 96660 547030
rect 96724 547028 96730 547092
rect 66805 546816 68938 546818
rect 66805 546760 66810 546816
rect 66866 546760 68938 546816
rect 66805 546758 68938 546760
rect 66805 546755 66871 546758
rect 66805 545458 66871 545461
rect 68878 545458 68938 546040
rect 94638 545730 94698 546312
rect 96705 545730 96771 545733
rect 94638 545728 96771 545730
rect 94638 545672 96710 545728
rect 96766 545672 96771 545728
rect 94638 545670 96771 545672
rect 96705 545667 96771 545670
rect 66805 545456 68938 545458
rect 66805 545400 66810 545456
rect 66866 545400 68938 545456
rect 66805 545398 68938 545400
rect 66805 545395 66871 545398
rect 66069 544098 66135 544101
rect 68878 544098 68938 544680
rect 94638 544370 94698 544952
rect 97073 544370 97139 544373
rect 94638 544368 97139 544370
rect 94638 544312 97078 544368
rect 97134 544312 97139 544368
rect 94638 544310 97139 544312
rect 97073 544307 97139 544310
rect 66069 544096 68938 544098
rect 66069 544040 66074 544096
rect 66130 544040 68938 544096
rect 66069 544038 68938 544040
rect 66069 544035 66135 544038
rect 68645 543554 68711 543557
rect 69422 543554 69428 543556
rect 68645 543552 69428 543554
rect 68645 543496 68650 543552
rect 68706 543496 69428 543552
rect 68645 543494 69428 543496
rect 68645 543491 68711 543494
rect 69422 543492 69428 543494
rect 69492 543492 69498 543556
rect 68369 543350 68435 543353
rect 68369 543348 68908 543350
rect 68369 543292 68374 543348
rect 68430 543292 68908 543348
rect 68369 543290 68908 543292
rect 68369 543287 68435 543290
rect 94638 543010 94698 543592
rect 97073 543010 97139 543013
rect 94638 543008 97139 543010
rect 94638 542952 97078 543008
rect 97134 542952 97139 543008
rect 94638 542950 97139 542952
rect 97073 542947 97139 542950
rect 66621 541378 66687 541381
rect 68878 541378 68938 541960
rect 94638 541650 94698 542232
rect 96613 541650 96679 541653
rect 94638 541648 96679 541650
rect 94638 541592 96618 541648
rect 96674 541592 96679 541648
rect 94638 541590 96679 541592
rect 96613 541587 96679 541590
rect 66621 541376 68938 541378
rect 66621 541320 66626 541376
rect 66682 541320 68938 541376
rect 66621 541318 68938 541320
rect 66621 541315 66687 541318
rect -960 540684 480 540924
rect 69430 539882 69490 540600
rect 69430 539822 69674 539882
rect 69614 539746 69674 539822
rect 94270 539749 94330 540872
rect 70301 539746 70367 539749
rect 69614 539744 70367 539746
rect 69614 539688 70306 539744
rect 70362 539688 70367 539744
rect 69614 539686 70367 539688
rect 94270 539744 94379 539749
rect 94270 539688 94318 539744
rect 94374 539688 94379 539744
rect 94270 539686 94379 539688
rect 70301 539683 70367 539686
rect 94313 539683 94379 539686
rect 75862 539548 75868 539612
rect 75932 539610 75938 539612
rect 76741 539610 76807 539613
rect 75932 539608 76807 539610
rect 75932 539552 76746 539608
rect 76802 539552 76807 539608
rect 75932 539550 76807 539552
rect 75932 539548 75938 539550
rect 76741 539547 76807 539550
rect 93945 538930 94011 538933
rect 94086 538930 94146 539512
rect 93945 538928 94146 538930
rect 93945 538872 93950 538928
rect 94006 538872 94146 538928
rect 93945 538870 94146 538872
rect 93945 538867 94011 538870
rect 65885 538794 65951 538797
rect 142153 538794 142219 538797
rect 65885 538792 142219 538794
rect 65885 538736 65890 538792
rect 65946 538736 142158 538792
rect 142214 538736 142219 538792
rect 65885 538734 142219 538736
rect 65885 538731 65951 538734
rect 142153 538731 142219 538734
rect 583109 537842 583175 537845
rect 583520 537842 584960 537932
rect 583109 537840 584960 537842
rect 583109 537784 583114 537840
rect 583170 537784 584960 537840
rect 583109 537782 584960 537784
rect 583109 537779 583175 537782
rect 583520 537692 584960 537782
rect 73286 537508 73292 537572
rect 73356 537570 73362 537572
rect 91686 537570 91692 537572
rect 73356 537510 91692 537570
rect 73356 537508 73362 537510
rect 91686 537508 91692 537510
rect 91756 537508 91762 537572
rect 69790 537372 69796 537436
rect 69860 537434 69866 537436
rect 115197 537434 115263 537437
rect 69860 537432 115263 537434
rect 69860 537376 115202 537432
rect 115258 537376 115263 537432
rect 69860 537374 115263 537376
rect 69860 537372 69866 537374
rect 115197 537371 115263 537374
rect 90357 536754 90423 536757
rect 136633 536754 136699 536757
rect 90357 536752 136699 536754
rect 90357 536696 90362 536752
rect 90418 536696 136638 536752
rect 136694 536696 136699 536752
rect 90357 536694 136699 536696
rect 90357 536691 90423 536694
rect 136633 536691 136699 536694
rect 88425 534850 88491 534853
rect 106406 534850 106412 534852
rect 88425 534848 106412 534850
rect 88425 534792 88430 534848
rect 88486 534792 106412 534848
rect 88425 534790 106412 534792
rect 88425 534787 88491 534790
rect 106406 534788 106412 534790
rect 106476 534788 106482 534852
rect 61837 534714 61903 534717
rect 96654 534714 96660 534716
rect 61837 534712 96660 534714
rect 61837 534656 61842 534712
rect 61898 534656 96660 534712
rect 61837 534654 96660 534656
rect 61837 534651 61903 534654
rect 96654 534652 96660 534654
rect 96724 534652 96730 534716
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 582925 524514 582991 524517
rect 583520 524514 584960 524604
rect 582925 524512 584960 524514
rect 582925 524456 582930 524512
rect 582986 524456 584960 524512
rect 582925 524454 584960 524456
rect 582925 524451 582991 524454
rect 583520 524364 584960 524454
rect 79726 523636 79732 523700
rect 79796 523698 79802 523700
rect 95325 523698 95391 523701
rect 79796 523696 95391 523698
rect 79796 523640 95330 523696
rect 95386 523640 95391 523696
rect 79796 523638 95391 523640
rect 79796 523636 79802 523638
rect 95325 523635 95391 523638
rect 72734 520916 72740 520980
rect 72804 520978 72810 520980
rect 94681 520978 94747 520981
rect 72804 520976 94747 520978
rect 72804 520920 94686 520976
rect 94742 520920 94747 520976
rect 72804 520918 94747 520920
rect 72804 520916 72810 520918
rect 94681 520915 94747 520918
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 583293 511322 583359 511325
rect 583520 511322 584960 511412
rect 583293 511320 584960 511322
rect 583293 511264 583298 511320
rect 583354 511264 584960 511320
rect 583293 511262 584960 511264
rect 583293 511259 583359 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 67725 479498 67791 479501
rect 96654 479498 96660 479500
rect 67725 479496 96660 479498
rect 67725 479440 67730 479496
rect 67786 479440 96660 479496
rect 67725 479438 96660 479440
rect 67725 479435 67791 479438
rect 96654 479436 96660 479438
rect 96724 479436 96730 479500
rect 75678 476716 75684 476780
rect 75748 476778 75754 476780
rect 90909 476778 90975 476781
rect 75748 476776 90975 476778
rect 75748 476720 90914 476776
rect 90970 476720 90975 476776
rect 75748 476718 90975 476720
rect 75748 476716 75754 476718
rect 90909 476715 90975 476718
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 81433 472562 81499 472565
rect 107694 472562 107700 472564
rect 81433 472560 107700 472562
rect 81433 472504 81438 472560
rect 81494 472504 107700 472560
rect 81433 472502 107700 472504
rect 81433 472499 81499 472502
rect 107694 472500 107700 472502
rect 107764 472500 107770 472564
rect 583201 471474 583267 471477
rect 583520 471474 584960 471564
rect 583201 471472 584960 471474
rect 583201 471416 583206 471472
rect 583262 471416 584960 471472
rect 583201 471414 584960 471416
rect 583201 471411 583267 471414
rect 583520 471324 584960 471414
rect 67766 468420 67772 468484
rect 67836 468482 67842 468484
rect 96705 468482 96771 468485
rect 67836 468480 96771 468482
rect 67836 468424 96710 468480
rect 96766 468424 96771 468480
rect 67836 468422 96771 468424
rect 67836 468420 67842 468422
rect 96705 468419 96771 468422
rect 69657 466580 69723 466581
rect 69606 466578 69612 466580
rect 69566 466518 69612 466578
rect 69676 466578 69723 466580
rect 194593 466578 194659 466581
rect 69676 466576 194659 466578
rect 69718 466520 194598 466576
rect 194654 466520 194659 466576
rect 69606 466516 69612 466518
rect 69676 466518 194659 466520
rect 69676 466516 69723 466518
rect 69657 466515 69723 466516
rect 194593 466515 194659 466518
rect 120717 465218 120783 465221
rect 259637 465218 259703 465221
rect 120717 465216 259703 465218
rect 120717 465160 120722 465216
rect 120778 465160 259642 465216
rect 259698 465160 259703 465216
rect 120717 465158 259703 465160
rect 120717 465155 120783 465158
rect 259637 465155 259703 465158
rect 72918 464340 72924 464404
rect 72988 464402 72994 464404
rect 113214 464402 113220 464404
rect 72988 464342 113220 464402
rect 72988 464340 72994 464342
rect 113214 464340 113220 464342
rect 113284 464340 113290 464404
rect 109677 463586 109743 463589
rect 110321 463586 110387 463589
rect 109677 463584 110387 463586
rect 109677 463528 109682 463584
rect 109738 463528 110326 463584
rect 110382 463528 110387 463584
rect 109677 463526 110387 463528
rect 109677 463523 109743 463526
rect 110321 463523 110387 463526
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 110321 462362 110387 462365
rect 262254 462362 262260 462364
rect 110321 462360 262260 462362
rect 110321 462304 110326 462360
rect 110382 462304 262260 462360
rect 110321 462302 262260 462304
rect 110321 462299 110387 462302
rect 262254 462300 262260 462302
rect 262324 462300 262330 462364
rect 88333 461546 88399 461549
rect 118693 461546 118759 461549
rect 88333 461544 118759 461546
rect 88333 461488 88338 461544
rect 88394 461488 118698 461544
rect 118754 461488 118759 461544
rect 88333 461486 118759 461488
rect 88333 461483 88399 461486
rect 118693 461483 118759 461486
rect 118693 461002 118759 461005
rect 253933 461002 253999 461005
rect 118693 461000 253999 461002
rect 118693 460944 118698 461000
rect 118754 460944 253938 461000
rect 253994 460944 253999 461000
rect 118693 460942 253999 460944
rect 118693 460939 118759 460942
rect 253933 460939 253999 460942
rect 83406 460124 83412 460188
rect 83476 460186 83482 460188
rect 97206 460186 97212 460188
rect 83476 460126 97212 460186
rect 83476 460124 83482 460126
rect 97206 460124 97212 460126
rect 97276 460124 97282 460188
rect 240133 460186 240199 460189
rect 280153 460186 280219 460189
rect 240133 460184 280219 460186
rect 240133 460128 240138 460184
rect 240194 460128 280158 460184
rect 280214 460128 280219 460184
rect 240133 460126 280219 460128
rect 240133 460123 240199 460126
rect 280153 460123 280219 460126
rect 75913 459642 75979 459645
rect 83590 459642 83596 459644
rect 75913 459640 83596 459642
rect 75913 459584 75918 459640
rect 75974 459584 83596 459640
rect 75913 459582 83596 459584
rect 75913 459579 75979 459582
rect 83590 459580 83596 459582
rect 83660 459580 83666 459644
rect 189717 459642 189783 459645
rect 216857 459642 216923 459645
rect 220077 459642 220143 459645
rect 189717 459640 220143 459642
rect 189717 459584 189722 459640
rect 189778 459584 216862 459640
rect 216918 459584 220082 459640
rect 220138 459584 220143 459640
rect 189717 459582 220143 459584
rect 189717 459579 189783 459582
rect 216857 459579 216923 459582
rect 220077 459579 220143 459582
rect 238753 459642 238819 459645
rect 240133 459642 240199 459645
rect 238753 459640 240199 459642
rect 238753 459584 238758 459640
rect 238814 459584 240138 459640
rect 240194 459584 240199 459640
rect 238753 459582 240199 459584
rect 238753 459579 238819 459582
rect 240133 459579 240199 459582
rect 76557 458826 76623 458829
rect 99966 458826 99972 458828
rect 76557 458824 99972 458826
rect 76557 458768 76562 458824
rect 76618 458768 99972 458824
rect 76557 458766 99972 458768
rect 76557 458763 76623 458766
rect 99966 458764 99972 458766
rect 100036 458764 100042 458828
rect 179229 458418 179295 458421
rect 210417 458418 210483 458421
rect 179229 458416 210483 458418
rect 179229 458360 179234 458416
rect 179290 458360 210422 458416
rect 210478 458360 210483 458416
rect 179229 458358 210483 458360
rect 179229 458355 179295 458358
rect 210417 458355 210483 458358
rect 195789 458284 195855 458285
rect 195789 458280 195836 458284
rect 195900 458282 195906 458284
rect 249241 458282 249307 458285
rect 284293 458282 284359 458285
rect 195789 458224 195794 458280
rect 195789 458220 195836 458224
rect 195900 458222 195946 458282
rect 249241 458280 284359 458282
rect 249241 458224 249246 458280
rect 249302 458224 284298 458280
rect 284354 458224 284359 458280
rect 249241 458222 284359 458224
rect 195900 458220 195906 458222
rect 195789 458219 195855 458220
rect 249241 458219 249307 458222
rect 284293 458219 284359 458222
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 173801 457058 173867 457061
rect 207565 457058 207631 457061
rect 173801 457056 207631 457058
rect 173801 457000 173806 457056
rect 173862 457000 207570 457056
rect 207626 457000 207631 457056
rect 173801 456998 207631 457000
rect 173801 456995 173867 456998
rect 207565 456995 207631 456998
rect 219801 457058 219867 457061
rect 247718 457058 247724 457060
rect 219801 457056 247724 457058
rect 219801 457000 219806 457056
rect 219862 457000 247724 457056
rect 219801 456998 247724 457000
rect 219801 456995 219867 456998
rect 247718 456996 247724 456998
rect 247788 456996 247794 457060
rect 116577 456922 116643 456925
rect 250621 456922 250687 456925
rect 116577 456920 250687 456922
rect 116577 456864 116582 456920
rect 116638 456864 250626 456920
rect 250682 456864 250687 456920
rect 116577 456862 250687 456864
rect 116577 456859 116643 456862
rect 250621 456859 250687 456862
rect 582649 456106 582715 456109
rect 287010 456104 582715 456106
rect 287010 456048 582654 456104
rect 582710 456048 582715 456104
rect 287010 456046 582715 456048
rect 192661 455698 192727 455701
rect 212717 455698 212783 455701
rect 192661 455696 212783 455698
rect 192661 455640 192666 455696
rect 192722 455640 212722 455696
rect 212778 455640 212783 455696
rect 192661 455638 212783 455640
rect 192661 455635 192727 455638
rect 212717 455635 212783 455638
rect 233233 455698 233299 455701
rect 252686 455698 252692 455700
rect 233233 455696 252692 455698
rect 233233 455640 233238 455696
rect 233294 455640 252692 455696
rect 233233 455638 252692 455640
rect 233233 455635 233299 455638
rect 252686 455636 252692 455638
rect 252756 455636 252762 455700
rect 187601 455562 187667 455565
rect 214557 455562 214623 455565
rect 187601 455560 214623 455562
rect 187601 455504 187606 455560
rect 187662 455504 214562 455560
rect 214618 455504 214623 455560
rect 187601 455502 214623 455504
rect 187601 455499 187667 455502
rect 214557 455499 214623 455502
rect 220813 455562 220879 455565
rect 284334 455562 284340 455564
rect 220813 455560 284340 455562
rect 220813 455504 220818 455560
rect 220874 455504 284340 455560
rect 220813 455502 284340 455504
rect 220813 455499 220879 455502
rect 284334 455500 284340 455502
rect 284404 455562 284410 455564
rect 287010 455562 287070 456046
rect 582649 456043 582715 456046
rect 284404 455502 287070 455562
rect 284404 455500 284410 455502
rect 180149 454474 180215 454477
rect 255497 454474 255563 454477
rect 180149 454472 255563 454474
rect 180149 454416 180154 454472
rect 180210 454416 255502 454472
rect 255558 454416 255563 454472
rect 180149 454414 255563 454416
rect 180149 454411 180215 454414
rect 255497 454411 255563 454414
rect 176653 454338 176719 454341
rect 177941 454338 178007 454341
rect 207105 454338 207171 454341
rect 176653 454336 207171 454338
rect 176653 454280 176658 454336
rect 176714 454280 177946 454336
rect 178002 454280 207110 454336
rect 207166 454280 207171 454336
rect 176653 454278 207171 454280
rect 176653 454275 176719 454278
rect 177941 454275 178007 454278
rect 207105 454275 207171 454278
rect 147581 454202 147647 454205
rect 197905 454202 197971 454205
rect 147581 454200 197971 454202
rect 147581 454144 147586 454200
rect 147642 454144 197910 454200
rect 197966 454144 197971 454200
rect 147581 454142 197971 454144
rect 147581 454139 147647 454142
rect 197905 454139 197971 454142
rect 231209 454202 231275 454205
rect 276238 454202 276244 454204
rect 231209 454200 276244 454202
rect 231209 454144 231214 454200
rect 231270 454144 276244 454200
rect 231209 454142 276244 454144
rect 231209 454139 231275 454142
rect 276238 454140 276244 454142
rect 276308 454140 276314 454204
rect 77385 454066 77451 454069
rect 176653 454066 176719 454069
rect 77385 454064 176719 454066
rect 77385 454008 77390 454064
rect 77446 454008 176658 454064
rect 176714 454008 176719 454064
rect 77385 454006 176719 454008
rect 77385 454003 77451 454006
rect 176653 454003 176719 454006
rect 234889 454066 234955 454069
rect 244774 454066 244780 454068
rect 234889 454064 244780 454066
rect 234889 454008 234894 454064
rect 234950 454008 244780 454064
rect 234889 454006 244780 454008
rect 234889 454003 234955 454006
rect 244774 454004 244780 454006
rect 244844 454004 244850 454068
rect 242157 453930 242223 453933
rect 243997 453930 244063 453933
rect 242157 453928 244063 453930
rect 242157 453872 242162 453928
rect 242218 453872 244002 453928
rect 244058 453872 244063 453928
rect 242157 453870 244063 453872
rect 242157 453867 242223 453870
rect 243997 453867 244063 453870
rect 225045 453250 225111 453253
rect 237373 453250 237439 453253
rect 225045 453248 237439 453250
rect 225045 453192 225050 453248
rect 225106 453192 237378 453248
rect 237434 453192 237439 453248
rect 225045 453190 237439 453192
rect 225045 453187 225111 453190
rect 237373 453187 237439 453190
rect 71037 453114 71103 453117
rect 194685 453114 194751 453117
rect 71037 453112 194751 453114
rect 71037 453056 71042 453112
rect 71098 453056 194690 453112
rect 194746 453056 194751 453112
rect 71037 453054 194751 453056
rect 71037 453051 71103 453054
rect 194685 453051 194751 453054
rect 197118 453052 197124 453116
rect 197188 453114 197194 453116
rect 203149 453114 203215 453117
rect 197188 453112 203215 453114
rect 197188 453056 203154 453112
rect 203210 453056 203215 453112
rect 197188 453054 203215 453056
rect 197188 453052 197194 453054
rect 203149 453051 203215 453054
rect 183461 452978 183527 452981
rect 195973 452978 196039 452981
rect 183461 452976 196039 452978
rect 183461 452920 183466 452976
rect 183522 452920 195978 452976
rect 196034 452920 196039 452976
rect 183461 452918 196039 452920
rect 183461 452915 183527 452918
rect 195973 452915 196039 452918
rect 243997 452978 244063 452981
rect 263593 452978 263659 452981
rect 243997 452976 263659 452978
rect 243997 452920 244002 452976
rect 244058 452920 263598 452976
rect 263654 452920 263659 452976
rect 243997 452918 263659 452920
rect 243997 452915 244063 452918
rect 263593 452915 263659 452918
rect 187509 452842 187575 452845
rect 205909 452842 205975 452845
rect 187509 452840 205975 452842
rect 187509 452784 187514 452840
rect 187570 452784 205914 452840
rect 205970 452784 205975 452840
rect 187509 452782 205975 452784
rect 187509 452779 187575 452782
rect 205909 452779 205975 452782
rect 212441 452706 212507 452709
rect 224125 452706 224191 452709
rect 212441 452704 224191 452706
rect 212441 452648 212446 452704
rect 212502 452648 224130 452704
rect 224186 452648 224191 452704
rect 212441 452646 224191 452648
rect 212441 452643 212507 452646
rect 224125 452643 224191 452646
rect 234429 452706 234495 452709
rect 242014 452706 242020 452708
rect 234429 452704 242020 452706
rect 234429 452648 234434 452704
rect 234490 452648 242020 452704
rect 234429 452646 242020 452648
rect 234429 452643 234495 452646
rect 242014 452644 242020 452646
rect 242084 452644 242090 452708
rect 250621 452706 250687 452709
rect 254526 452706 254532 452708
rect 250621 452704 254532 452706
rect 250621 452648 250626 452704
rect 250682 452648 254532 452704
rect 250621 452646 254532 452648
rect 250621 452643 250687 452646
rect 254526 452644 254532 452646
rect 254596 452644 254602 452708
rect 124121 451890 124187 451893
rect 211613 451890 211679 451893
rect 124121 451888 211679 451890
rect 124121 451832 124126 451888
rect 124182 451832 211618 451888
rect 211674 451832 211679 451888
rect 124121 451830 211679 451832
rect 124121 451827 124187 451830
rect 211613 451827 211679 451830
rect 236729 451890 236795 451893
rect 298093 451890 298159 451893
rect 236729 451888 298159 451890
rect 236729 451832 236734 451888
rect 236790 451832 298098 451888
rect 298154 451832 298159 451888
rect 236729 451830 298159 451832
rect 236729 451827 236795 451830
rect 298093 451827 298159 451830
rect 191097 451482 191163 451485
rect 209773 451482 209839 451485
rect 191097 451480 209839 451482
rect 191097 451424 191102 451480
rect 191158 451424 209778 451480
rect 209834 451424 209839 451480
rect 191097 451422 209839 451424
rect 191097 451419 191163 451422
rect 209773 451419 209839 451422
rect 122097 451346 122163 451349
rect 247861 451346 247927 451349
rect 122097 451344 247927 451346
rect 122097 451288 122102 451344
rect 122158 451288 247866 451344
rect 247922 451288 247927 451344
rect 122097 451286 247927 451288
rect 122097 451283 122163 451286
rect 247861 451283 247927 451286
rect 228081 450394 228147 450397
rect 277393 450394 277459 450397
rect 228081 450392 277459 450394
rect 228081 450336 228086 450392
rect 228142 450336 277398 450392
rect 277454 450336 277459 450392
rect 228081 450334 277459 450336
rect 228081 450331 228147 450334
rect 277393 450331 277459 450334
rect 187141 450258 187207 450261
rect 230473 450258 230539 450261
rect 187141 450256 230539 450258
rect 187141 450200 187146 450256
rect 187202 450200 230478 450256
rect 230534 450200 230539 450256
rect 187141 450198 230539 450200
rect 187141 450195 187207 450198
rect 230473 450195 230539 450198
rect 133137 450122 133203 450125
rect 244549 450122 244615 450125
rect 255957 450122 256023 450125
rect 133137 450120 256023 450122
rect 133137 450064 133142 450120
rect 133198 450064 244554 450120
rect 244610 450064 255962 450120
rect 256018 450064 256023 450120
rect 133137 450062 256023 450064
rect 133137 450059 133203 450062
rect 244549 450059 244615 450062
rect 255957 450059 256023 450062
rect 86217 449986 86283 449989
rect 88374 449986 88380 449988
rect 86217 449984 88380 449986
rect 86217 449928 86222 449984
rect 86278 449928 88380 449984
rect 86217 449926 88380 449928
rect 86217 449923 86283 449926
rect 88374 449924 88380 449926
rect 88444 449924 88450 449988
rect 88517 449986 88583 449989
rect 220813 449986 220879 449989
rect 88517 449984 220879 449986
rect 88517 449928 88522 449984
rect 88578 449928 220818 449984
rect 220874 449928 220879 449984
rect 88517 449926 220879 449928
rect 88382 449850 88442 449924
rect 88517 449923 88583 449926
rect 220813 449923 220879 449926
rect 238477 449986 238543 449989
rect 248505 449988 248571 449989
rect 241646 449986 241652 449988
rect 238477 449984 241652 449986
rect 238477 449928 238482 449984
rect 238538 449928 241652 449984
rect 238477 449926 241652 449928
rect 238477 449923 238543 449926
rect 241646 449924 241652 449926
rect 241716 449924 241722 449988
rect 248454 449986 248460 449988
rect 248414 449926 248460 449986
rect 248524 449984 248571 449988
rect 248566 449928 248571 449984
rect 248454 449924 248460 449926
rect 248524 449924 248571 449928
rect 248505 449923 248571 449924
rect 179229 449850 179295 449853
rect 88382 449848 179295 449850
rect 88382 449792 179234 449848
rect 179290 449792 179295 449848
rect 88382 449790 179295 449792
rect 179229 449787 179295 449790
rect 193489 449716 193555 449717
rect 245745 449716 245811 449717
rect 193438 449714 193444 449716
rect -960 449578 480 449668
rect 193398 449654 193444 449714
rect 193508 449712 193555 449716
rect 245694 449714 245700 449716
rect 193550 449656 193555 449712
rect 193438 449652 193444 449654
rect 193508 449652 193555 449656
rect 245654 449654 245700 449714
rect 245764 449712 245811 449716
rect 245806 449656 245811 449712
rect 245694 449652 245700 449654
rect 245764 449652 245811 449656
rect 193489 449651 193555 449652
rect 245745 449651 245811 449652
rect 3233 449578 3299 449581
rect -960 449576 3299 449578
rect -960 449520 3238 449576
rect 3294 449520 3299 449576
rect -960 449518 3299 449520
rect -960 449428 480 449518
rect 3233 449515 3299 449518
rect 191649 449170 191715 449173
rect 191649 449168 193660 449170
rect 191649 449112 191654 449168
rect 191710 449112 193660 449168
rect 191649 449110 193660 449112
rect 191649 449107 191715 449110
rect 255497 448898 255563 448901
rect 253460 448896 255563 448898
rect 253460 448840 255502 448896
rect 255558 448840 255563 448896
rect 253460 448838 255563 448840
rect 255497 448835 255563 448838
rect 100753 448626 100819 448629
rect 101254 448626 101260 448628
rect 100753 448624 101260 448626
rect 100753 448568 100758 448624
rect 100814 448568 101260 448624
rect 100753 448566 101260 448568
rect 100753 448563 100819 448566
rect 101254 448564 101260 448566
rect 101324 448564 101330 448628
rect 179229 448626 179295 448629
rect 180057 448626 180123 448629
rect 179229 448624 180123 448626
rect 179229 448568 179234 448624
rect 179290 448568 180062 448624
rect 180118 448568 180123 448624
rect 179229 448566 180123 448568
rect 179229 448563 179295 448566
rect 180057 448563 180123 448566
rect 117957 448490 118023 448493
rect 187049 448490 187115 448493
rect 117957 448488 187115 448490
rect 117957 448432 117962 448488
rect 118018 448432 187054 448488
rect 187110 448432 187115 448488
rect 117957 448430 187115 448432
rect 117957 448427 118023 448430
rect 187049 448427 187115 448430
rect 182081 447946 182147 447949
rect 192661 447946 192727 447949
rect 182081 447944 192727 447946
rect 182081 447888 182086 447944
rect 182142 447888 192666 447944
rect 192722 447888 192727 447944
rect 182081 447886 192727 447888
rect 182081 447883 182147 447886
rect 192661 447883 192727 447886
rect 191005 447810 191071 447813
rect 191005 447808 193660 447810
rect 191005 447752 191010 447808
rect 191066 447752 193660 447808
rect 191005 447750 193660 447752
rect 191005 447747 191071 447750
rect 255405 447538 255471 447541
rect 253460 447536 255471 447538
rect 253460 447480 255410 447536
rect 255466 447480 255471 447536
rect 253460 447478 255471 447480
rect 255405 447475 255471 447478
rect 66110 446388 66116 446452
rect 66180 446450 66186 446452
rect 86953 446450 87019 446453
rect 66180 446448 87019 446450
rect 66180 446392 86958 446448
rect 87014 446392 87019 446448
rect 66180 446390 87019 446392
rect 66180 446388 66186 446390
rect 86953 446387 87019 446390
rect 191649 446450 191715 446453
rect 191649 446448 193660 446450
rect 191649 446392 191654 446448
rect 191710 446392 193660 446448
rect 191649 446390 193660 446392
rect 191649 446387 191715 446390
rect 253933 446178 253999 446181
rect 254669 446178 254735 446181
rect 253460 446176 254735 446178
rect 253460 446120 253938 446176
rect 253994 446120 254674 446176
rect 254730 446120 254735 446176
rect 253460 446118 254735 446120
rect 253933 446115 253999 446118
rect 254669 446115 254735 446118
rect 69749 445634 69815 445637
rect 70301 445634 70367 445637
rect 193438 445634 193444 445636
rect 69749 445632 193444 445634
rect 69749 445576 69754 445632
rect 69810 445576 70306 445632
rect 70362 445576 193444 445632
rect 69749 445574 193444 445576
rect 69749 445571 69815 445574
rect 70301 445571 70367 445574
rect 193438 445572 193444 445574
rect 193508 445572 193514 445636
rect 193121 445090 193187 445093
rect 193121 445088 193660 445090
rect 193121 445032 193126 445088
rect 193182 445032 193660 445088
rect 193121 445030 193660 445032
rect 193121 445027 193187 445030
rect 255405 444818 255471 444821
rect 253460 444816 255471 444818
rect 253460 444760 255410 444816
rect 255466 444760 255471 444816
rect 253460 444758 255471 444760
rect 255405 444755 255471 444758
rect 583520 444668 584960 444908
rect 69606 442988 69612 443052
rect 69676 443050 69682 443052
rect 193630 443050 193690 443700
rect 255405 443458 255471 443461
rect 253460 443456 255471 443458
rect 253460 443400 255410 443456
rect 255466 443400 255471 443456
rect 253460 443398 255471 443400
rect 255405 443395 255471 443398
rect 69676 442990 193690 443050
rect 69676 442988 69682 442990
rect 110321 442370 110387 442373
rect 117497 442370 117563 442373
rect 110321 442368 117563 442370
rect 110321 442312 110326 442368
rect 110382 442312 117502 442368
rect 117558 442312 117563 442368
rect 110321 442310 117563 442312
rect 110321 442307 110387 442310
rect 117497 442307 117563 442310
rect 50981 442234 51047 442237
rect 95325 442234 95391 442237
rect 50981 442232 95391 442234
rect 50981 442176 50986 442232
rect 51042 442176 95330 442232
rect 95386 442176 95391 442232
rect 50981 442174 95391 442176
rect 50981 442171 51047 442174
rect 95325 442171 95391 442174
rect 100017 442234 100083 442237
rect 114737 442234 114803 442237
rect 100017 442232 114803 442234
rect 100017 442176 100022 442232
rect 100078 442176 114742 442232
rect 114798 442176 114803 442232
rect 100017 442174 114803 442176
rect 100017 442171 100083 442174
rect 114737 442171 114803 442174
rect 191649 442098 191715 442101
rect 255405 442098 255471 442101
rect 191649 442096 193660 442098
rect 191649 442040 191654 442096
rect 191710 442040 193660 442096
rect 191649 442038 193660 442040
rect 253460 442096 255471 442098
rect 253460 442040 255410 442096
rect 255466 442040 255471 442096
rect 253460 442038 255471 442040
rect 191649 442035 191715 442038
rect 255405 442035 255471 442038
rect 122833 441690 122899 441693
rect 191649 441690 191715 441693
rect 122833 441688 191715 441690
rect 122833 441632 122838 441688
rect 122894 441632 191654 441688
rect 191710 441632 191715 441688
rect 122833 441630 191715 441632
rect 122833 441627 122899 441630
rect 191649 441627 191715 441630
rect 21357 441554 21423 441557
rect 104249 441554 104315 441557
rect 21357 441552 104315 441554
rect 21357 441496 21362 441552
rect 21418 441496 104254 441552
rect 104310 441496 104315 441552
rect 21357 441494 104315 441496
rect 21357 441491 21423 441494
rect 104249 441491 104315 441494
rect 191373 440738 191439 440741
rect 191373 440736 193660 440738
rect 191373 440680 191378 440736
rect 191434 440680 193660 440736
rect 191373 440678 193660 440680
rect 191373 440675 191439 440678
rect 253933 440466 253999 440469
rect 253460 440464 253999 440466
rect 253460 440408 253938 440464
rect 253994 440408 253999 440464
rect 253460 440406 253999 440408
rect 253933 440403 253999 440406
rect 66069 439650 66135 439653
rect 82813 439650 82879 439653
rect 66069 439648 82879 439650
rect 66069 439592 66074 439648
rect 66130 439592 82818 439648
rect 82874 439592 82879 439648
rect 66069 439590 82879 439592
rect 66069 439587 66135 439590
rect 82813 439587 82879 439590
rect 83590 439452 83596 439516
rect 83660 439514 83666 439516
rect 184197 439514 184263 439517
rect 83660 439512 184263 439514
rect 83660 439456 184202 439512
rect 184258 439456 184263 439512
rect 83660 439454 184263 439456
rect 83660 439452 83666 439454
rect 184197 439451 184263 439454
rect 191373 439378 191439 439381
rect 191373 439376 193660 439378
rect 191373 439320 191378 439376
rect 191434 439320 193660 439376
rect 191373 439318 193660 439320
rect 191373 439315 191439 439318
rect 255313 439106 255379 439109
rect 253460 439104 255379 439106
rect 253460 439048 255318 439104
rect 255374 439048 255379 439104
rect 253460 439046 255379 439048
rect 255313 439043 255379 439046
rect 98637 438154 98703 438157
rect 107878 438154 107884 438156
rect 98637 438152 107884 438154
rect 98637 438096 98642 438152
rect 98698 438096 107884 438152
rect 98637 438094 107884 438096
rect 98637 438091 98703 438094
rect 107878 438092 107884 438094
rect 107948 438092 107954 438156
rect 191557 438018 191623 438021
rect 191557 438016 193660 438018
rect 191557 437960 191562 438016
rect 191618 437960 193660 438016
rect 191557 437958 193660 437960
rect 191557 437955 191623 437958
rect 255405 437746 255471 437749
rect 253460 437744 255471 437746
rect 253460 437688 255410 437744
rect 255466 437688 255471 437744
rect 253460 437686 255471 437688
rect 255405 437683 255471 437686
rect 133137 437474 133203 437477
rect 122790 437472 133203 437474
rect 122790 437416 133142 437472
rect 133198 437416 133203 437472
rect 122790 437414 133203 437416
rect 106917 437338 106983 437341
rect 122790 437338 122850 437414
rect 133137 437411 133203 437414
rect 106917 437336 122850 437338
rect 106917 437280 106922 437336
rect 106978 437280 122850 437336
rect 106917 437278 122850 437280
rect 106917 437275 106983 437278
rect 110781 437066 110847 437069
rect 116577 437066 116643 437069
rect 110781 437064 116643 437066
rect 110781 437008 110786 437064
rect 110842 437008 116582 437064
rect 116638 437008 116643 437064
rect 110781 437006 116643 437008
rect 110781 437003 110847 437006
rect 116577 437003 116643 437006
rect 113265 436930 113331 436933
rect 262305 436932 262371 436933
rect 263409 436932 263475 436933
rect 114318 436930 114324 436932
rect 113265 436928 114324 436930
rect 113265 436872 113270 436928
rect 113326 436872 114324 436928
rect 113265 436870 114324 436872
rect 113265 436867 113331 436870
rect 114318 436868 114324 436870
rect 114388 436868 114394 436932
rect 262254 436930 262260 436932
rect 262178 436870 262260 436930
rect 262324 436930 262371 436932
rect 263358 436930 263364 436932
rect 262324 436928 263364 436930
rect 263428 436930 263475 436932
rect 263428 436928 263556 436930
rect 262366 436872 263364 436928
rect 263470 436872 263556 436928
rect 262254 436868 262260 436870
rect 262324 436870 263364 436872
rect 262324 436868 262371 436870
rect 263358 436868 263364 436870
rect 263428 436870 263556 436872
rect 263428 436868 263475 436870
rect 262305 436867 262371 436868
rect 263409 436867 263475 436868
rect 95601 436794 95667 436797
rect 187141 436794 187207 436797
rect 95601 436792 187207 436794
rect -960 436508 480 436748
rect 95601 436736 95606 436792
rect 95662 436736 187146 436792
rect 187202 436736 187207 436792
rect 95601 436734 187207 436736
rect 95601 436731 95667 436734
rect 187141 436731 187207 436734
rect 192477 436658 192543 436661
rect 192477 436656 193660 436658
rect 192477 436600 192482 436656
rect 192538 436600 193660 436656
rect 192477 436598 193660 436600
rect 192477 436595 192543 436598
rect 255405 436386 255471 436389
rect 253460 436384 255471 436386
rect 253460 436328 255410 436384
rect 255466 436328 255471 436384
rect 253460 436326 255471 436328
rect 255405 436323 255471 436326
rect 61929 436250 61995 436253
rect 80973 436250 81039 436253
rect 61929 436248 81039 436250
rect 61929 436192 61934 436248
rect 61990 436192 80978 436248
rect 81034 436192 81039 436248
rect 61929 436190 81039 436192
rect 61929 436187 61995 436190
rect 80973 436187 81039 436190
rect 94630 436188 94636 436252
rect 94700 436250 94706 436252
rect 101213 436250 101279 436253
rect 94700 436248 101279 436250
rect 94700 436192 101218 436248
rect 101274 436192 101279 436248
rect 94700 436190 101279 436192
rect 94700 436188 94706 436190
rect 101213 436187 101279 436190
rect 71865 436116 71931 436117
rect 71814 436114 71820 436116
rect 71738 436054 71820 436114
rect 71884 436114 71931 436116
rect 72693 436114 72759 436117
rect 71884 436112 72759 436114
rect 71926 436056 72698 436112
rect 72754 436056 72759 436112
rect 71814 436052 71820 436054
rect 71884 436054 72759 436056
rect 71884 436052 71931 436054
rect 71865 436051 71931 436052
rect 72693 436051 72759 436054
rect 80329 436114 80395 436117
rect 81014 436114 81020 436116
rect 80329 436112 81020 436114
rect 80329 436056 80334 436112
rect 80390 436056 81020 436112
rect 80329 436054 81020 436056
rect 80329 436051 80395 436054
rect 81014 436052 81020 436054
rect 81084 436114 81090 436116
rect 81341 436114 81407 436117
rect 81084 436112 81407 436114
rect 81084 436056 81346 436112
rect 81402 436056 81407 436112
rect 81084 436054 81407 436056
rect 81084 436052 81090 436054
rect 81341 436051 81407 436054
rect 83089 436114 83155 436117
rect 83590 436114 83596 436116
rect 83089 436112 83596 436114
rect 83089 436056 83094 436112
rect 83150 436056 83596 436112
rect 83089 436054 83596 436056
rect 83089 436051 83155 436054
rect 83590 436052 83596 436054
rect 83660 436052 83666 436116
rect 94446 436052 94452 436116
rect 94516 436114 94522 436116
rect 96889 436114 96955 436117
rect 94516 436112 96955 436114
rect 94516 436056 96894 436112
rect 96950 436056 96955 436112
rect 94516 436054 96955 436056
rect 94516 436052 94522 436054
rect 96889 436051 96955 436054
rect 73654 435372 73660 435436
rect 73724 435434 73730 435436
rect 75821 435434 75887 435437
rect 73724 435432 75887 435434
rect 73724 435376 75826 435432
rect 75882 435376 75887 435432
rect 73724 435374 75887 435376
rect 73724 435372 73730 435374
rect 75821 435371 75887 435374
rect 72601 435298 72667 435301
rect 132493 435298 132559 435301
rect 72601 435296 132559 435298
rect 72601 435240 72606 435296
rect 72662 435240 132498 435296
rect 132554 435240 132559 435296
rect 72601 435238 132559 435240
rect 72601 435235 72667 435238
rect 132493 435235 132559 435238
rect 191557 435298 191623 435301
rect 191557 435296 193660 435298
rect 191557 435240 191562 435296
rect 191618 435240 193660 435296
rect 191557 435238 193660 435240
rect 191557 435235 191623 435238
rect 255405 435026 255471 435029
rect 253460 435024 255471 435026
rect 253460 434968 255410 435024
rect 255466 434968 255471 435024
rect 253460 434966 255471 434968
rect 255405 434963 255471 434966
rect 71221 434890 71287 434893
rect 71630 434890 71636 434892
rect 71221 434888 71636 434890
rect 71221 434832 71226 434888
rect 71282 434832 71636 434888
rect 71221 434830 71636 434832
rect 71221 434827 71287 434830
rect 71630 434828 71636 434830
rect 71700 434890 71706 434892
rect 71700 434830 74550 434890
rect 71700 434828 71706 434830
rect 68001 434754 68067 434757
rect 73797 434754 73863 434757
rect 74165 434754 74231 434757
rect 68001 434752 74231 434754
rect 68001 434696 68006 434752
rect 68062 434696 73802 434752
rect 73858 434696 74170 434752
rect 74226 434696 74231 434752
rect 68001 434694 74231 434696
rect 74490 434754 74550 434830
rect 116577 434754 116643 434757
rect 74490 434752 116643 434754
rect 74490 434696 116582 434752
rect 116638 434696 116643 434752
rect 74490 434694 116643 434696
rect 68001 434691 68067 434694
rect 73797 434691 73863 434694
rect 74165 434691 74231 434694
rect 116577 434691 116643 434694
rect 67398 434556 67404 434620
rect 67468 434618 67474 434620
rect 71221 434618 71287 434621
rect 67468 434616 71287 434618
rect 67468 434560 71226 434616
rect 71282 434560 71287 434616
rect 67468 434558 71287 434560
rect 67468 434556 67474 434558
rect 71221 434555 71287 434558
rect 102726 434556 102732 434620
rect 102796 434618 102802 434620
rect 104893 434618 104959 434621
rect 102796 434616 104959 434618
rect 102796 434560 104898 434616
rect 104954 434560 104959 434616
rect 102796 434558 104959 434560
rect 102796 434556 102802 434558
rect 104893 434555 104959 434558
rect 69054 434284 69060 434348
rect 69124 434346 69130 434348
rect 69197 434346 69263 434349
rect 69124 434344 69263 434346
rect 69124 434288 69202 434344
rect 69258 434288 69263 434344
rect 69124 434286 69263 434288
rect 69124 434284 69130 434286
rect 69197 434283 69263 434286
rect 76373 434348 76439 434349
rect 81893 434348 81959 434349
rect 83089 434348 83155 434349
rect 76373 434344 76420 434348
rect 76484 434346 76490 434348
rect 76373 434288 76378 434344
rect 76373 434284 76420 434288
rect 76484 434286 76530 434346
rect 81893 434344 81940 434348
rect 82004 434346 82010 434348
rect 83038 434346 83044 434348
rect 81893 434288 81898 434344
rect 76484 434284 76490 434286
rect 81893 434284 81940 434288
rect 82004 434286 82050 434346
rect 82998 434286 83044 434346
rect 83108 434344 83155 434348
rect 83150 434288 83155 434344
rect 82004 434284 82010 434286
rect 83038 434284 83044 434286
rect 83108 434284 83155 434288
rect 76373 434283 76439 434284
rect 81893 434283 81959 434284
rect 83089 434283 83155 434284
rect 84653 434348 84719 434349
rect 85849 434348 85915 434349
rect 84653 434344 84700 434348
rect 84764 434346 84770 434348
rect 85798 434346 85804 434348
rect 84653 434288 84658 434344
rect 84653 434284 84700 434288
rect 84764 434286 84810 434346
rect 85758 434286 85804 434346
rect 85868 434344 85915 434348
rect 85910 434288 85915 434344
rect 84764 434284 84770 434286
rect 85798 434284 85804 434286
rect 85868 434284 85915 434288
rect 84653 434283 84719 434284
rect 85849 434283 85915 434284
rect 96245 434348 96311 434349
rect 96245 434344 96292 434348
rect 96356 434346 96362 434348
rect 100385 434346 100451 434349
rect 100518 434346 100524 434348
rect 96245 434288 96250 434344
rect 96245 434284 96292 434288
rect 96356 434286 96402 434346
rect 100385 434344 100524 434346
rect 100385 434288 100390 434344
rect 100446 434288 100524 434344
rect 100385 434286 100524 434288
rect 96356 434284 96362 434286
rect 96245 434283 96311 434284
rect 100385 434283 100451 434286
rect 100518 434284 100524 434286
rect 100588 434284 100594 434348
rect 92841 434210 92907 434213
rect 92974 434210 92980 434212
rect 92841 434208 92980 434210
rect 92841 434152 92846 434208
rect 92902 434152 92980 434208
rect 92841 434150 92980 434152
rect 92841 434147 92907 434150
rect 92974 434148 92980 434150
rect 93044 434148 93050 434212
rect 83222 434012 83228 434076
rect 83292 434074 83298 434076
rect 83825 434074 83891 434077
rect 83292 434072 83891 434074
rect 83292 434016 83830 434072
rect 83886 434016 83891 434072
rect 83292 434014 83891 434016
rect 83292 434012 83298 434014
rect 83825 434011 83891 434014
rect 85849 434074 85915 434077
rect 85849 434072 93870 434074
rect 85849 434016 85854 434072
rect 85910 434016 93870 434072
rect 85849 434014 93870 434016
rect 85849 434011 85915 434014
rect 67950 433876 67956 433940
rect 68020 433938 68026 433940
rect 68020 433878 93226 433938
rect 68020 433876 68026 433878
rect 70894 433740 70900 433804
rect 70964 433802 70970 433804
rect 77109 433802 77175 433805
rect 70964 433800 77175 433802
rect 70964 433744 77114 433800
rect 77170 433744 77175 433800
rect 70964 433742 77175 433744
rect 70964 433740 70970 433742
rect 77109 433739 77175 433742
rect 74574 433604 74580 433668
rect 74644 433666 74650 433668
rect 75453 433666 75519 433669
rect 74644 433664 75519 433666
rect 74644 433608 75458 433664
rect 75514 433608 75519 433664
rect 74644 433606 75519 433608
rect 74644 433604 74650 433606
rect 75453 433603 75519 433606
rect 77334 433604 77340 433668
rect 77404 433666 77410 433668
rect 77477 433666 77543 433669
rect 77404 433664 77543 433666
rect 77404 433608 77482 433664
rect 77538 433608 77543 433664
rect 77404 433606 77543 433608
rect 77404 433604 77410 433606
rect 77477 433603 77543 433606
rect 87086 433604 87092 433668
rect 87156 433666 87162 433668
rect 87229 433666 87295 433669
rect 87156 433664 87295 433666
rect 87156 433608 87234 433664
rect 87290 433608 87295 433664
rect 87156 433606 87295 433608
rect 87156 433604 87162 433606
rect 87229 433603 87295 433606
rect 87454 433604 87460 433668
rect 87524 433666 87530 433668
rect 87965 433666 88031 433669
rect 87524 433664 88031 433666
rect 87524 433608 87970 433664
rect 88026 433608 88031 433664
rect 87524 433606 88031 433608
rect 87524 433604 87530 433606
rect 87965 433603 88031 433606
rect 89621 433668 89687 433669
rect 90081 433668 90147 433669
rect 89621 433664 89668 433668
rect 89732 433666 89738 433668
rect 90030 433666 90036 433668
rect 89621 433608 89626 433664
rect 89621 433604 89668 433608
rect 89732 433606 89778 433666
rect 89990 433606 90036 433666
rect 90100 433664 90147 433668
rect 91277 433668 91343 433669
rect 91553 433668 91619 433669
rect 91277 433666 91324 433668
rect 90142 433608 90147 433664
rect 89732 433604 89738 433606
rect 90030 433604 90036 433606
rect 90100 433604 90147 433608
rect 91232 433664 91324 433666
rect 91232 433608 91282 433664
rect 91232 433606 91324 433608
rect 89621 433603 89687 433604
rect 90081 433603 90147 433604
rect 91277 433604 91324 433606
rect 91388 433604 91394 433668
rect 91502 433666 91508 433668
rect 91462 433606 91508 433666
rect 91572 433664 91619 433668
rect 91614 433608 91619 433664
rect 91502 433604 91508 433606
rect 91572 433604 91619 433608
rect 92790 433604 92796 433668
rect 92860 433666 92866 433668
rect 92933 433666 92999 433669
rect 92860 433664 92999 433666
rect 92860 433608 92938 433664
rect 92994 433608 92999 433664
rect 92860 433606 92999 433608
rect 93166 433666 93226 433878
rect 93810 433802 93870 434014
rect 97717 433938 97783 433941
rect 101121 433938 101187 433941
rect 97717 433936 101187 433938
rect 97717 433880 97722 433936
rect 97778 433880 101126 433936
rect 101182 433880 101187 433936
rect 97717 433878 101187 433880
rect 97717 433875 97783 433878
rect 101121 433875 101187 433878
rect 105353 433938 105419 433941
rect 110137 433938 110203 433941
rect 105353 433936 110203 433938
rect 105353 433880 105358 433936
rect 105414 433880 110142 433936
rect 110198 433880 110203 433936
rect 105353 433878 110203 433880
rect 105353 433875 105419 433878
rect 110137 433875 110203 433878
rect 118877 433802 118943 433805
rect 93810 433800 118943 433802
rect 93810 433744 118882 433800
rect 118938 433744 118943 433800
rect 93810 433742 118943 433744
rect 118877 433739 118943 433742
rect 97717 433666 97783 433669
rect 93166 433664 97783 433666
rect 93166 433608 97722 433664
rect 97778 433608 97783 433664
rect 93166 433606 97783 433608
rect 92860 433604 92866 433606
rect 91277 433603 91343 433604
rect 91553 433603 91619 433604
rect 92933 433603 92999 433606
rect 97717 433603 97783 433606
rect 97942 433604 97948 433668
rect 98012 433666 98018 433668
rect 98361 433666 98427 433669
rect 98012 433664 98427 433666
rect 98012 433608 98366 433664
rect 98422 433608 98427 433664
rect 98012 433606 98427 433608
rect 98012 433604 98018 433606
rect 98361 433603 98427 433606
rect 98494 433604 98500 433668
rect 98564 433666 98570 433668
rect 99189 433666 99255 433669
rect 98564 433664 99255 433666
rect 98564 433608 99194 433664
rect 99250 433608 99255 433664
rect 98564 433606 99255 433608
rect 98564 433604 98570 433606
rect 99189 433603 99255 433606
rect 100661 433668 100727 433669
rect 100661 433664 100708 433668
rect 100772 433666 100778 433668
rect 101121 433666 101187 433669
rect 105353 433666 105419 433669
rect 100661 433608 100666 433664
rect 100661 433604 100708 433608
rect 100772 433606 100818 433666
rect 101121 433664 105419 433666
rect 101121 433608 101126 433664
rect 101182 433608 105358 433664
rect 105414 433608 105419 433664
rect 101121 433606 105419 433608
rect 100772 433604 100778 433606
rect 100661 433603 100727 433604
rect 101121 433603 101187 433606
rect 105353 433603 105419 433606
rect 105486 433604 105492 433668
rect 105556 433666 105562 433668
rect 106733 433666 106799 433669
rect 109033 433668 109099 433669
rect 108982 433666 108988 433668
rect 105556 433664 106799 433666
rect 105556 433608 106738 433664
rect 106794 433608 106799 433664
rect 105556 433606 106799 433608
rect 108942 433606 108988 433666
rect 109052 433664 109099 433668
rect 109094 433608 109099 433664
rect 105556 433604 105562 433606
rect 106733 433603 106799 433606
rect 108982 433604 108988 433606
rect 109052 433604 109099 433608
rect 109033 433603 109099 433604
rect 110137 433666 110203 433669
rect 255405 433666 255471 433669
rect 110137 433664 193660 433666
rect 110137 433608 110142 433664
rect 110198 433608 193660 433664
rect 110137 433606 193660 433608
rect 253460 433664 255471 433666
rect 253460 433608 255410 433664
rect 255466 433608 255471 433664
rect 253460 433606 255471 433608
rect 110137 433603 110203 433606
rect 255405 433603 255471 433606
rect 66805 433394 66871 433397
rect 115749 433394 115815 433397
rect 66805 433392 68908 433394
rect 66805 433336 66810 433392
rect 66866 433336 68908 433392
rect 66805 433334 68908 433336
rect 112700 433392 115815 433394
rect 112700 433336 115754 433392
rect 115810 433336 115815 433392
rect 112700 433334 115815 433336
rect 66805 433331 66871 433334
rect 115749 433331 115815 433334
rect 68645 433122 68711 433125
rect 68645 433120 68938 433122
rect 68645 433064 68650 433120
rect 68706 433064 68938 433120
rect 68645 433062 68938 433064
rect 68645 433059 68711 433062
rect 67541 432578 67607 432581
rect 68878 432578 68938 433062
rect 67541 432576 68938 432578
rect 67541 432520 67546 432576
rect 67602 432548 68938 432576
rect 67602 432520 68908 432548
rect 67541 432518 68908 432520
rect 67541 432515 67607 432518
rect 115841 432306 115907 432309
rect 112700 432304 115907 432306
rect 112700 432248 115846 432304
rect 115902 432248 115907 432304
rect 112700 432246 115907 432248
rect 115841 432243 115907 432246
rect 190637 432306 190703 432309
rect 190637 432304 193660 432306
rect 190637 432248 190642 432304
rect 190698 432248 193660 432304
rect 190637 432246 193660 432248
rect 190637 432243 190703 432246
rect 255405 432034 255471 432037
rect 253460 432032 255471 432034
rect 253460 431976 255410 432032
rect 255466 431976 255471 432032
rect 253460 431974 255471 431976
rect 255405 431971 255471 431974
rect 68369 431898 68435 431901
rect 68369 431896 68938 431898
rect 68369 431840 68374 431896
rect 68430 431840 68938 431896
rect 68369 431838 68938 431840
rect 68369 431835 68435 431838
rect 68878 430810 68938 431838
rect 582465 431626 582531 431629
rect 583520 431626 584960 431716
rect 582465 431624 584960 431626
rect 582465 431568 582470 431624
rect 582526 431568 584960 431624
rect 582465 431566 584960 431568
rect 582465 431563 582531 431566
rect 583520 431476 584960 431566
rect 115841 431218 115907 431221
rect 112700 431216 115907 431218
rect 112700 431160 115846 431216
rect 115902 431160 115907 431216
rect 112700 431158 115907 431160
rect 115841 431155 115907 431158
rect 254669 431218 254735 431221
rect 281574 431218 281580 431220
rect 254669 431216 281580 431218
rect 254669 431160 254674 431216
rect 254730 431160 281580 431216
rect 254669 431158 281580 431160
rect 254669 431155 254735 431158
rect 281574 431156 281580 431158
rect 281644 431156 281650 431220
rect 191097 430946 191163 430949
rect 191097 430944 193660 430946
rect 191097 430888 191102 430944
rect 191158 430888 193660 430944
rect 191097 430886 193660 430888
rect 191097 430883 191163 430886
rect 64830 430750 68938 430810
rect 58893 430674 58959 430677
rect 64830 430674 64890 430750
rect 255405 430674 255471 430677
rect 58893 430672 64890 430674
rect 58893 430616 58898 430672
rect 58954 430616 64890 430672
rect 58893 430614 64890 430616
rect 253460 430672 255471 430674
rect 253460 430616 255410 430672
rect 255466 430616 255471 430672
rect 253460 430614 255471 430616
rect 58893 430611 58959 430614
rect 255405 430611 255471 430614
rect 66069 430402 66135 430405
rect 66069 430400 68908 430402
rect 66069 430344 66074 430400
rect 66130 430344 68908 430400
rect 66069 430342 68908 430344
rect 66069 430339 66135 430342
rect 114553 430130 114619 430133
rect 112700 430128 114619 430130
rect 112700 430072 114558 430128
rect 114614 430072 114619 430128
rect 112700 430070 114619 430072
rect 114553 430067 114619 430070
rect 69422 429796 69428 429860
rect 69492 429796 69498 429860
rect 112713 429858 112779 429861
rect 112670 429856 112779 429858
rect 112670 429800 112718 429856
rect 112774 429800 112779 429856
rect 61653 429314 61719 429317
rect 69430 429314 69490 429796
rect 61653 429312 69490 429314
rect 61653 429256 61658 429312
rect 61714 429284 69490 429312
rect 112670 429795 112779 429800
rect 112670 429284 112730 429795
rect 191189 429586 191255 429589
rect 191189 429584 193660 429586
rect 191189 429528 191194 429584
rect 191250 429528 193660 429584
rect 191189 429526 193660 429528
rect 191189 429523 191255 429526
rect 255497 429314 255563 429317
rect 253460 429312 255563 429314
rect 61714 429256 69460 429284
rect 61653 429254 69460 429256
rect 253460 429256 255502 429312
rect 255558 429256 255563 429312
rect 253460 429254 255563 429256
rect 61653 429251 61719 429254
rect 255497 429251 255563 429254
rect 67081 428226 67147 428229
rect 115841 428226 115907 428229
rect 67081 428224 68908 428226
rect 67081 428168 67086 428224
rect 67142 428168 68908 428224
rect 67081 428166 68908 428168
rect 112700 428224 115907 428226
rect 112700 428168 115846 428224
rect 115902 428168 115907 428224
rect 112700 428166 115907 428168
rect 67081 428163 67147 428166
rect 115841 428163 115907 428166
rect 191741 428226 191807 428229
rect 191741 428224 193660 428226
rect 191741 428168 191746 428224
rect 191802 428168 193660 428224
rect 191741 428166 193660 428168
rect 191741 428163 191807 428166
rect 255405 427954 255471 427957
rect 253460 427952 255471 427954
rect 253460 427896 255410 427952
rect 255466 427896 255471 427952
rect 253460 427894 255471 427896
rect 255405 427891 255471 427894
rect 66989 427410 67055 427413
rect 67265 427410 67331 427413
rect 66989 427408 68908 427410
rect 66989 427352 66994 427408
rect 67050 427352 67270 427408
rect 67326 427352 68908 427408
rect 66989 427350 68908 427352
rect 66989 427347 67055 427350
rect 67265 427347 67331 427350
rect 112118 426596 112178 427108
rect 190637 426866 190703 426869
rect 190637 426864 193660 426866
rect 190637 426808 190642 426864
rect 190698 426808 193660 426864
rect 190637 426806 193660 426808
rect 190637 426803 190703 426806
rect 112110 426532 112116 426596
rect 112180 426532 112186 426596
rect 255497 426594 255563 426597
rect 253460 426592 255563 426594
rect 253460 426536 255502 426592
rect 255558 426536 255563 426592
rect 253460 426534 255563 426536
rect 255497 426531 255563 426534
rect 67265 426322 67331 426325
rect 67541 426322 67607 426325
rect 67265 426320 68908 426322
rect 67265 426264 67270 426320
rect 67326 426264 67546 426320
rect 67602 426264 68908 426320
rect 67265 426262 68908 426264
rect 67265 426259 67331 426262
rect 67541 426259 67607 426262
rect 113357 426050 113423 426053
rect 115381 426050 115447 426053
rect 112700 426048 115447 426050
rect 112700 425992 113362 426048
rect 113418 425992 115386 426048
rect 115442 425992 115447 426048
rect 112700 425990 115447 425992
rect 113357 425987 113423 425990
rect 115381 425987 115447 425990
rect 191741 425506 191807 425509
rect 191741 425504 193660 425506
rect 191741 425448 191746 425504
rect 191802 425448 193660 425504
rect 191741 425446 193660 425448
rect 191741 425443 191807 425446
rect 65977 425234 66043 425237
rect 255865 425234 255931 425237
rect 65977 425232 68908 425234
rect 65977 425176 65982 425232
rect 66038 425176 68908 425232
rect 65977 425174 68908 425176
rect 253460 425232 255931 425234
rect 253460 425176 255870 425232
rect 255926 425176 255931 425232
rect 253460 425174 255931 425176
rect 65977 425171 66043 425174
rect 255865 425171 255931 425174
rect 115381 424962 115447 424965
rect 112700 424960 115447 424962
rect 112700 424904 115386 424960
rect 115442 424904 115447 424960
rect 112700 424902 115447 424904
rect 115381 424899 115447 424902
rect 66621 424146 66687 424149
rect 115013 424146 115079 424149
rect 66621 424144 68908 424146
rect 66621 424088 66626 424144
rect 66682 424088 68908 424144
rect 66621 424086 68908 424088
rect 112700 424144 115079 424146
rect 112700 424088 115018 424144
rect 115074 424088 115079 424144
rect 112700 424086 115079 424088
rect 66621 424083 66687 424086
rect 115013 424083 115079 424086
rect 193814 423740 193874 423844
rect -960 423602 480 423692
rect 193806 423676 193812 423740
rect 193876 423676 193882 423740
rect 3417 423602 3483 423605
rect 255497 423602 255563 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect 253460 423600 255563 423602
rect 253460 423544 255502 423600
rect 255558 423544 255563 423600
rect 253460 423542 255563 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 255497 423539 255563 423542
rect 66805 423330 66871 423333
rect 66805 423328 68908 423330
rect 66805 423272 66810 423328
rect 66866 423272 68908 423328
rect 66805 423270 68908 423272
rect 66805 423267 66871 423270
rect 115013 423058 115079 423061
rect 112700 423056 115079 423058
rect 112700 423000 115018 423056
rect 115074 423000 115079 423056
rect 112700 422998 115079 423000
rect 115013 422995 115079 422998
rect 190637 422514 190703 422517
rect 190637 422512 193660 422514
rect 190637 422456 190642 422512
rect 190698 422456 193660 422512
rect 190637 422454 193660 422456
rect 190637 422451 190703 422454
rect 67081 422242 67147 422245
rect 67950 422242 67956 422244
rect 67081 422240 67956 422242
rect 67081 422184 67086 422240
rect 67142 422184 67956 422240
rect 67081 422182 67956 422184
rect 67081 422179 67147 422182
rect 67950 422180 67956 422182
rect 68020 422242 68026 422244
rect 255497 422242 255563 422245
rect 68020 422182 68908 422242
rect 253460 422240 255563 422242
rect 253460 422184 255502 422240
rect 255558 422184 255563 422240
rect 253460 422182 255563 422184
rect 68020 422180 68026 422182
rect 255497 422179 255563 422182
rect 115197 421970 115263 421973
rect 112700 421968 115263 421970
rect 112700 421912 115202 421968
rect 115258 421912 115263 421968
rect 112700 421910 115263 421912
rect 115197 421907 115263 421910
rect 66621 421154 66687 421157
rect 66621 421152 68908 421154
rect 66621 421096 66626 421152
rect 66682 421096 68908 421152
rect 66621 421094 68908 421096
rect 66621 421091 66687 421094
rect 190361 421018 190427 421021
rect 193630 421018 193690 421124
rect 190361 421016 193690 421018
rect 190361 420960 190366 421016
rect 190422 420960 193690 421016
rect 190361 420958 193690 420960
rect 190361 420955 190427 420958
rect 115749 420882 115815 420885
rect 255497 420882 255563 420885
rect 112700 420880 115815 420882
rect 112700 420824 115754 420880
rect 115810 420824 115815 420880
rect 112700 420822 115815 420824
rect 253460 420880 255563 420882
rect 253460 420824 255502 420880
rect 255558 420824 255563 420880
rect 253460 420822 255563 420824
rect 115749 420819 115815 420822
rect 255497 420819 255563 420822
rect 66805 420066 66871 420069
rect 113541 420066 113607 420069
rect 66805 420064 68908 420066
rect 66805 420008 66810 420064
rect 66866 420008 68908 420064
rect 66805 420006 68908 420008
rect 112700 420064 113607 420066
rect 112700 420008 113546 420064
rect 113602 420008 113607 420064
rect 112700 420006 113607 420008
rect 66805 420003 66871 420006
rect 113541 420003 113607 420006
rect 191741 419794 191807 419797
rect 191741 419792 193660 419794
rect 191741 419736 191746 419792
rect 191802 419736 193660 419792
rect 191741 419734 193660 419736
rect 191741 419731 191807 419734
rect 255405 419522 255471 419525
rect 253460 419520 255471 419522
rect 253460 419464 255410 419520
rect 255466 419464 255471 419520
rect 253460 419462 255471 419464
rect 255405 419459 255471 419462
rect 66805 418978 66871 418981
rect 66805 418976 68908 418978
rect 66805 418920 66810 418976
rect 66866 418920 68908 418976
rect 66805 418918 68908 418920
rect 66805 418915 66871 418918
rect 112670 418437 112730 418948
rect 112670 418432 112779 418437
rect 112670 418376 112718 418432
rect 112774 418376 112779 418432
rect 112670 418374 112779 418376
rect 112713 418371 112779 418374
rect 191741 418434 191807 418437
rect 191741 418432 193660 418434
rect 191741 418376 191746 418432
rect 191802 418376 193660 418432
rect 191741 418374 193660 418376
rect 191741 418371 191807 418374
rect 583017 418298 583083 418301
rect 583520 418298 584960 418388
rect 583017 418296 584960 418298
rect 583017 418240 583022 418296
rect 583078 418240 584960 418296
rect 583017 418238 584960 418240
rect 583017 418235 583083 418238
rect 67081 418162 67147 418165
rect 67449 418162 67515 418165
rect 255497 418162 255563 418165
rect 67081 418160 68908 418162
rect 67081 418104 67086 418160
rect 67142 418104 67454 418160
rect 67510 418104 68908 418160
rect 67081 418102 68908 418104
rect 253460 418160 255563 418162
rect 253460 418104 255502 418160
rect 255558 418104 255563 418160
rect 583520 418148 584960 418238
rect 253460 418102 255563 418104
rect 67081 418099 67147 418102
rect 67449 418099 67515 418102
rect 255497 418099 255563 418102
rect 114645 417890 114711 417893
rect 112700 417888 114711 417890
rect 112700 417832 114650 417888
rect 114706 417832 114711 417888
rect 112700 417830 114711 417832
rect 114645 417827 114711 417830
rect 41321 417482 41387 417485
rect 66294 417482 66300 417484
rect 41321 417480 66300 417482
rect 41321 417424 41326 417480
rect 41382 417424 66300 417480
rect 41321 417422 66300 417424
rect 41321 417419 41387 417422
rect 66294 417420 66300 417422
rect 66364 417420 66370 417484
rect 67633 417074 67699 417077
rect 191741 417074 191807 417077
rect 67633 417072 68908 417074
rect 67633 417016 67638 417072
rect 67694 417016 68908 417072
rect 67633 417014 68908 417016
rect 191741 417072 193660 417074
rect 191741 417016 191746 417072
rect 191802 417016 193660 417072
rect 191741 417014 193660 417016
rect 67633 417011 67699 417014
rect 191741 417011 191807 417014
rect 113265 416802 113331 416805
rect 113909 416802 113975 416805
rect 255405 416802 255471 416805
rect 112700 416800 113975 416802
rect 112700 416744 113270 416800
rect 113326 416744 113914 416800
rect 113970 416744 113975 416800
rect 112700 416742 113975 416744
rect 253460 416800 255471 416802
rect 253460 416744 255410 416800
rect 255466 416744 255471 416800
rect 253460 416742 255471 416744
rect 113265 416739 113331 416742
rect 113909 416739 113975 416742
rect 255405 416739 255471 416742
rect 66253 415986 66319 415989
rect 66253 415984 68908 415986
rect 66253 415928 66258 415984
rect 66314 415928 68908 415984
rect 66253 415926 68908 415928
rect 66253 415923 66319 415926
rect 177246 415924 177252 415988
rect 177316 415986 177322 415988
rect 187693 415986 187759 415989
rect 177316 415984 187759 415986
rect 177316 415928 187698 415984
rect 187754 415928 187759 415984
rect 177316 415926 187759 415928
rect 177316 415924 177322 415926
rect 187693 415923 187759 415926
rect 115841 415714 115907 415717
rect 112700 415712 115907 415714
rect 112700 415656 115846 415712
rect 115902 415656 115907 415712
rect 112700 415654 115907 415656
rect 115841 415651 115907 415654
rect 190637 415442 190703 415445
rect 190637 415440 193660 415442
rect 190637 415384 190642 415440
rect 190698 415384 193660 415440
rect 190637 415382 193660 415384
rect 190637 415379 190703 415382
rect 254025 415170 254091 415173
rect 253460 415168 254091 415170
rect 253460 415112 254030 415168
rect 254086 415112 254091 415168
rect 253460 415110 254091 415112
rect 254025 415107 254091 415110
rect 66805 414898 66871 414901
rect 115841 414898 115907 414901
rect 66805 414896 68908 414898
rect 66805 414840 66810 414896
rect 66866 414840 68908 414896
rect 66805 414838 68908 414840
rect 112700 414896 115907 414898
rect 112700 414840 115846 414896
rect 115902 414840 115907 414896
rect 112700 414838 115907 414840
rect 66805 414835 66871 414838
rect 115841 414835 115907 414838
rect 61745 414354 61811 414357
rect 66253 414354 66319 414357
rect 61745 414352 66319 414354
rect 61745 414296 61750 414352
rect 61806 414296 66258 414352
rect 66314 414296 66319 414352
rect 61745 414294 66319 414296
rect 61745 414291 61811 414294
rect 66253 414291 66319 414294
rect 66897 414082 66963 414085
rect 191741 414082 191807 414085
rect 66897 414080 68908 414082
rect 66897 414024 66902 414080
rect 66958 414024 68908 414080
rect 66897 414022 68908 414024
rect 191741 414080 193660 414082
rect 191741 414024 191746 414080
rect 191802 414024 193660 414080
rect 191741 414022 193660 414024
rect 66897 414019 66963 414022
rect 191741 414019 191807 414022
rect 113173 413810 113239 413813
rect 255405 413810 255471 413813
rect 112700 413808 113239 413810
rect 112700 413752 113178 413808
rect 113234 413752 113239 413808
rect 112700 413750 113239 413752
rect 253460 413808 255471 413810
rect 253460 413752 255410 413808
rect 255466 413752 255471 413808
rect 253460 413750 255471 413752
rect 113173 413747 113239 413750
rect 255405 413747 255471 413750
rect 66253 412996 66319 412997
rect 66253 412994 66300 412996
rect 66172 412992 66300 412994
rect 66364 412994 66370 412996
rect 66172 412936 66258 412992
rect 66172 412934 66300 412936
rect 66253 412932 66300 412934
rect 66364 412934 68908 412994
rect 66364 412932 66370 412934
rect 66253 412931 66319 412932
rect 115289 412722 115355 412725
rect 112700 412720 115355 412722
rect 112700 412664 115294 412720
rect 115350 412664 115355 412720
rect 112700 412662 115355 412664
rect 115289 412659 115355 412662
rect 191598 412660 191604 412724
rect 191668 412722 191674 412724
rect 191668 412662 193660 412722
rect 191668 412660 191674 412662
rect 254117 412450 254183 412453
rect 253460 412448 254183 412450
rect 253460 412392 254122 412448
rect 254178 412392 254183 412448
rect 253460 412390 254183 412392
rect 254117 412387 254183 412390
rect 66110 411844 66116 411908
rect 66180 411906 66186 411908
rect 66253 411906 66319 411909
rect 66180 411904 68908 411906
rect 66180 411848 66258 411904
rect 66314 411848 68908 411904
rect 66180 411846 68908 411848
rect 66180 411844 66186 411846
rect 66253 411843 66319 411846
rect 115841 411634 115907 411637
rect 112700 411632 115907 411634
rect 112700 411576 115846 411632
rect 115902 411576 115907 411632
rect 112700 411574 115907 411576
rect 115841 411571 115907 411574
rect 191741 411362 191807 411365
rect 191741 411360 193660 411362
rect 191741 411304 191746 411360
rect 191802 411304 193660 411360
rect 191741 411302 193660 411304
rect 191741 411299 191807 411302
rect 255405 411090 255471 411093
rect 253460 411088 255471 411090
rect 253460 411032 255410 411088
rect 255466 411032 255471 411088
rect 253460 411030 255471 411032
rect 255405 411027 255471 411030
rect 66621 410818 66687 410821
rect 66621 410816 68908 410818
rect 66621 410760 66626 410816
rect 66682 410760 68908 410816
rect 66621 410758 68908 410760
rect 66621 410755 66687 410758
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect 114737 410546 114803 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect 112700 410544 114803 410546
rect 112700 410488 114742 410544
rect 114798 410488 114803 410544
rect 112700 410486 114803 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 114737 410483 114803 410486
rect 151077 410138 151143 410141
rect 122790 410136 151143 410138
rect 122790 410080 151082 410136
rect 151138 410080 151143 410136
rect 122790 410078 151143 410080
rect 115054 409940 115060 410004
rect 115124 409940 115130 410004
rect 122790 410002 122850 410078
rect 151077 410075 151143 410078
rect 115798 409942 122850 410002
rect 191005 410002 191071 410005
rect 191005 410000 193660 410002
rect 191005 409944 191010 410000
rect 191066 409944 193660 410000
rect 191005 409942 193660 409944
rect 115062 409866 115122 409940
rect 115798 409866 115858 409942
rect 191005 409939 191071 409942
rect 113130 409806 115858 409866
rect 67398 409668 67404 409732
rect 67468 409730 67474 409732
rect 113130 409730 113190 409806
rect 255405 409730 255471 409733
rect 67468 409670 68908 409730
rect 112700 409670 113190 409730
rect 253460 409728 255471 409730
rect 253460 409672 255410 409728
rect 255466 409672 255471 409728
rect 253460 409670 255471 409672
rect 67468 409668 67474 409670
rect 255405 409667 255471 409670
rect 66805 408914 66871 408917
rect 66805 408912 68908 408914
rect 66805 408856 66810 408912
rect 66866 408856 68908 408912
rect 66805 408854 68908 408856
rect 66805 408851 66871 408854
rect 115841 408642 115907 408645
rect 112700 408640 115907 408642
rect 112700 408584 115846 408640
rect 115902 408584 115907 408640
rect 112700 408582 115907 408584
rect 115841 408579 115907 408582
rect 191005 408642 191071 408645
rect 191005 408640 193660 408642
rect 191005 408584 191010 408640
rect 191066 408584 193660 408640
rect 191005 408582 193660 408584
rect 191005 408579 191071 408582
rect 255313 408370 255379 408373
rect 253460 408368 255379 408370
rect 253460 408312 255318 408368
rect 255374 408312 255379 408368
rect 253460 408310 255379 408312
rect 255313 408307 255379 408310
rect 66897 407826 66963 407829
rect 66897 407824 68908 407826
rect 66897 407768 66902 407824
rect 66958 407768 68908 407824
rect 66897 407766 68908 407768
rect 66897 407763 66963 407766
rect 115381 407554 115447 407557
rect 112700 407552 115447 407554
rect 112700 407496 115386 407552
rect 115442 407496 115447 407552
rect 112700 407494 115447 407496
rect 115381 407491 115447 407494
rect 191741 407010 191807 407013
rect 255405 407010 255471 407013
rect 191741 407008 193660 407010
rect 191741 406952 191746 407008
rect 191802 406952 193660 407008
rect 191741 406950 193660 406952
rect 253460 407008 255471 407010
rect 253460 406952 255410 407008
rect 255466 406952 255471 407008
rect 253460 406950 255471 406952
rect 191741 406947 191807 406950
rect 255405 406947 255471 406950
rect 66805 406738 66871 406741
rect 66805 406736 68908 406738
rect 66805 406680 66810 406736
rect 66866 406680 68908 406736
rect 66805 406678 68908 406680
rect 66805 406675 66871 406678
rect 115197 406466 115263 406469
rect 112700 406464 115263 406466
rect 112700 406408 115202 406464
rect 115258 406408 115263 406464
rect 112700 406406 115263 406408
rect 115197 406403 115263 406406
rect 67357 405650 67423 405653
rect 115749 405650 115815 405653
rect 67357 405648 68908 405650
rect 67357 405592 67362 405648
rect 67418 405592 68908 405648
rect 67357 405590 68908 405592
rect 112700 405648 115815 405650
rect 112700 405592 115754 405648
rect 115810 405592 115815 405648
rect 112700 405590 115815 405592
rect 67357 405587 67423 405590
rect 115749 405587 115815 405590
rect 191741 405650 191807 405653
rect 191741 405648 193660 405650
rect 191741 405592 191746 405648
rect 191802 405592 193660 405648
rect 191741 405590 193660 405592
rect 191741 405587 191807 405590
rect 114318 405452 114324 405516
rect 114388 405514 114394 405516
rect 114921 405514 114987 405517
rect 114388 405512 114987 405514
rect 114388 405456 114926 405512
rect 114982 405456 114987 405512
rect 114388 405454 114987 405456
rect 114388 405452 114394 405454
rect 114921 405451 114987 405454
rect 254209 405378 254275 405381
rect 253460 405376 254275 405378
rect 253460 405320 254214 405376
rect 254270 405320 254275 405376
rect 253460 405318 254275 405320
rect 254209 405315 254275 405318
rect 583293 404970 583359 404973
rect 583520 404970 584960 405060
rect 583293 404968 584960 404970
rect 583293 404912 583298 404968
rect 583354 404912 584960 404968
rect 583293 404910 584960 404912
rect 583293 404907 583359 404910
rect 583520 404820 584960 404910
rect 66805 404562 66871 404565
rect 115841 404562 115907 404565
rect 66805 404560 68908 404562
rect 66805 404504 66810 404560
rect 66866 404504 68908 404560
rect 66805 404502 68908 404504
rect 112700 404560 115907 404562
rect 112700 404504 115846 404560
rect 115902 404504 115907 404560
rect 112700 404502 115907 404504
rect 66805 404499 66871 404502
rect 115841 404499 115907 404502
rect 114921 404426 114987 404429
rect 169201 404426 169267 404429
rect 114921 404424 169267 404426
rect 114921 404368 114926 404424
rect 114982 404368 169206 404424
rect 169262 404368 169267 404424
rect 114921 404366 169267 404368
rect 114921 404363 114987 404366
rect 169201 404363 169267 404366
rect 191741 404290 191807 404293
rect 191741 404288 193660 404290
rect 191741 404232 191746 404288
rect 191802 404232 193660 404288
rect 191741 404230 193660 404232
rect 191741 404227 191807 404230
rect 256785 404018 256851 404021
rect 253460 404016 256851 404018
rect 253460 403960 256790 404016
rect 256846 403960 256851 404016
rect 253460 403958 256851 403960
rect 256785 403955 256851 403958
rect 66805 403746 66871 403749
rect 66805 403744 68908 403746
rect 66805 403688 66810 403744
rect 66866 403688 68908 403744
rect 66805 403686 68908 403688
rect 66805 403683 66871 403686
rect 115841 403474 115907 403477
rect 112700 403472 115907 403474
rect 112700 403416 115846 403472
rect 115902 403416 115907 403472
rect 112700 403414 115907 403416
rect 115841 403411 115907 403414
rect 67173 402658 67239 402661
rect 67173 402656 68908 402658
rect 67173 402600 67178 402656
rect 67234 402600 68908 402656
rect 67173 402598 68908 402600
rect 67173 402595 67239 402598
rect 113449 402386 113515 402389
rect 112700 402384 113515 402386
rect 112700 402328 113454 402384
rect 113510 402328 113515 402384
rect 112700 402326 113515 402328
rect 113449 402323 113515 402326
rect 191649 402386 191715 402389
rect 193630 402386 193690 402900
rect 191649 402384 193690 402386
rect 191649 402328 191654 402384
rect 191710 402328 193690 402384
rect 191649 402326 193690 402328
rect 191649 402323 191715 402326
rect 253430 402114 253490 402628
rect 253565 402114 253631 402117
rect 253430 402112 253631 402114
rect 253430 402056 253570 402112
rect 253626 402056 253631 402112
rect 253430 402054 253631 402056
rect 253565 402051 253631 402054
rect 66662 401644 66668 401708
rect 66732 401706 66738 401708
rect 67173 401706 67239 401709
rect 66732 401704 67239 401706
rect 66732 401648 67178 401704
rect 67234 401648 67239 401704
rect 66732 401646 67239 401648
rect 66732 401644 66738 401646
rect 67173 401643 67239 401646
rect 66713 401570 66779 401573
rect 66713 401568 68908 401570
rect 66713 401512 66718 401568
rect 66774 401512 68908 401568
rect 66713 401510 68908 401512
rect 66713 401507 66779 401510
rect 115565 401298 115631 401301
rect 112700 401296 115631 401298
rect 112700 401240 115570 401296
rect 115626 401240 115631 401296
rect 112700 401238 115631 401240
rect 115565 401235 115631 401238
rect 67541 400482 67607 400485
rect 114737 400482 114803 400485
rect 67541 400480 68908 400482
rect 67541 400424 67546 400480
rect 67602 400424 68908 400480
rect 67541 400422 68908 400424
rect 112700 400480 114803 400482
rect 112700 400424 114742 400480
rect 114798 400424 114803 400480
rect 112700 400422 114803 400424
rect 67541 400419 67607 400422
rect 114737 400419 114803 400422
rect 188838 400420 188844 400484
rect 188908 400482 188914 400484
rect 193630 400482 193690 401540
rect 255405 401298 255471 401301
rect 253460 401296 255471 401298
rect 253460 401240 255410 401296
rect 255466 401240 255471 401296
rect 253460 401238 255471 401240
rect 255405 401235 255471 401238
rect 188908 400422 193690 400482
rect 188908 400420 188914 400422
rect 191741 400210 191807 400213
rect 191741 400208 193660 400210
rect 191741 400152 191746 400208
rect 191802 400152 193660 400208
rect 191741 400150 193660 400152
rect 191741 400147 191807 400150
rect 255405 399938 255471 399941
rect 253460 399936 255471 399938
rect 253460 399880 255410 399936
rect 255466 399880 255471 399936
rect 253460 399878 255471 399880
rect 255405 399875 255471 399878
rect 66805 399666 66871 399669
rect 66805 399664 68908 399666
rect 66805 399608 66810 399664
rect 66866 399608 68908 399664
rect 66805 399606 68908 399608
rect 66805 399603 66871 399606
rect 57881 399530 57947 399533
rect 65885 399530 65951 399533
rect 57881 399528 65951 399530
rect 57881 399472 57886 399528
rect 57942 399472 65890 399528
rect 65946 399472 65951 399528
rect 57881 399470 65951 399472
rect 57881 399467 57947 399470
rect 65885 399467 65951 399470
rect 115841 399394 115907 399397
rect 112700 399392 115907 399394
rect 112700 399336 115846 399392
rect 115902 399336 115907 399392
rect 112700 399334 115907 399336
rect 115841 399331 115907 399334
rect 65885 398850 65951 398853
rect 65885 398848 68938 398850
rect 65885 398792 65890 398848
rect 65946 398792 68938 398848
rect 65885 398790 68938 398792
rect 65885 398787 65951 398790
rect 68878 398548 68938 398790
rect 190821 398578 190887 398581
rect 190821 398576 193660 398578
rect 190821 398520 190826 398576
rect 190882 398520 193660 398576
rect 190821 398518 193660 398520
rect 190821 398515 190887 398518
rect 115381 398306 115447 398309
rect 112700 398304 115447 398306
rect 112700 398248 115386 398304
rect 115442 398248 115447 398304
rect 112700 398246 115447 398248
rect 115381 398243 115447 398246
rect 253430 398034 253490 398548
rect 255998 398034 256004 398036
rect 253430 397974 256004 398034
rect 255998 397972 256004 397974
rect 256068 398034 256074 398036
rect 582557 398034 582623 398037
rect 256068 398032 582623 398034
rect 256068 397976 582562 398032
rect 582618 397976 582623 398032
rect 256068 397974 582623 397976
rect 256068 397972 256074 397974
rect 582557 397971 582623 397974
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 67173 397490 67239 397493
rect 67766 397490 67772 397492
rect 67173 397488 67772 397490
rect 67173 397432 67178 397488
rect 67234 397432 67772 397488
rect 67173 397430 67772 397432
rect 67173 397427 67239 397430
rect 67766 397428 67772 397430
rect 67836 397490 67842 397492
rect 67836 397430 68908 397490
rect 67836 397428 67842 397430
rect 115197 397354 115263 397357
rect 115749 397354 115815 397357
rect 115197 397352 115815 397354
rect 115197 397296 115202 397352
rect 115258 397296 115754 397352
rect 115810 397296 115815 397352
rect 115197 397294 115815 397296
rect 115197 397291 115263 397294
rect 115749 397291 115815 397294
rect 113214 397218 113220 397220
rect 112700 397158 113220 397218
rect 113214 397156 113220 397158
rect 113284 397218 113290 397220
rect 115289 397218 115355 397221
rect 113284 397216 115355 397218
rect 113284 397160 115294 397216
rect 115350 397160 115355 397216
rect 113284 397158 115355 397160
rect 113284 397156 113290 397158
rect 115289 397155 115355 397158
rect 191741 397218 191807 397221
rect 191741 397216 193660 397218
rect 191741 397160 191746 397216
rect 191802 397160 193660 397216
rect 191741 397158 193660 397160
rect 191741 397155 191807 397158
rect 255313 396946 255379 396949
rect 253460 396944 255379 396946
rect 253460 396888 255318 396944
rect 255374 396888 255379 396944
rect 253460 396886 255379 396888
rect 255313 396883 255379 396886
rect 258717 396674 258783 396677
rect 270534 396674 270540 396676
rect 258717 396672 270540 396674
rect 258717 396616 258722 396672
rect 258778 396616 270540 396672
rect 258717 396614 270540 396616
rect 258717 396611 258783 396614
rect 270534 396612 270540 396614
rect 270604 396612 270610 396676
rect 193990 396538 193996 396540
rect 180750 396478 193996 396538
rect 67817 396402 67883 396405
rect 114921 396402 114987 396405
rect 67817 396400 68908 396402
rect 67817 396344 67822 396400
rect 67878 396344 68908 396400
rect 67817 396342 68908 396344
rect 112700 396400 114987 396402
rect 112700 396344 114926 396400
rect 114982 396344 114987 396400
rect 112700 396342 114987 396344
rect 67817 396339 67883 396342
rect 114921 396339 114987 396342
rect 115749 396266 115815 396269
rect 180750 396266 180810 396478
rect 193990 396476 193996 396478
rect 194060 396476 194066 396540
rect 115749 396264 180810 396266
rect 115749 396208 115754 396264
rect 115810 396208 180810 396264
rect 115749 396206 180810 396208
rect 115749 396203 115815 396206
rect 190821 395858 190887 395861
rect 190821 395856 193660 395858
rect 190821 395800 190826 395856
rect 190882 395800 193660 395856
rect 190821 395798 193660 395800
rect 190821 395795 190887 395798
rect 255497 395586 255563 395589
rect 253460 395584 255563 395586
rect 253460 395528 255502 395584
rect 255558 395528 255563 395584
rect 253460 395526 255563 395528
rect 255497 395523 255563 395526
rect 67173 395314 67239 395317
rect 67909 395314 67975 395317
rect 115841 395314 115907 395317
rect 67173 395312 68908 395314
rect 67173 395256 67178 395312
rect 67234 395256 67914 395312
rect 67970 395256 68908 395312
rect 67173 395254 68908 395256
rect 112700 395312 115907 395314
rect 112700 395256 115846 395312
rect 115902 395256 115907 395312
rect 112700 395254 115907 395256
rect 67173 395251 67239 395254
rect 67909 395251 67975 395254
rect 115841 395251 115907 395254
rect 190821 394498 190887 394501
rect 190821 394496 193660 394498
rect 69430 393956 69490 394468
rect 190821 394440 190826 394496
rect 190882 394440 193660 394496
rect 190821 394438 193660 394440
rect 190821 394435 190887 394438
rect 115749 394226 115815 394229
rect 256877 394226 256943 394229
rect 112700 394224 115815 394226
rect 112700 394168 115754 394224
rect 115810 394168 115815 394224
rect 112700 394166 115815 394168
rect 253460 394224 256943 394226
rect 253460 394168 256882 394224
rect 256938 394168 256943 394224
rect 253460 394166 256943 394168
rect 115749 394163 115815 394166
rect 256877 394163 256943 394166
rect 69422 393892 69428 393956
rect 69492 393892 69498 393956
rect 112846 393484 112852 393548
rect 112916 393546 112922 393548
rect 112916 393486 161490 393546
rect 112916 393484 112922 393486
rect 67633 393410 67699 393413
rect 161430 393410 161490 393486
rect 165521 393410 165587 393413
rect 190453 393410 190519 393413
rect 67633 393408 68908 393410
rect 67633 393352 67638 393408
rect 67694 393352 68908 393408
rect 67633 393350 68908 393352
rect 161430 393408 190519 393410
rect 161430 393352 165526 393408
rect 165582 393352 190458 393408
rect 190514 393352 190519 393408
rect 161430 393350 190519 393352
rect 67633 393347 67699 393350
rect 165521 393347 165587 393350
rect 190453 393347 190519 393350
rect 115565 393138 115631 393141
rect 112700 393136 115631 393138
rect 112700 393080 115570 393136
rect 115626 393080 115631 393136
rect 112700 393078 115631 393080
rect 115565 393075 115631 393078
rect 191557 393138 191623 393141
rect 191557 393136 193660 393138
rect 191557 393080 191562 393136
rect 191618 393080 193660 393136
rect 191557 393078 193660 393080
rect 191557 393075 191623 393078
rect 255589 392866 255655 392869
rect 253460 392864 255655 392866
rect 253460 392808 255594 392864
rect 255650 392808 255655 392864
rect 253460 392806 255655 392808
rect 255589 392803 255655 392806
rect 66805 392322 66871 392325
rect 66805 392320 68908 392322
rect 66805 392264 66810 392320
rect 66866 392264 68908 392320
rect 66805 392262 68908 392264
rect 66805 392259 66871 392262
rect 115749 392050 115815 392053
rect 112700 392048 115815 392050
rect 112700 391992 115754 392048
rect 115810 391992 115815 392048
rect 112700 391990 115815 391992
rect 115749 391987 115815 391990
rect 190453 391778 190519 391781
rect 190453 391776 193660 391778
rect 190453 391720 190458 391776
rect 190514 391720 193660 391776
rect 190453 391718 193660 391720
rect 190453 391715 190519 391718
rect 583520 391628 584960 391868
rect 114829 391234 114895 391237
rect 112700 391232 114895 391234
rect 69430 390690 69490 391204
rect 112700 391176 114834 391232
rect 114890 391176 114895 391232
rect 112700 391174 114895 391176
rect 114829 391171 114895 391174
rect 117221 391098 117287 391101
rect 73294 391096 117287 391098
rect 73294 391040 117226 391096
rect 117282 391040 117287 391096
rect 73294 391038 117287 391040
rect 70393 390962 70459 390965
rect 71681 390962 71747 390965
rect 73294 390962 73354 391038
rect 117221 391035 117287 391038
rect 70393 390960 73354 390962
rect 70393 390904 70398 390960
rect 70454 390904 71686 390960
rect 71742 390904 73354 390960
rect 70393 390902 73354 390904
rect 70393 390899 70459 390902
rect 71681 390899 71747 390902
rect 73470 390900 73476 390964
rect 73540 390962 73546 390964
rect 73981 390962 74047 390965
rect 73540 390960 74047 390962
rect 73540 390904 73986 390960
rect 74042 390904 74047 390960
rect 73540 390902 74047 390904
rect 73540 390900 73546 390902
rect 73981 390899 74047 390902
rect 111977 390962 112043 390965
rect 193489 390962 193555 390965
rect 111977 390960 193555 390962
rect 111977 390904 111982 390960
rect 112038 390904 193494 390960
rect 193550 390904 193555 390960
rect 111977 390902 193555 390904
rect 111977 390899 112043 390902
rect 193489 390899 193555 390902
rect 252553 390962 252619 390965
rect 252878 390962 252938 391476
rect 252553 390960 252938 390962
rect 252553 390904 252558 390960
rect 252614 390904 252938 390960
rect 252553 390902 252938 390904
rect 252553 390899 252619 390902
rect 91277 390826 91343 390829
rect 223481 390826 223547 390829
rect 91277 390824 223547 390826
rect 91277 390768 91282 390824
rect 91338 390768 223486 390824
rect 223542 390768 223547 390824
rect 91277 390766 223547 390768
rect 91277 390763 91343 390766
rect 223481 390763 223547 390766
rect 107929 390692 107995 390693
rect 107878 390690 107884 390692
rect 69430 390630 107762 390690
rect 107838 390630 107884 390690
rect 107948 390688 107995 390692
rect 112846 390690 112852 390692
rect 107990 390632 107995 390688
rect 96654 390492 96660 390556
rect 96724 390554 96730 390556
rect 96981 390554 97047 390557
rect 96724 390552 97047 390554
rect 96724 390496 96986 390552
rect 97042 390496 97047 390552
rect 96724 390494 97047 390496
rect 96724 390492 96730 390494
rect 96981 390491 97047 390494
rect 101029 390554 101095 390557
rect 101254 390554 101260 390556
rect 101029 390552 101260 390554
rect 101029 390496 101034 390552
rect 101090 390496 101260 390552
rect 101029 390494 101260 390496
rect 101029 390491 101095 390494
rect 101254 390492 101260 390494
rect 101324 390492 101330 390556
rect 107702 390554 107762 390630
rect 107878 390628 107884 390630
rect 107948 390628 107995 390632
rect 107929 390627 107995 390628
rect 108070 390630 112852 390690
rect 108070 390554 108130 390630
rect 112846 390628 112852 390630
rect 112916 390628 112922 390692
rect 107702 390494 108130 390554
rect 193990 390492 193996 390556
rect 194060 390554 194066 390556
rect 254117 390554 254183 390557
rect 194060 390552 254183 390554
rect 194060 390496 254122 390552
rect 254178 390496 254183 390552
rect 194060 390494 254183 390496
rect 194060 390492 194066 390494
rect 254117 390491 254183 390494
rect 99649 390418 99715 390421
rect 99966 390418 99972 390420
rect 99649 390416 99972 390418
rect 99649 390360 99654 390416
rect 99710 390360 99972 390416
rect 99649 390358 99972 390360
rect 99649 390355 99715 390358
rect 99966 390356 99972 390358
rect 100036 390356 100042 390420
rect 104934 390356 104940 390420
rect 105004 390418 105010 390420
rect 105261 390418 105327 390421
rect 105004 390416 105327 390418
rect 105004 390360 105266 390416
rect 105322 390360 105327 390416
rect 105004 390358 105327 390360
rect 105004 390356 105010 390358
rect 105261 390355 105327 390358
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106733 390418 106799 390421
rect 107745 390420 107811 390421
rect 107694 390418 107700 390420
rect 106476 390416 106799 390418
rect 106476 390360 106738 390416
rect 106794 390360 106799 390416
rect 106476 390358 106799 390360
rect 107654 390358 107700 390418
rect 107764 390416 107811 390420
rect 107806 390360 107811 390416
rect 106476 390356 106482 390358
rect 106733 390355 106799 390358
rect 107694 390356 107700 390358
rect 107764 390356 107811 390360
rect 107745 390355 107811 390356
rect 69105 390146 69171 390149
rect 70071 390146 70137 390149
rect 69105 390144 70137 390146
rect 69105 390088 69110 390144
rect 69166 390088 70076 390144
rect 70132 390088 70137 390144
rect 69105 390086 70137 390088
rect 69105 390083 69171 390086
rect 70071 390083 70137 390086
rect 238017 389874 238083 389877
rect 248454 389874 248460 389876
rect 238017 389872 248460 389874
rect 238017 389816 238022 389872
rect 238078 389816 248460 389872
rect 238017 389814 248460 389816
rect 238017 389811 238083 389814
rect 248454 389812 248460 389814
rect 248524 389812 248530 389876
rect 78581 389466 78647 389469
rect 110597 389466 110663 389469
rect 78581 389464 113190 389466
rect 78581 389408 78586 389464
rect 78642 389408 110602 389464
rect 110658 389408 113190 389464
rect 78581 389406 113190 389408
rect 78581 389403 78647 389406
rect 110597 389403 110663 389406
rect 7649 389330 7715 389333
rect 107837 389330 107903 389333
rect 7649 389328 107903 389330
rect 7649 389272 7654 389328
rect 7710 389272 107842 389328
rect 107898 389272 107903 389328
rect 7649 389270 107903 389272
rect 113130 389330 113190 389406
rect 205541 389330 205607 389333
rect 113130 389328 205607 389330
rect 113130 389272 205546 389328
rect 205602 389272 205607 389328
rect 113130 389270 205607 389272
rect 7649 389267 7715 389270
rect 107837 389267 107903 389270
rect 205541 389267 205607 389270
rect 69105 389194 69171 389197
rect 195421 389194 195487 389197
rect 69105 389192 195487 389194
rect 69105 389136 69110 389192
rect 69166 389136 195426 389192
rect 195482 389136 195487 389192
rect 69105 389134 195487 389136
rect 69105 389131 69171 389134
rect 195421 389131 195487 389134
rect 72417 389058 72483 389061
rect 72734 389058 72740 389060
rect 72417 389056 72740 389058
rect 72417 389000 72422 389056
rect 72478 389000 72740 389056
rect 72417 388998 72740 389000
rect 72417 388995 72483 388998
rect 72734 388996 72740 388998
rect 72804 389058 72810 389060
rect 73061 389058 73127 389061
rect 72804 389056 73127 389058
rect 72804 389000 73066 389056
rect 73122 389000 73127 389056
rect 72804 388998 73127 389000
rect 72804 388996 72810 388998
rect 73061 388995 73127 388998
rect 79133 389058 79199 389061
rect 79726 389058 79732 389060
rect 79133 389056 79732 389058
rect 79133 389000 79138 389056
rect 79194 389000 79732 389056
rect 79133 388998 79732 389000
rect 79133 388995 79199 388998
rect 79726 388996 79732 388998
rect 79796 389058 79802 389060
rect 79869 389058 79935 389061
rect 79796 389056 79935 389058
rect 79796 389000 79874 389056
rect 79930 389000 79935 389056
rect 79796 388998 79935 389000
rect 79796 388996 79802 388998
rect 79869 388995 79935 388998
rect 80053 389060 80119 389061
rect 80053 389056 80100 389060
rect 80164 389058 80170 389060
rect 80973 389058 81039 389061
rect 80164 389056 81039 389058
rect 80053 389000 80058 389056
rect 80164 389000 80978 389056
rect 81034 389000 81039 389056
rect 80053 388996 80100 389000
rect 80164 388998 81039 389000
rect 80164 388996 80170 388998
rect 80053 388995 80119 388996
rect 80973 388995 81039 388998
rect 97441 389058 97507 389061
rect 97901 389058 97967 389061
rect 97441 389056 97967 389058
rect 97441 389000 97446 389056
rect 97502 389000 97906 389056
rect 97962 389000 97967 389056
rect 97441 388998 97967 389000
rect 97441 388995 97507 388998
rect 97901 388995 97967 388998
rect 178033 389058 178099 389061
rect 178769 389058 178835 389061
rect 194501 389058 194567 389061
rect 178033 389056 194567 389058
rect 178033 389000 178038 389056
rect 178094 389000 178774 389056
rect 178830 389000 194506 389056
rect 194562 389000 194567 389056
rect 178033 388998 194567 389000
rect 178033 388995 178099 388998
rect 178769 388995 178835 388998
rect 194501 388995 194567 388998
rect 242249 389058 242315 389061
rect 282821 389058 282887 389061
rect 287329 389058 287395 389061
rect 242249 389056 287395 389058
rect 242249 389000 242254 389056
rect 242310 389000 282826 389056
rect 282882 389000 287334 389056
rect 287390 389000 287395 389056
rect 242249 388998 287395 389000
rect 242249 388995 242315 388998
rect 282821 388995 282887 388998
rect 287329 388995 287395 388998
rect 96889 388922 96955 388925
rect 97206 388922 97212 388924
rect 96889 388920 97212 388922
rect 96889 388864 96894 388920
rect 96950 388864 97212 388920
rect 96889 388862 97212 388864
rect 96889 388859 96955 388862
rect 97206 388860 97212 388862
rect 97276 388922 97282 388924
rect 105537 388922 105603 388925
rect 97276 388920 105603 388922
rect 97276 388864 105542 388920
rect 105598 388864 105603 388920
rect 97276 388862 105603 388864
rect 97276 388860 97282 388862
rect 105537 388859 105603 388862
rect 247033 388922 247099 388925
rect 247585 388922 247651 388925
rect 273897 388922 273963 388925
rect 247033 388920 273963 388922
rect 247033 388864 247038 388920
rect 247094 388864 247590 388920
rect 247646 388864 273902 388920
rect 273958 388864 273963 388920
rect 247033 388862 273963 388864
rect 247033 388859 247099 388862
rect 247585 388859 247651 388862
rect 273897 388859 273963 388862
rect 74441 388786 74507 388789
rect 167729 388786 167795 388789
rect 74441 388784 171150 388786
rect 74441 388728 74446 388784
rect 74502 388728 167734 388784
rect 167790 388728 171150 388784
rect 74441 388726 171150 388728
rect 74441 388723 74507 388726
rect 167729 388723 167795 388726
rect 122097 388514 122163 388517
rect 125593 388514 125659 388517
rect 122097 388512 125659 388514
rect 122097 388456 122102 388512
rect 122158 388456 125598 388512
rect 125654 388456 125659 388512
rect 122097 388454 125659 388456
rect 171090 388514 171150 388726
rect 201125 388514 201191 388517
rect 171090 388512 201191 388514
rect 171090 388456 201130 388512
rect 201186 388456 201191 388512
rect 171090 388454 201191 388456
rect 122097 388451 122163 388454
rect 125593 388451 125659 388454
rect 201125 388451 201191 388454
rect 51441 388378 51507 388381
rect 79961 388378 80027 388381
rect 51441 388376 80027 388378
rect 51441 388320 51446 388376
rect 51502 388320 79966 388376
rect 80022 388320 80027 388376
rect 51441 388318 80027 388320
rect 51441 388315 51507 388318
rect 79961 388315 80027 388318
rect 82997 388378 83063 388381
rect 173065 388378 173131 388381
rect 177297 388378 177363 388381
rect 213453 388378 213519 388381
rect 82997 388376 161490 388378
rect 82997 388320 83002 388376
rect 83058 388320 161490 388376
rect 82997 388318 161490 388320
rect 82997 388315 83063 388318
rect 161430 388242 161490 388318
rect 173065 388376 177363 388378
rect 173065 388320 173070 388376
rect 173126 388320 177302 388376
rect 177358 388320 177363 388376
rect 173065 388318 177363 388320
rect 173065 388315 173131 388318
rect 177297 388315 177363 388318
rect 180750 388376 213519 388378
rect 180750 388320 213458 388376
rect 213514 388320 213519 388376
rect 180750 388318 213519 388320
rect 180241 388242 180307 388245
rect 180750 388242 180810 388318
rect 213453 388315 213519 388318
rect 228357 388378 228423 388381
rect 238109 388378 238175 388381
rect 228357 388376 238175 388378
rect 228357 388320 228362 388376
rect 228418 388320 238114 388376
rect 238170 388320 238175 388376
rect 228357 388318 238175 388320
rect 228357 388315 228423 388318
rect 238109 388315 238175 388318
rect 161430 388240 180810 388242
rect 161430 388184 180246 388240
rect 180302 388184 180810 388240
rect 161430 388182 180810 388184
rect 180241 388179 180307 388182
rect 116669 388106 116735 388109
rect 121453 388106 121519 388109
rect 116669 388104 121519 388106
rect 116669 388048 116674 388104
rect 116730 388048 121458 388104
rect 121514 388048 121519 388104
rect 116669 388046 121519 388048
rect 116669 388043 116735 388046
rect 121453 388043 121519 388046
rect 91093 387834 91159 387837
rect 91318 387834 91324 387836
rect 91093 387832 91324 387834
rect 91093 387776 91098 387832
rect 91154 387776 91324 387832
rect 91093 387774 91324 387776
rect 91093 387771 91159 387774
rect 91318 387772 91324 387774
rect 91388 387772 91394 387836
rect 128353 387834 128419 387837
rect 128997 387834 129063 387837
rect 170489 387834 170555 387837
rect 128353 387832 170555 387834
rect 128353 387776 128358 387832
rect 128414 387776 129002 387832
rect 129058 387776 170494 387832
rect 170550 387776 170555 387832
rect 128353 387774 170555 387776
rect 128353 387771 128419 387774
rect 128997 387771 129063 387774
rect 170489 387771 170555 387774
rect 205541 387834 205607 387837
rect 206829 387834 206895 387837
rect 205541 387832 206895 387834
rect 205541 387776 205546 387832
rect 205602 387776 206834 387832
rect 206890 387776 206895 387832
rect 205541 387774 206895 387776
rect 205541 387771 205607 387774
rect 206829 387771 206895 387774
rect 214557 387834 214623 387837
rect 218237 387834 218303 387837
rect 214557 387832 218303 387834
rect 214557 387776 214562 387832
rect 214618 387776 218242 387832
rect 218298 387776 218303 387832
rect 214557 387774 218303 387776
rect 214557 387771 214623 387774
rect 218237 387771 218303 387774
rect 129733 387698 129799 387701
rect 130469 387698 130535 387701
rect 122790 387696 130535 387698
rect 122790 387640 129738 387696
rect 129794 387640 130474 387696
rect 130530 387640 130535 387696
rect 122790 387638 130535 387640
rect 98913 387562 98979 387565
rect 122790 387562 122850 387638
rect 129733 387635 129799 387638
rect 130469 387635 130535 387638
rect 187049 387698 187115 387701
rect 288617 387698 288683 387701
rect 187049 387696 288683 387698
rect 187049 387640 187054 387696
rect 187110 387640 288622 387696
rect 288678 387640 288683 387696
rect 187049 387638 288683 387640
rect 187049 387635 187115 387638
rect 288617 387635 288683 387638
rect 98913 387560 122850 387562
rect 98913 387504 98918 387560
rect 98974 387504 122850 387560
rect 98913 387502 122850 387504
rect 173157 387562 173223 387565
rect 269297 387562 269363 387565
rect 269430 387562 269436 387564
rect 173157 387560 269436 387562
rect 173157 387504 173162 387560
rect 173218 387504 269302 387560
rect 269358 387504 269436 387560
rect 173157 387502 269436 387504
rect 98913 387499 98979 387502
rect 173157 387499 173223 387502
rect 269297 387499 269363 387502
rect 269430 387500 269436 387502
rect 269500 387500 269506 387564
rect 86861 387426 86927 387429
rect 116669 387426 116735 387429
rect 86861 387424 116735 387426
rect 86861 387368 86866 387424
rect 86922 387368 116674 387424
rect 116730 387368 116735 387424
rect 86861 387366 116735 387368
rect 86861 387363 86927 387366
rect 116669 387363 116735 387366
rect 67357 387290 67423 387293
rect 188521 387290 188587 387293
rect 67357 387288 188587 387290
rect 67357 387232 67362 387288
rect 67418 387232 188526 387288
rect 188582 387232 188587 387288
rect 67357 387230 188587 387232
rect 67357 387227 67423 387230
rect 188521 387227 188587 387230
rect 79317 387018 79383 387021
rect 87454 387018 87460 387020
rect 79317 387016 87460 387018
rect 79317 386960 79322 387016
rect 79378 386960 87460 387016
rect 79317 386958 87460 386960
rect 79317 386955 79383 386958
rect 87454 386956 87460 386958
rect 87524 386956 87530 387020
rect 77201 386338 77267 386341
rect 128353 386338 128419 386341
rect 77201 386336 128419 386338
rect 77201 386280 77206 386336
rect 77262 386280 128358 386336
rect 128414 386280 128419 386336
rect 77201 386278 128419 386280
rect 77201 386275 77267 386278
rect 128353 386275 128419 386278
rect 231117 386338 231183 386341
rect 234245 386338 234311 386341
rect 231117 386336 234311 386338
rect 231117 386280 231122 386336
rect 231178 386280 234250 386336
rect 234306 386280 234311 386336
rect 231117 386278 234311 386280
rect 231117 386275 231183 386278
rect 234245 386275 234311 386278
rect 75821 386202 75887 386205
rect 81934 386202 81940 386204
rect 75821 386200 81940 386202
rect 75821 386144 75826 386200
rect 75882 386144 81940 386200
rect 75821 386142 81940 386144
rect 75821 386139 75887 386142
rect 81934 386140 81940 386142
rect 82004 386140 82010 386204
rect 115974 386202 115980 386204
rect 84150 386142 115980 386202
rect 59077 385658 59143 385661
rect 80421 385658 80487 385661
rect 84150 385658 84210 386142
rect 115974 386140 115980 386142
rect 116044 386140 116050 386204
rect 100845 385794 100911 385797
rect 188429 385794 188495 385797
rect 200205 385794 200271 385797
rect 100845 385792 103530 385794
rect 100845 385736 100850 385792
rect 100906 385736 103530 385792
rect 100845 385734 103530 385736
rect 100845 385731 100911 385734
rect 59077 385656 84210 385658
rect 59077 385600 59082 385656
rect 59138 385600 80426 385656
rect 80482 385600 84210 385656
rect 59077 385598 84210 385600
rect 89621 385658 89687 385661
rect 100702 385658 100708 385660
rect 89621 385656 100708 385658
rect 89621 385600 89626 385656
rect 89682 385600 100708 385656
rect 89621 385598 100708 385600
rect 59077 385595 59143 385598
rect 80421 385595 80487 385598
rect 89621 385595 89687 385598
rect 100702 385596 100708 385598
rect 100772 385596 100778 385660
rect 103470 385658 103530 385734
rect 188429 385792 200271 385794
rect 188429 385736 188434 385792
rect 188490 385736 200210 385792
rect 200266 385736 200271 385792
rect 188429 385734 200271 385736
rect 188429 385731 188495 385734
rect 200205 385731 200271 385734
rect 234613 385658 234679 385661
rect 103470 385656 234679 385658
rect 103470 385600 234618 385656
rect 234674 385600 234679 385656
rect 103470 385598 234679 385600
rect 234613 385595 234679 385598
rect 242893 385658 242959 385661
rect 258390 385658 258396 385660
rect 242893 385656 258396 385658
rect 242893 385600 242898 385656
rect 242954 385600 258396 385656
rect 242893 385598 258396 385600
rect 242893 385595 242959 385598
rect 258390 385596 258396 385598
rect 258460 385596 258466 385660
rect 197353 385114 197419 385117
rect 289905 385114 289971 385117
rect 197353 385112 289971 385114
rect 197353 385056 197358 385112
rect 197414 385056 289910 385112
rect 289966 385056 289971 385112
rect 197353 385054 289971 385056
rect 197353 385051 197419 385054
rect 289905 385051 289971 385054
rect 109677 384978 109743 384981
rect 124213 384978 124279 384981
rect 249057 384978 249123 384981
rect 249517 384978 249583 384981
rect 109677 384976 249583 384978
rect 109677 384920 109682 384976
rect 109738 384920 124218 384976
rect 124274 384920 249062 384976
rect 249118 384920 249522 384976
rect 249578 384920 249583 384976
rect 109677 384918 249583 384920
rect 109677 384915 109743 384918
rect 124213 384915 124279 384918
rect 249057 384915 249123 384918
rect 249517 384915 249583 384918
rect -960 384284 480 384524
rect 83457 384298 83523 384301
rect 90030 384298 90036 384300
rect 83457 384296 90036 384298
rect 83457 384240 83462 384296
rect 83518 384240 90036 384296
rect 83457 384238 90036 384240
rect 83457 384235 83523 384238
rect 90030 384236 90036 384238
rect 90100 384236 90106 384300
rect 101254 384236 101260 384300
rect 101324 384298 101330 384300
rect 113357 384298 113423 384301
rect 101324 384296 113423 384298
rect 101324 384240 113362 384296
rect 113418 384240 113423 384296
rect 101324 384238 113423 384240
rect 101324 384236 101330 384238
rect 113357 384235 113423 384238
rect 91001 383754 91067 383757
rect 94630 383754 94636 383756
rect 91001 383752 94636 383754
rect 91001 383696 91006 383752
rect 91062 383696 94636 383752
rect 91001 383694 94636 383696
rect 91001 383691 91067 383694
rect 94630 383692 94636 383694
rect 94700 383692 94706 383756
rect 73061 383618 73127 383621
rect 197353 383618 197419 383621
rect 73061 383616 197419 383618
rect 73061 383560 73066 383616
rect 73122 383560 197358 383616
rect 197414 383560 197419 383616
rect 73061 383558 197419 383560
rect 73061 383555 73127 383558
rect 197353 383555 197419 383558
rect 187141 383482 187207 383485
rect 273345 383482 273411 383485
rect 187141 383480 273411 383482
rect 187141 383424 187146 383480
rect 187202 383424 273350 383480
rect 273406 383424 273411 383480
rect 187141 383422 273411 383424
rect 187141 383419 187207 383422
rect 273345 383419 273411 383422
rect 81014 382876 81020 382940
rect 81084 382938 81090 382940
rect 88977 382938 89043 382941
rect 81084 382936 89043 382938
rect 81084 382880 88982 382936
rect 89038 382880 89043 382936
rect 81084 382878 89043 382880
rect 81084 382876 81090 382878
rect 88977 382875 89043 382878
rect 79869 382258 79935 382261
rect 173065 382258 173131 382261
rect 79869 382256 173131 382258
rect 79869 382200 79874 382256
rect 79930 382200 173070 382256
rect 173126 382200 173131 382256
rect 79869 382198 173131 382200
rect 79869 382195 79935 382198
rect 173065 382195 173131 382198
rect 180149 382258 180215 382261
rect 266445 382258 266511 382261
rect 180149 382256 266511 382258
rect 180149 382200 180154 382256
rect 180210 382200 266450 382256
rect 266506 382200 266511 382256
rect 180149 382198 266511 382200
rect 180149 382195 180215 382198
rect 266445 382195 266511 382198
rect 55121 382122 55187 382125
rect 103697 382122 103763 382125
rect 104249 382122 104315 382125
rect 55121 382120 104315 382122
rect 55121 382064 55126 382120
rect 55182 382064 103702 382120
rect 103758 382064 104254 382120
rect 104310 382064 104315 382120
rect 55121 382062 104315 382064
rect 55121 382059 55187 382062
rect 103697 382059 103763 382062
rect 104249 382059 104315 382062
rect 195830 381516 195836 381580
rect 195900 381578 195906 381580
rect 204345 381578 204411 381581
rect 195900 381576 204411 381578
rect 195900 381520 204350 381576
rect 204406 381520 204411 381576
rect 195900 381518 204411 381520
rect 195900 381516 195906 381518
rect 204345 381515 204411 381518
rect 72509 380898 72575 380901
rect 72509 380896 180810 380898
rect 72509 380840 72514 380896
rect 72570 380840 180810 380896
rect 72509 380838 180810 380840
rect 72509 380835 72575 380838
rect 180750 380762 180810 380838
rect 197118 380836 197124 380900
rect 197188 380898 197194 380900
rect 200205 380898 200271 380901
rect 260833 380898 260899 380901
rect 261661 380898 261727 380901
rect 197188 380838 200130 380898
rect 197188 380836 197194 380838
rect 198733 380762 198799 380765
rect 180750 380760 198799 380762
rect 180750 380704 198738 380760
rect 198794 380704 198799 380760
rect 180750 380702 198799 380704
rect 200070 380762 200130 380838
rect 200205 380896 261727 380898
rect 200205 380840 200210 380896
rect 200266 380840 260838 380896
rect 260894 380840 261666 380896
rect 261722 380840 261727 380896
rect 200205 380838 261727 380840
rect 200205 380835 200271 380838
rect 260833 380835 260899 380838
rect 261661 380835 261727 380838
rect 202137 380762 202203 380765
rect 200070 380760 202203 380762
rect 200070 380704 202142 380760
rect 202198 380704 202203 380760
rect 200070 380702 202203 380704
rect 198733 380699 198799 380702
rect 202137 380699 202203 380702
rect 168373 380218 168439 380221
rect 169109 380218 169175 380221
rect 200113 380218 200179 380221
rect 168373 380216 200179 380218
rect 168373 380160 168378 380216
rect 168434 380160 169114 380216
rect 169170 380160 200118 380216
rect 200174 380160 200179 380216
rect 168373 380158 200179 380160
rect 168373 380155 168439 380158
rect 169109 380155 169175 380158
rect 200113 380155 200179 380158
rect 234613 380218 234679 380221
rect 274582 380218 274588 380220
rect 234613 380216 274588 380218
rect 234613 380160 234618 380216
rect 234674 380160 274588 380216
rect 234613 380158 274588 380160
rect 234613 380155 234679 380158
rect 274582 380156 274588 380158
rect 274652 380218 274658 380220
rect 274725 380218 274791 380221
rect 274652 380216 274791 380218
rect 274652 380160 274730 380216
rect 274786 380160 274791 380216
rect 274652 380158 274791 380160
rect 274652 380156 274658 380158
rect 274725 380155 274791 380158
rect 50797 379402 50863 379405
rect 178677 379402 178743 379405
rect 50797 379400 178743 379402
rect 50797 379344 50802 379400
rect 50858 379344 178682 379400
rect 178738 379344 178743 379400
rect 50797 379342 178743 379344
rect 50797 379339 50863 379342
rect 178677 379339 178743 379342
rect 191598 379340 191604 379404
rect 191668 379402 191674 379404
rect 583017 379402 583083 379405
rect 191668 379400 583083 379402
rect 191668 379344 583022 379400
rect 583078 379344 583083 379400
rect 191668 379342 583083 379344
rect 191668 379340 191674 379342
rect 583017 379339 583083 379342
rect 261661 379266 261727 379269
rect 266302 379266 266308 379268
rect 261661 379264 266308 379266
rect 261661 379208 261666 379264
rect 261722 379208 266308 379264
rect 261661 379206 266308 379208
rect 261661 379203 261727 379206
rect 266302 379204 266308 379206
rect 266372 379204 266378 379268
rect 191598 378932 191604 378996
rect 191668 378994 191674 378996
rect 191741 378994 191807 378997
rect 191668 378992 191807 378994
rect 191668 378936 191746 378992
rect 191802 378936 191807 378992
rect 191668 378934 191807 378936
rect 191668 378932 191674 378934
rect 191741 378931 191807 378934
rect 85021 378722 85087 378725
rect 96654 378722 96660 378724
rect 85021 378720 96660 378722
rect 85021 378664 85026 378720
rect 85082 378664 96660 378720
rect 85021 378662 96660 378664
rect 85021 378659 85087 378662
rect 96654 378660 96660 378662
rect 96724 378660 96730 378724
rect 582557 378450 582623 378453
rect 583520 378450 584960 378540
rect 582557 378448 584960 378450
rect 582557 378392 582562 378448
rect 582618 378392 584960 378448
rect 582557 378390 584960 378392
rect 582557 378387 582623 378390
rect 583520 378300 584960 378390
rect 48129 378042 48195 378045
rect 130377 378042 130443 378045
rect 48129 378040 130443 378042
rect 48129 377984 48134 378040
rect 48190 377984 130382 378040
rect 130438 377984 130443 378040
rect 48129 377982 130443 377984
rect 48129 377979 48195 377982
rect 130377 377979 130443 377982
rect 151077 378042 151143 378045
rect 265065 378042 265131 378045
rect 265750 378042 265756 378044
rect 151077 378040 265756 378042
rect 151077 377984 151082 378040
rect 151138 377984 265070 378040
rect 265126 377984 265756 378040
rect 151077 377982 265756 377984
rect 151077 377979 151143 377982
rect 265065 377979 265131 377982
rect 265750 377980 265756 377982
rect 265820 377980 265826 378044
rect 119429 377362 119495 377365
rect 255814 377362 255820 377364
rect 119429 377360 255820 377362
rect 119429 377304 119434 377360
rect 119490 377304 255820 377360
rect 119429 377302 255820 377304
rect 119429 377299 119495 377302
rect 255814 377300 255820 377302
rect 255884 377362 255890 377364
rect 258257 377362 258323 377365
rect 255884 377360 258323 377362
rect 255884 377304 258262 377360
rect 258318 377304 258323 377360
rect 255884 377302 258323 377304
rect 255884 377300 255890 377302
rect 258257 377299 258323 377302
rect 148409 376002 148475 376005
rect 255681 376002 255747 376005
rect 148409 376000 255747 376002
rect 148409 375944 148414 376000
rect 148470 375944 255686 376000
rect 255742 375944 255747 376000
rect 148409 375942 255747 375944
rect 148409 375939 148475 375942
rect 255681 375939 255747 375942
rect 69606 375260 69612 375324
rect 69676 375322 69682 375324
rect 157977 375322 158043 375325
rect 69676 375320 158043 375322
rect 69676 375264 157982 375320
rect 158038 375264 158043 375320
rect 69676 375262 158043 375264
rect 69676 375260 69682 375262
rect 157977 375259 158043 375262
rect 188521 375322 188587 375325
rect 279417 375322 279483 375325
rect 188521 375320 279483 375322
rect 188521 375264 188526 375320
rect 188582 375264 279422 375320
rect 279478 375264 279483 375320
rect 188521 375262 279483 375264
rect 188521 375259 188587 375262
rect 279417 375259 279483 375262
rect 65885 373962 65951 373965
rect 188838 373962 188844 373964
rect 65885 373960 188844 373962
rect 65885 373904 65890 373960
rect 65946 373904 188844 373960
rect 65885 373902 188844 373904
rect 65885 373899 65951 373902
rect 188838 373900 188844 373902
rect 188908 373900 188914 373964
rect 72417 373282 72483 373285
rect 77334 373282 77340 373284
rect 72417 373280 77340 373282
rect 72417 373224 72422 373280
rect 72478 373224 77340 373280
rect 72417 373222 77340 373224
rect 72417 373219 72483 373222
rect 77334 373220 77340 373222
rect 77404 373220 77410 373284
rect 191741 373282 191807 373285
rect 252502 373282 252508 373284
rect 191741 373280 252508 373282
rect 191741 373224 191746 373280
rect 191802 373224 252508 373280
rect 191741 373222 252508 373224
rect 191741 373219 191807 373222
rect 252502 373220 252508 373222
rect 252572 373220 252578 373284
rect 188838 372812 188844 372876
rect 188908 372874 188914 372876
rect 191741 372874 191807 372877
rect 188908 372872 191807 372874
rect 188908 372816 191746 372872
rect 191802 372816 191807 372872
rect 188908 372814 191807 372816
rect 188908 372812 188914 372814
rect 191741 372811 191807 372814
rect 67909 372602 67975 372605
rect 160737 372602 160803 372605
rect 67909 372600 160803 372602
rect 67909 372544 67914 372600
rect 67970 372544 160742 372600
rect 160798 372544 160803 372600
rect 67909 372542 160803 372544
rect 67909 372539 67975 372542
rect 160737 372539 160803 372542
rect 170489 372058 170555 372061
rect 171041 372058 171107 372061
rect 204253 372058 204319 372061
rect 170489 372056 204319 372058
rect 170489 372000 170494 372056
rect 170550 372000 171046 372056
rect 171102 372000 204258 372056
rect 204314 372000 204319 372056
rect 170489 371998 204319 372000
rect 170489 371995 170555 371998
rect 171041 371995 171107 371998
rect 204253 371995 204319 371998
rect 193806 371860 193812 371924
rect 193876 371922 193882 371924
rect 242157 371922 242223 371925
rect 193876 371920 242223 371922
rect 193876 371864 242162 371920
rect 242218 371864 242223 371920
rect 193876 371862 242223 371864
rect 193876 371860 193882 371862
rect 242157 371859 242223 371862
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 160185 371378 160251 371381
rect 160737 371378 160803 371381
rect 160185 371376 160803 371378
rect 160185 371320 160190 371376
rect 160246 371320 160742 371376
rect 160798 371320 160803 371376
rect 160185 371318 160803 371320
rect 160185 371315 160251 371318
rect 160737 371315 160803 371318
rect 242014 371316 242020 371380
rect 242084 371378 242090 371380
rect 244917 371378 244983 371381
rect 242084 371376 244983 371378
rect 242084 371320 244922 371376
rect 244978 371320 244983 371376
rect 242084 371318 244983 371320
rect 242084 371316 242090 371318
rect 244917 371315 244983 371318
rect 67817 371242 67883 371245
rect 159541 371242 159607 371245
rect 67817 371240 159607 371242
rect 67817 371184 67822 371240
rect 67878 371184 159546 371240
rect 159602 371184 159607 371240
rect 67817 371182 159607 371184
rect 67817 371179 67883 371182
rect 159541 371179 159607 371182
rect 193121 370562 193187 370565
rect 242985 370562 243051 370565
rect 193121 370560 243051 370562
rect 193121 370504 193126 370560
rect 193182 370504 242990 370560
rect 243046 370504 243051 370560
rect 193121 370502 243051 370504
rect 193121 370499 193187 370502
rect 242985 370499 243051 370502
rect 243537 370562 243603 370565
rect 260833 370562 260899 370565
rect 243537 370560 260899 370562
rect 243537 370504 243542 370560
rect 243598 370504 260838 370560
rect 260894 370504 260899 370560
rect 243537 370502 260899 370504
rect 243537 370499 243603 370502
rect 260833 370499 260899 370502
rect 66662 369684 66668 369748
rect 66732 369746 66738 369748
rect 159357 369746 159423 369749
rect 66732 369744 159423 369746
rect 66732 369688 159362 369744
rect 159418 369688 159423 369744
rect 66732 369686 159423 369688
rect 66732 369684 66738 369686
rect 159357 369683 159423 369686
rect 169201 369746 169267 369749
rect 255998 369746 256004 369748
rect 169201 369744 256004 369746
rect 169201 369688 169206 369744
rect 169262 369688 256004 369744
rect 169201 369686 256004 369688
rect 169201 369683 169267 369686
rect 255998 369684 256004 369686
rect 256068 369746 256074 369748
rect 256068 369686 258090 369746
rect 256068 369684 256074 369686
rect 258030 369066 258090 369686
rect 273294 369066 273300 369068
rect 258030 369006 273300 369066
rect 273294 369004 273300 369006
rect 273364 369004 273370 369068
rect 191741 367706 191807 367709
rect 254577 367706 254643 367709
rect 191741 367704 254643 367706
rect 191741 367648 191746 367704
rect 191802 367648 254582 367704
rect 254638 367648 254643 367704
rect 191741 367646 254643 367648
rect 191741 367643 191807 367646
rect 254577 367643 254643 367646
rect 238661 366482 238727 366485
rect 241646 366482 241652 366484
rect 238661 366480 241652 366482
rect 238661 366424 238666 366480
rect 238722 366424 241652 366480
rect 238661 366422 241652 366424
rect 238661 366419 238727 366422
rect 241646 366420 241652 366422
rect 241716 366420 241722 366484
rect 233877 366346 233943 366349
rect 252686 366346 252692 366348
rect 233877 366344 252692 366346
rect 233877 366288 233882 366344
rect 233938 366288 252692 366344
rect 233877 366286 252692 366288
rect 233877 366283 233943 366286
rect 252686 366284 252692 366286
rect 252756 366284 252762 366348
rect 181345 365802 181411 365805
rect 220721 365802 220787 365805
rect 181345 365800 220787 365802
rect 181345 365744 181350 365800
rect 181406 365744 220726 365800
rect 220782 365744 220787 365800
rect 181345 365742 220787 365744
rect 181345 365739 181411 365742
rect 220721 365739 220787 365742
rect 214557 365666 214623 365669
rect 215201 365666 215267 365669
rect 214557 365664 215267 365666
rect 214557 365608 214562 365664
rect 214618 365608 215206 365664
rect 215262 365608 215267 365664
rect 214557 365606 215267 365608
rect 214557 365603 214623 365606
rect 215201 365603 215267 365606
rect 582465 365122 582531 365125
rect 583520 365122 584960 365212
rect 582465 365120 584960 365122
rect 582465 365064 582470 365120
rect 582526 365064 584960 365120
rect 582465 365062 584960 365064
rect 582465 365059 582531 365062
rect 116669 364986 116735 364989
rect 215201 364986 215267 364989
rect 116669 364984 215267 364986
rect 116669 364928 116674 364984
rect 116730 364928 215206 364984
rect 215262 364928 215267 364984
rect 583520 364972 584960 365062
rect 116669 364926 215267 364928
rect 116669 364923 116735 364926
rect 215201 364923 215267 364926
rect 104249 363626 104315 363629
rect 213821 363626 213887 363629
rect 104249 363624 213887 363626
rect 104249 363568 104254 363624
rect 104310 363568 213826 363624
rect 213882 363568 213887 363624
rect 104249 363566 213887 363568
rect 104249 363563 104315 363566
rect 213821 363563 213887 363566
rect 215201 363626 215267 363629
rect 267774 363626 267780 363628
rect 215201 363624 267780 363626
rect 215201 363568 215206 363624
rect 215262 363568 267780 363624
rect 215201 363566 267780 363568
rect 215201 363563 215267 363566
rect 267774 363564 267780 363566
rect 267844 363564 267850 363628
rect 240041 361722 240107 361725
rect 245694 361722 245700 361724
rect 240041 361720 245700 361722
rect 240041 361664 240046 361720
rect 240102 361664 245700 361720
rect 240041 361662 245700 361664
rect 240041 361659 240107 361662
rect 245694 361660 245700 361662
rect 245764 361660 245770 361724
rect 213821 361586 213887 361589
rect 242249 361586 242315 361589
rect 213821 361584 242315 361586
rect 213821 361528 213826 361584
rect 213882 361528 242254 361584
rect 242310 361528 242315 361584
rect 213821 361526 242315 361528
rect 213821 361523 213887 361526
rect 242249 361523 242315 361526
rect 231117 359410 231183 359413
rect 277158 359410 277164 359412
rect 231117 359408 277164 359410
rect 231117 359352 231122 359408
rect 231178 359352 277164 359408
rect 231117 359350 277164 359352
rect 231117 359347 231183 359350
rect 277158 359348 277164 359350
rect 277228 359348 277234 359412
rect 124857 358730 124923 358733
rect 258390 358730 258396 358732
rect 124857 358728 258396 358730
rect 124857 358672 124862 358728
rect 124918 358672 258396 358728
rect 124857 358670 258396 358672
rect 124857 358667 124923 358670
rect 258390 358668 258396 358670
rect 258460 358668 258466 358732
rect -960 358458 480 358548
rect 2773 358458 2839 358461
rect -960 358456 2839 358458
rect -960 358400 2778 358456
rect 2834 358400 2839 358456
rect -960 358398 2839 358400
rect -960 358308 480 358398
rect 2773 358395 2839 358398
rect 122097 356690 122163 356693
rect 228357 356690 228423 356693
rect 122097 356688 228423 356690
rect 122097 356632 122102 356688
rect 122158 356632 228362 356688
rect 228418 356632 228423 356688
rect 122097 356630 228423 356632
rect 122097 356627 122163 356630
rect 228357 356627 228423 356630
rect 582649 351930 582715 351933
rect 583520 351930 584960 352020
rect 582649 351928 584960 351930
rect 582649 351872 582654 351928
rect 582710 351872 584960 351928
rect 582649 351870 584960 351872
rect 582649 351867 582715 351870
rect 583520 351780 584960 351870
rect 135989 347850 136055 347853
rect 263685 347850 263751 347853
rect 135989 347848 263751 347850
rect 135989 347792 135994 347848
rect 136050 347792 263690 347848
rect 263746 347792 263751 347848
rect 135989 347790 263751 347792
rect 135989 347787 136055 347790
rect 263685 347787 263751 347790
rect 191598 346972 191604 347036
rect 191668 347034 191674 347036
rect 253933 347034 253999 347037
rect 191668 347032 253999 347034
rect 191668 346976 253938 347032
rect 253994 346976 253999 347032
rect 191668 346974 253999 346976
rect 191668 346972 191674 346974
rect 253933 346971 253999 346974
rect 205541 345674 205607 345677
rect 250294 345674 250300 345676
rect 205541 345672 250300 345674
rect 205541 345616 205546 345672
rect 205602 345616 250300 345672
rect 205541 345614 250300 345616
rect 205541 345611 205607 345614
rect 250294 345612 250300 345614
rect 250364 345612 250370 345676
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 202137 344314 202203 344317
rect 241646 344314 241652 344316
rect 202137 344312 241652 344314
rect 202137 344256 202142 344312
rect 202198 344256 241652 344312
rect 202137 344254 241652 344256
rect 202137 344251 202203 344254
rect 241646 344252 241652 344254
rect 241716 344252 241722 344316
rect 148409 342274 148475 342277
rect 231209 342274 231275 342277
rect 148409 342272 231275 342274
rect 148409 342216 148414 342272
rect 148470 342216 231214 342272
rect 231270 342216 231275 342272
rect 148409 342214 231275 342216
rect 148409 342211 148475 342214
rect 231209 342211 231275 342214
rect 47577 340914 47643 340917
rect 205633 340914 205699 340917
rect 47577 340912 205699 340914
rect 47577 340856 47582 340912
rect 47638 340856 205638 340912
rect 205694 340856 205699 340912
rect 47577 340854 205699 340856
rect 47577 340851 47643 340854
rect 205633 340851 205699 340854
rect 48221 339554 48287 339557
rect 205725 339554 205791 339557
rect 48221 339552 205791 339554
rect 48221 339496 48226 339552
rect 48282 339496 205730 339552
rect 205786 339496 205791 339552
rect 48221 339494 205791 339496
rect 48221 339491 48287 339494
rect 205725 339491 205791 339494
rect 184197 338738 184263 338741
rect 269246 338738 269252 338740
rect 184197 338736 269252 338738
rect 184197 338680 184202 338736
rect 184258 338680 269252 338736
rect 184197 338678 269252 338680
rect 184197 338675 184263 338678
rect 269246 338676 269252 338678
rect 269316 338676 269322 338740
rect 583520 338452 584960 338692
rect 128997 336834 129063 336837
rect 227713 336834 227779 336837
rect 128997 336832 227779 336834
rect 128997 336776 129002 336832
rect 129058 336776 227718 336832
rect 227774 336776 227779 336832
rect 128997 336774 227779 336776
rect 128997 336771 129063 336774
rect 227713 336771 227779 336774
rect 31661 335474 31727 335477
rect 222285 335474 222351 335477
rect 31661 335472 222351 335474
rect 31661 335416 31666 335472
rect 31722 335416 222290 335472
rect 222346 335416 222351 335472
rect 31661 335414 222351 335416
rect 31661 335411 31727 335414
rect 222285 335411 222351 335414
rect 35801 334114 35867 334117
rect 213177 334114 213243 334117
rect 35801 334112 213243 334114
rect 35801 334056 35806 334112
rect 35862 334056 213182 334112
rect 213238 334056 213243 334112
rect 35801 334054 213243 334056
rect 35801 334051 35867 334054
rect 213177 334051 213243 334054
rect 221549 333298 221615 333301
rect 260925 333298 260991 333301
rect 221549 333296 260991 333298
rect 221549 333240 221554 333296
rect 221610 333240 260930 333296
rect 260986 333240 260991 333296
rect 221549 333238 260991 333240
rect 221549 333235 221615 333238
rect 260925 333235 260991 333238
rect 13721 332618 13787 332621
rect 219433 332618 219499 332621
rect 13721 332616 219499 332618
rect 13721 332560 13726 332616
rect 13782 332560 219438 332616
rect 219494 332560 219499 332616
rect 13721 332558 219499 332560
rect 13721 332555 13787 332558
rect 219433 332555 219499 332558
rect -960 332196 480 332436
rect 122189 331394 122255 331397
rect 228449 331394 228515 331397
rect 122189 331392 228515 331394
rect 122189 331336 122194 331392
rect 122250 331336 228454 331392
rect 228510 331336 228515 331392
rect 122189 331334 228515 331336
rect 122189 331331 122255 331334
rect 228449 331331 228515 331334
rect 34421 331258 34487 331261
rect 199377 331258 199443 331261
rect 34421 331256 199443 331258
rect 34421 331200 34426 331256
rect 34482 331200 199382 331256
rect 199438 331200 199443 331256
rect 34421 331198 199443 331200
rect 34421 331195 34487 331198
rect 199377 331195 199443 331198
rect 220077 330442 220143 330445
rect 253933 330442 253999 330445
rect 220077 330440 253999 330442
rect 220077 330384 220082 330440
rect 220138 330384 253938 330440
rect 253994 330384 253999 330440
rect 220077 330382 253999 330384
rect 220077 330379 220143 330382
rect 253933 330379 253999 330382
rect 127617 330034 127683 330037
rect 213269 330034 213335 330037
rect 127617 330032 213335 330034
rect 127617 329976 127622 330032
rect 127678 329976 213274 330032
rect 213330 329976 213335 330032
rect 127617 329974 213335 329976
rect 127617 329971 127683 329974
rect 213269 329971 213335 329974
rect 22001 329898 22067 329901
rect 201677 329898 201743 329901
rect 22001 329896 201743 329898
rect 22001 329840 22006 329896
rect 22062 329840 201682 329896
rect 201738 329840 201743 329896
rect 22001 329838 201743 329840
rect 22001 329835 22067 329838
rect 201677 329835 201743 329838
rect 93761 329082 93827 329085
rect 102726 329082 102732 329084
rect 93761 329080 102732 329082
rect 93761 329024 93766 329080
rect 93822 329024 102732 329080
rect 93761 329022 102732 329024
rect 93761 329019 93827 329022
rect 102726 329020 102732 329022
rect 102796 329020 102802 329084
rect 184381 328674 184447 328677
rect 258717 328674 258783 328677
rect 184381 328672 258783 328674
rect 184381 328616 184386 328672
rect 184442 328616 258722 328672
rect 258778 328616 258783 328672
rect 184381 328614 258783 328616
rect 184381 328611 184447 328614
rect 258717 328611 258783 328614
rect 147029 328538 147095 328541
rect 225137 328538 225203 328541
rect 147029 328536 225203 328538
rect 147029 328480 147034 328536
rect 147090 328480 225142 328536
rect 225198 328480 225203 328536
rect 147029 328478 225203 328480
rect 147029 328475 147095 328478
rect 225137 328475 225203 328478
rect 254526 328340 254532 328404
rect 254596 328402 254602 328404
rect 254761 328402 254827 328405
rect 254596 328400 254827 328402
rect 254596 328344 254766 328400
rect 254822 328344 254827 328400
rect 254596 328342 254827 328344
rect 254596 328340 254602 328342
rect 254761 328339 254827 328342
rect 158069 327722 158135 327725
rect 188889 327722 188955 327725
rect 246389 327722 246455 327725
rect 158069 327720 246455 327722
rect 158069 327664 158074 327720
rect 158130 327664 188894 327720
rect 188950 327664 246394 327720
rect 246450 327664 246455 327720
rect 158069 327662 246455 327664
rect 158069 327659 158135 327662
rect 188889 327659 188955 327662
rect 246389 327659 246455 327662
rect 189073 327314 189139 327317
rect 190361 327314 190427 327317
rect 254761 327314 254827 327317
rect 189073 327312 254827 327314
rect 189073 327256 189078 327312
rect 189134 327256 190366 327312
rect 190422 327256 254766 327312
rect 254822 327256 254827 327312
rect 189073 327254 254827 327256
rect 189073 327251 189139 327254
rect 190361 327251 190427 327254
rect 254761 327251 254827 327254
rect 126329 327178 126395 327181
rect 216029 327178 216095 327181
rect 126329 327176 216095 327178
rect 126329 327120 126334 327176
rect 126390 327120 216034 327176
rect 216090 327120 216095 327176
rect 126329 327118 216095 327120
rect 126329 327115 126395 327118
rect 216029 327115 216095 327118
rect 133137 325954 133203 325957
rect 215937 325954 216003 325957
rect 133137 325952 216003 325954
rect 133137 325896 133142 325952
rect 133198 325896 215942 325952
rect 215998 325896 216003 325952
rect 133137 325894 216003 325896
rect 133137 325891 133203 325894
rect 215937 325891 216003 325894
rect 38561 325818 38627 325821
rect 223665 325818 223731 325821
rect 38561 325816 223731 325818
rect 38561 325760 38566 325816
rect 38622 325760 223670 325816
rect 223726 325760 223731 325816
rect 38561 325758 223731 325760
rect 38561 325755 38627 325758
rect 223665 325755 223731 325758
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect 97257 325002 97323 325005
rect 162761 325002 162827 325005
rect 263869 325002 263935 325005
rect 97257 325000 263935 325002
rect 97257 324944 97262 325000
rect 97318 324944 162766 325000
rect 162822 324944 263874 325000
rect 263930 324944 263935 325000
rect 97257 324942 263935 324944
rect 97257 324939 97323 324942
rect 162761 324939 162827 324942
rect 263869 324939 263935 324942
rect 140129 324458 140195 324461
rect 215845 324458 215911 324461
rect 256877 324458 256943 324461
rect 140129 324456 256943 324458
rect 140129 324400 140134 324456
rect 140190 324400 215850 324456
rect 215906 324400 256882 324456
rect 256938 324400 256943 324456
rect 140129 324398 256943 324400
rect 140129 324395 140195 324398
rect 215845 324395 215911 324398
rect 256877 324395 256943 324398
rect 259453 323644 259519 323645
rect 259453 323642 259500 323644
rect 259408 323640 259500 323642
rect 259408 323584 259458 323640
rect 259408 323582 259500 323584
rect 259453 323580 259500 323582
rect 259564 323580 259570 323644
rect 259453 323579 259519 323580
rect 159357 323098 159423 323101
rect 222929 323098 222995 323101
rect 159357 323096 222995 323098
rect 159357 323040 159362 323096
rect 159418 323040 222934 323096
rect 222990 323040 222995 323096
rect 159357 323038 222995 323040
rect 159357 323035 159423 323038
rect 222929 323035 222995 323038
rect 25497 322962 25563 322965
rect 198825 322962 198891 322965
rect 25497 322960 198891 322962
rect 25497 322904 25502 322960
rect 25558 322904 198830 322960
rect 198886 322904 198891 322960
rect 25497 322902 198891 322904
rect 25497 322899 25563 322902
rect 198825 322899 198891 322902
rect 78581 322826 78647 322829
rect 85798 322826 85804 322828
rect 78581 322824 85804 322826
rect 78581 322768 78586 322824
rect 78642 322768 85804 322824
rect 78581 322766 85804 322768
rect 78581 322763 78647 322766
rect 85798 322764 85804 322766
rect 85868 322764 85874 322828
rect 149789 321738 149855 321741
rect 207105 321738 207171 321741
rect 149789 321736 207171 321738
rect 149789 321680 149794 321736
rect 149850 321680 207110 321736
rect 207166 321680 207171 321736
rect 149789 321678 207171 321680
rect 149789 321675 149855 321678
rect 207105 321675 207171 321678
rect 186957 321602 187023 321605
rect 187601 321602 187667 321605
rect 258809 321602 258875 321605
rect 186957 321600 258875 321602
rect 186957 321544 186962 321600
rect 187018 321544 187606 321600
rect 187662 321544 258814 321600
rect 258870 321544 258875 321600
rect 186957 321542 258875 321544
rect 186957 321539 187023 321542
rect 187601 321539 187667 321542
rect 258809 321539 258875 321542
rect 170489 320378 170555 320381
rect 239397 320378 239463 320381
rect 170489 320376 239463 320378
rect 170489 320320 170494 320376
rect 170550 320320 239402 320376
rect 239458 320320 239463 320376
rect 170489 320318 239463 320320
rect 170489 320315 170555 320318
rect 239397 320315 239463 320318
rect 151077 320242 151143 320245
rect 266353 320242 266419 320245
rect 151077 320240 266419 320242
rect 151077 320184 151082 320240
rect 151138 320184 266358 320240
rect 266414 320184 266419 320240
rect 151077 320182 266419 320184
rect 151077 320179 151143 320182
rect 266353 320179 266419 320182
rect 75913 320106 75979 320109
rect 84694 320106 84700 320108
rect 75913 320104 84700 320106
rect 75913 320048 75918 320104
rect 75974 320048 84700 320104
rect 75913 320046 84700 320048
rect 75913 320043 75979 320046
rect 84694 320044 84700 320046
rect 84764 320106 84770 320108
rect 182081 320106 182147 320109
rect 84764 320104 182147 320106
rect 84764 320048 182086 320104
rect 182142 320048 182147 320104
rect 84764 320046 182147 320048
rect 84764 320044 84770 320046
rect 182081 320043 182147 320046
rect 86861 319426 86927 319429
rect 94446 319426 94452 319428
rect 86861 319424 94452 319426
rect -960 319290 480 319380
rect 86861 319368 86866 319424
rect 86922 319368 94452 319424
rect 86861 319366 94452 319368
rect 86861 319363 86927 319366
rect 94446 319364 94452 319366
rect 94516 319364 94522 319428
rect 95141 319426 95207 319429
rect 105486 319426 105492 319428
rect 95141 319424 105492 319426
rect 95141 319368 95146 319424
rect 95202 319368 105492 319424
rect 95141 319366 105492 319368
rect 95141 319363 95207 319366
rect 105486 319364 105492 319366
rect 105556 319364 105562 319428
rect 151169 319426 151235 319429
rect 258349 319426 258415 319429
rect 259361 319426 259427 319429
rect 151169 319424 259427 319426
rect 151169 319368 151174 319424
rect 151230 319368 258354 319424
rect 258410 319368 259366 319424
rect 259422 319368 259427 319424
rect 151169 319366 259427 319368
rect 151169 319363 151235 319366
rect 258349 319363 258415 319366
rect 259361 319363 259427 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 178953 318882 179019 318885
rect 233325 318882 233391 318885
rect 178953 318880 233391 318882
rect 178953 318824 178958 318880
rect 179014 318824 233330 318880
rect 233386 318824 233391 318880
rect 178953 318822 233391 318824
rect 178953 318819 179019 318822
rect 233325 318819 233391 318822
rect 284293 318746 284359 318749
rect 284569 318746 284635 318749
rect 284293 318744 284635 318746
rect 284293 318688 284298 318744
rect 284354 318688 284574 318744
rect 284630 318688 284635 318744
rect 284293 318686 284635 318688
rect 284293 318683 284359 318686
rect 284569 318683 284635 318686
rect 79961 318066 80027 318069
rect 87086 318066 87092 318068
rect 79961 318064 87092 318066
rect 79961 318008 79966 318064
rect 80022 318008 87092 318064
rect 79961 318006 87092 318008
rect 79961 318003 80027 318006
rect 87086 318004 87092 318006
rect 87156 318004 87162 318068
rect 88149 318066 88215 318069
rect 97942 318066 97948 318068
rect 88149 318064 97948 318066
rect 88149 318008 88154 318064
rect 88210 318008 97948 318064
rect 88149 318006 97948 318008
rect 88149 318003 88215 318006
rect 97942 318004 97948 318006
rect 98012 318004 98018 318068
rect 188470 317732 188476 317796
rect 188540 317794 188546 317796
rect 209037 317794 209103 317797
rect 188540 317792 209103 317794
rect 188540 317736 209042 317792
rect 209098 317736 209103 317792
rect 188540 317734 209103 317736
rect 188540 317732 188546 317734
rect 209037 317731 209103 317734
rect 134609 317658 134675 317661
rect 229921 317658 229987 317661
rect 134609 317656 229987 317658
rect 134609 317600 134614 317656
rect 134670 317600 229926 317656
rect 229982 317600 229987 317656
rect 134609 317598 229987 317600
rect 134609 317595 134675 317598
rect 229921 317595 229987 317598
rect 262857 317658 262923 317661
rect 267958 317658 267964 317660
rect 262857 317656 267964 317658
rect 262857 317600 262862 317656
rect 262918 317600 267964 317656
rect 262857 317598 267964 317600
rect 262857 317595 262923 317598
rect 267958 317596 267964 317598
rect 268028 317596 268034 317660
rect 188337 317522 188403 317525
rect 284569 317522 284635 317525
rect 188337 317520 284635 317522
rect 188337 317464 188342 317520
rect 188398 317464 284574 317520
rect 284630 317464 284635 317520
rect 188337 317462 284635 317464
rect 188337 317459 188403 317462
rect 284569 317459 284635 317462
rect 75177 317386 75243 317389
rect 83038 317386 83044 317388
rect 75177 317384 83044 317386
rect 75177 317328 75182 317384
rect 75238 317328 83044 317384
rect 75177 317326 83044 317328
rect 75177 317323 75243 317326
rect 83038 317324 83044 317326
rect 83108 317324 83114 317388
rect 84510 317324 84516 317388
rect 84580 317386 84586 317388
rect 87045 317386 87111 317389
rect 84580 317384 87111 317386
rect 84580 317328 87050 317384
rect 87106 317328 87111 317384
rect 84580 317326 87111 317328
rect 84580 317324 84586 317326
rect 87045 317323 87111 317326
rect 166257 316298 166323 316301
rect 226977 316298 227043 316301
rect 166257 316296 227043 316298
rect 166257 316240 166262 316296
rect 166318 316240 226982 316296
rect 227038 316240 227043 316296
rect 166257 316238 227043 316240
rect 166257 316235 166323 316238
rect 226977 316235 227043 316238
rect 69289 316162 69355 316165
rect 74574 316162 74580 316164
rect 69289 316160 74580 316162
rect 69289 316104 69294 316160
rect 69350 316104 74580 316160
rect 69289 316102 74580 316104
rect 69289 316099 69355 316102
rect 74574 316100 74580 316102
rect 74644 316100 74650 316164
rect 94497 316162 94563 316165
rect 256693 316162 256759 316165
rect 257429 316162 257495 316165
rect 94497 316160 257495 316162
rect 94497 316104 94502 316160
rect 94558 316104 256698 316160
rect 256754 316104 257434 316160
rect 257490 316104 257495 316160
rect 94497 316102 257495 316104
rect 94497 316099 94563 316102
rect 256693 316099 256759 316102
rect 257429 316099 257495 316102
rect 211797 315346 211863 315349
rect 258390 315346 258396 315348
rect 211797 315344 258396 315346
rect 211797 315288 211802 315344
rect 211858 315288 258396 315344
rect 211797 315286 258396 315288
rect 211797 315283 211863 315286
rect 258390 315284 258396 315286
rect 258460 315284 258466 315348
rect 192569 315074 192635 315077
rect 193213 315074 193279 315077
rect 192569 315072 193279 315074
rect 192569 315016 192574 315072
rect 192630 315016 193218 315072
rect 193274 315016 193279 315072
rect 192569 315014 193279 315016
rect 192569 315011 192635 315014
rect 193213 315011 193279 315014
rect 142797 314938 142863 314941
rect 209773 314938 209839 314941
rect 142797 314936 209839 314938
rect 142797 314880 142802 314936
rect 142858 314880 209778 314936
rect 209834 314880 209839 314936
rect 142797 314878 209839 314880
rect 142797 314875 142863 314878
rect 209773 314875 209839 314878
rect 149697 314802 149763 314805
rect 218697 314802 218763 314805
rect 149697 314800 218763 314802
rect 149697 314744 149702 314800
rect 149758 314744 218702 314800
rect 218758 314744 218763 314800
rect 149697 314742 218763 314744
rect 149697 314739 149763 314742
rect 218697 314739 218763 314742
rect 192661 313986 192727 313989
rect 204345 313986 204411 313989
rect 243077 313986 243143 313989
rect 192661 313984 243143 313986
rect 192661 313928 192666 313984
rect 192722 313928 204350 313984
rect 204406 313928 243082 313984
rect 243138 313928 243143 313984
rect 192661 313926 243143 313928
rect 192661 313923 192727 313926
rect 204345 313923 204411 313926
rect 243077 313923 243143 313926
rect 41321 313442 41387 313445
rect 204713 313442 204779 313445
rect 41321 313440 204779 313442
rect 41321 313384 41326 313440
rect 41382 313384 204718 313440
rect 204774 313384 204779 313440
rect 41321 313382 204779 313384
rect 41321 313379 41387 313382
rect 204713 313379 204779 313382
rect 254761 313442 254827 313445
rect 255497 313442 255563 313445
rect 254761 313440 255563 313442
rect 254761 313384 254766 313440
rect 254822 313384 255502 313440
rect 255558 313384 255563 313440
rect 254761 313382 255563 313384
rect 254761 313379 254827 313382
rect 255497 313379 255563 313382
rect 82905 313306 82971 313309
rect 277393 313306 277459 313309
rect 82905 313304 277459 313306
rect 82905 313248 82910 313304
rect 82966 313248 277398 313304
rect 277454 313248 277459 313304
rect 82905 313246 277459 313248
rect 82905 313243 82971 313246
rect 277393 313243 277459 313246
rect 169201 312218 169267 312221
rect 269297 312218 269363 312221
rect 169201 312216 269363 312218
rect 169201 312160 169206 312216
rect 169262 312160 269302 312216
rect 269358 312160 269363 312216
rect 169201 312158 269363 312160
rect 169201 312155 169267 312158
rect 269297 312155 269363 312158
rect 32397 312082 32463 312085
rect 220905 312082 220971 312085
rect 32397 312080 220971 312082
rect 32397 312024 32402 312080
rect 32458 312024 220910 312080
rect 220966 312024 220971 312080
rect 32397 312022 220971 312024
rect 32397 312019 32463 312022
rect 220905 312019 220971 312022
rect 582649 312082 582715 312085
rect 583520 312082 584960 312172
rect 582649 312080 584960 312082
rect 582649 312024 582654 312080
rect 582710 312024 584960 312080
rect 582649 312022 584960 312024
rect 582649 312019 582715 312022
rect 23381 311946 23447 311949
rect 220997 311946 221063 311949
rect 23381 311944 221063 311946
rect 23381 311888 23386 311944
rect 23442 311888 221002 311944
rect 221058 311888 221063 311944
rect 583520 311932 584960 312022
rect 23381 311886 221063 311888
rect 23381 311883 23447 311886
rect 220997 311883 221063 311886
rect 249057 311266 249123 311269
rect 263542 311266 263548 311268
rect 249057 311264 263548 311266
rect 249057 311208 249062 311264
rect 249118 311208 263548 311264
rect 249057 311206 263548 311208
rect 249057 311203 249123 311206
rect 263542 311204 263548 311206
rect 263612 311204 263618 311268
rect 52177 311130 52243 311133
rect 52361 311130 52427 311133
rect 280286 311130 280292 311132
rect 52177 311128 280292 311130
rect 52177 311072 52182 311128
rect 52238 311072 52366 311128
rect 52422 311072 280292 311128
rect 52177 311070 280292 311072
rect 52177 311067 52243 311070
rect 52361 311067 52427 311070
rect 280286 311068 280292 311070
rect 280356 311130 280362 311132
rect 280797 311130 280863 311133
rect 280356 311128 280863 311130
rect 280356 311072 280802 311128
rect 280858 311072 280863 311128
rect 280356 311070 280863 311072
rect 280356 311068 280362 311070
rect 280797 311067 280863 311070
rect 171777 310722 171843 310725
rect 211429 310722 211495 310725
rect 171777 310720 211495 310722
rect 171777 310664 171782 310720
rect 171838 310664 211434 310720
rect 211490 310664 211495 310720
rect 171777 310662 211495 310664
rect 171777 310659 171843 310662
rect 211429 310659 211495 310662
rect 30281 310586 30347 310589
rect 203057 310586 203123 310589
rect 30281 310584 203123 310586
rect 30281 310528 30286 310584
rect 30342 310528 203062 310584
rect 203118 310528 203123 310584
rect 30281 310526 203123 310528
rect 30281 310523 30347 310526
rect 203057 310523 203123 310526
rect 81341 309906 81407 309909
rect 89662 309906 89668 309908
rect 81341 309904 89668 309906
rect 81341 309848 81346 309904
rect 81402 309848 89668 309904
rect 81341 309846 89668 309848
rect 81341 309843 81407 309846
rect 89662 309844 89668 309846
rect 89732 309844 89738 309908
rect 86769 309770 86835 309773
rect 96286 309770 96292 309772
rect 86769 309768 96292 309770
rect 86769 309712 86774 309768
rect 86830 309712 96292 309768
rect 86769 309710 96292 309712
rect 86769 309707 86835 309710
rect 96286 309708 96292 309710
rect 96356 309708 96362 309772
rect 96521 309770 96587 309773
rect 108982 309770 108988 309772
rect 96521 309768 108988 309770
rect 96521 309712 96526 309768
rect 96582 309712 108988 309768
rect 96521 309710 108988 309712
rect 96521 309707 96587 309710
rect 108982 309708 108988 309710
rect 109052 309708 109058 309772
rect 227069 309770 227135 309773
rect 260966 309770 260972 309772
rect 227069 309768 260972 309770
rect 227069 309712 227074 309768
rect 227130 309712 260972 309768
rect 227069 309710 260972 309712
rect 227069 309707 227135 309710
rect 260966 309708 260972 309710
rect 261036 309708 261042 309772
rect 173249 309498 173315 309501
rect 210233 309498 210299 309501
rect 173249 309496 210299 309498
rect 173249 309440 173254 309496
rect 173310 309440 210238 309496
rect 210294 309440 210299 309496
rect 173249 309438 210299 309440
rect 173249 309435 173315 309438
rect 210233 309435 210299 309438
rect 122741 309362 122807 309365
rect 218513 309362 218579 309365
rect 122741 309360 218579 309362
rect 122741 309304 122746 309360
rect 122802 309304 218518 309360
rect 218574 309304 218579 309360
rect 122741 309302 218579 309304
rect 122741 309299 122807 309302
rect 218513 309299 218579 309302
rect 119981 309226 120047 309229
rect 237373 309226 237439 309229
rect 119981 309224 237439 309226
rect 119981 309168 119986 309224
rect 120042 309168 237378 309224
rect 237434 309168 237439 309224
rect 119981 309166 237439 309168
rect 119981 309163 120047 309166
rect 237373 309163 237439 309166
rect 244917 309226 244983 309229
rect 285857 309226 285923 309229
rect 244917 309224 285923 309226
rect 244917 309168 244922 309224
rect 244978 309168 285862 309224
rect 285918 309168 285923 309224
rect 244917 309166 285923 309168
rect 244917 309163 244983 309166
rect 285857 309163 285923 309166
rect 242801 308410 242867 308413
rect 270769 308410 270835 308413
rect 242801 308408 270835 308410
rect 242801 308352 242806 308408
rect 242862 308352 270774 308408
rect 270830 308352 270835 308408
rect 242801 308350 270835 308352
rect 242801 308347 242867 308350
rect 270769 308347 270835 308350
rect 186814 308076 186820 308140
rect 186884 308138 186890 308140
rect 233969 308138 234035 308141
rect 186884 308136 234035 308138
rect 186884 308080 233974 308136
rect 234030 308080 234035 308136
rect 186884 308078 234035 308080
rect 186884 308076 186890 308078
rect 233969 308075 234035 308078
rect 141417 308002 141483 308005
rect 213637 308002 213703 308005
rect 141417 308000 213703 308002
rect 141417 307944 141422 308000
rect 141478 307944 213642 308000
rect 213698 307944 213703 308000
rect 141417 307942 213703 307944
rect 141417 307939 141483 307942
rect 213637 307939 213703 307942
rect 17861 307866 17927 307869
rect 201585 307866 201651 307869
rect 17861 307864 201651 307866
rect 17861 307808 17866 307864
rect 17922 307808 201590 307864
rect 201646 307808 201651 307864
rect 17861 307806 201651 307808
rect 17861 307803 17927 307806
rect 201585 307803 201651 307806
rect 250805 307866 250871 307869
rect 289813 307866 289879 307869
rect 250805 307864 289879 307866
rect 250805 307808 250810 307864
rect 250866 307808 289818 307864
rect 289874 307808 289879 307864
rect 250805 307806 289879 307808
rect 250805 307803 250871 307806
rect 289813 307803 289879 307806
rect 224217 307050 224283 307053
rect 255681 307050 255747 307053
rect 224217 307048 255747 307050
rect 224217 306992 224222 307048
rect 224278 306992 255686 307048
rect 255742 306992 255747 307048
rect 224217 306990 255747 306992
rect 224217 306987 224283 306990
rect 255681 306987 255747 306990
rect 124121 306914 124187 306917
rect 238201 306914 238267 306917
rect 124121 306912 238267 306914
rect 124121 306856 124126 306912
rect 124182 306856 238206 306912
rect 238262 306856 238267 306912
rect 124121 306854 238267 306856
rect 124121 306851 124187 306854
rect 238201 306851 238267 306854
rect 197353 306778 197419 306781
rect 219617 306778 219683 306781
rect 197353 306776 219683 306778
rect 197353 306720 197358 306776
rect 197414 306720 219622 306776
rect 219678 306720 219683 306776
rect 197353 306718 219683 306720
rect 197353 306715 197419 306718
rect 219617 306715 219683 306718
rect 166206 306580 166212 306644
rect 166276 306642 166282 306644
rect 226517 306642 226583 306645
rect 166276 306640 226583 306642
rect 166276 306584 226522 306640
rect 226578 306584 226583 306640
rect 166276 306582 226583 306584
rect 166276 306580 166282 306582
rect 226517 306579 226583 306582
rect 192518 306444 192524 306508
rect 192588 306506 192594 306508
rect 197905 306506 197971 306509
rect 192588 306504 197971 306506
rect 192588 306448 197910 306504
rect 197966 306448 197971 306504
rect 192588 306446 197971 306448
rect 192588 306444 192594 306446
rect 197905 306443 197971 306446
rect 249609 306506 249675 306509
rect 275001 306506 275067 306509
rect 249609 306504 275067 306506
rect 249609 306448 249614 306504
rect 249670 306448 275006 306504
rect 275062 306448 275067 306504
rect 249609 306446 275067 306448
rect 249609 306443 249675 306446
rect 275001 306443 275067 306446
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 230473 305690 230539 305693
rect 253289 305690 253355 305693
rect 230473 305688 253355 305690
rect 230473 305632 230478 305688
rect 230534 305632 253294 305688
rect 253350 305632 253355 305688
rect 230473 305630 253355 305632
rect 230473 305627 230539 305630
rect 253289 305627 253355 305630
rect 100518 305220 100524 305284
rect 100588 305282 100594 305284
rect 131849 305282 131915 305285
rect 100588 305280 131915 305282
rect 100588 305224 131854 305280
rect 131910 305224 131915 305280
rect 100588 305222 131915 305224
rect 100588 305220 100594 305222
rect 131849 305219 131915 305222
rect 184197 305282 184263 305285
rect 197353 305282 197419 305285
rect 184197 305280 197419 305282
rect 184197 305224 184202 305280
rect 184258 305224 197358 305280
rect 197414 305224 197419 305280
rect 184197 305222 197419 305224
rect 184197 305219 184263 305222
rect 197353 305219 197419 305222
rect 130377 305146 130443 305149
rect 214833 305146 214899 305149
rect 130377 305144 214899 305146
rect 130377 305088 130382 305144
rect 130438 305088 214838 305144
rect 214894 305088 214899 305144
rect 130377 305086 214899 305088
rect 130377 305083 130443 305086
rect 214833 305083 214899 305086
rect 257286 305084 257292 305148
rect 257356 305146 257362 305148
rect 258390 305146 258396 305148
rect 257356 305086 258396 305146
rect 257356 305084 257362 305086
rect 258390 305084 258396 305086
rect 258460 305084 258466 305148
rect 126237 305010 126303 305013
rect 215385 305010 215451 305013
rect 126237 305008 215451 305010
rect 126237 304952 126242 305008
rect 126298 304952 215390 305008
rect 215446 304952 215451 305008
rect 126237 304950 215451 304952
rect 126237 304947 126303 304950
rect 215385 304947 215451 304950
rect 240593 305010 240659 305013
rect 267917 305010 267983 305013
rect 274633 305010 274699 305013
rect 240593 305008 274699 305010
rect 240593 304952 240598 305008
rect 240654 304952 267922 305008
rect 267978 304952 274638 305008
rect 274694 304952 274699 305008
rect 240593 304950 274699 304952
rect 240593 304947 240659 304950
rect 267917 304947 267983 304950
rect 274633 304947 274699 304950
rect 244774 304540 244780 304604
rect 244844 304602 244850 304604
rect 248965 304602 249031 304605
rect 244844 304600 249031 304602
rect 244844 304544 248970 304600
rect 249026 304544 249031 304600
rect 244844 304542 249031 304544
rect 244844 304540 244850 304542
rect 248965 304539 249031 304542
rect 88425 304194 88491 304197
rect 100518 304194 100524 304196
rect 88425 304192 100524 304194
rect 88425 304136 88430 304192
rect 88486 304136 100524 304192
rect 88425 304134 100524 304136
rect 88425 304131 88491 304134
rect 100518 304132 100524 304134
rect 100588 304132 100594 304196
rect 104433 304194 104499 304197
rect 122833 304194 122899 304197
rect 104433 304192 122899 304194
rect 104433 304136 104438 304192
rect 104494 304136 122838 304192
rect 122894 304136 122899 304192
rect 104433 304134 122899 304136
rect 104433 304131 104499 304134
rect 122833 304131 122899 304134
rect 228449 304194 228515 304197
rect 232773 304194 232839 304197
rect 228449 304192 232839 304194
rect 228449 304136 228454 304192
rect 228510 304136 232778 304192
rect 232834 304136 232839 304192
rect 228449 304134 232839 304136
rect 228449 304131 228515 304134
rect 232773 304131 232839 304134
rect 155217 304058 155283 304061
rect 227437 304058 227503 304061
rect 155217 304056 227503 304058
rect 155217 304000 155222 304056
rect 155278 304000 227442 304056
rect 227498 304000 227503 304056
rect 155217 303998 227503 304000
rect 155217 303995 155283 303998
rect 227437 303995 227503 303998
rect 188286 303860 188292 303924
rect 188356 303922 188362 303924
rect 212993 303922 213059 303925
rect 188356 303920 213059 303922
rect 188356 303864 212998 303920
rect 213054 303864 213059 303920
rect 188356 303862 213059 303864
rect 188356 303860 188362 303862
rect 212993 303859 213059 303862
rect 238845 303922 238911 303925
rect 583109 303922 583175 303925
rect 238845 303920 583175 303922
rect 238845 303864 238850 303920
rect 238906 303864 583114 303920
rect 583170 303864 583175 303920
rect 238845 303862 583175 303864
rect 238845 303859 238911 303862
rect 583109 303859 583175 303862
rect 189942 303724 189948 303788
rect 190012 303786 190018 303788
rect 229185 303786 229251 303789
rect 190012 303784 229251 303786
rect 190012 303728 229190 303784
rect 229246 303728 229251 303784
rect 190012 303726 229251 303728
rect 190012 303724 190018 303726
rect 229185 303723 229251 303726
rect 242433 303786 242499 303789
rect 273437 303786 273503 303789
rect 242433 303784 273503 303786
rect 242433 303728 242438 303784
rect 242494 303728 273442 303784
rect 273498 303728 273503 303784
rect 242433 303726 273503 303728
rect 242433 303723 242499 303726
rect 273437 303723 273503 303726
rect 68829 303650 68895 303653
rect 71814 303650 71820 303652
rect 68829 303648 71820 303650
rect 68829 303592 68834 303648
rect 68890 303592 71820 303648
rect 68829 303590 71820 303592
rect 68829 303587 68895 303590
rect 71814 303588 71820 303590
rect 71884 303588 71890 303652
rect 196617 303650 196683 303653
rect 197118 303650 197124 303652
rect 196617 303648 197124 303650
rect 196617 303592 196622 303648
rect 196678 303592 197124 303648
rect 196617 303590 197124 303592
rect 196617 303587 196683 303590
rect 197118 303588 197124 303590
rect 197188 303588 197194 303652
rect 231209 303650 231275 303653
rect 234613 303650 234679 303653
rect 231209 303648 234679 303650
rect 231209 303592 231214 303648
rect 231270 303592 234618 303648
rect 234674 303592 234679 303648
rect 231209 303590 234679 303592
rect 231209 303587 231275 303590
rect 234613 303587 234679 303590
rect 247718 303588 247724 303652
rect 247788 303650 247794 303652
rect 247861 303650 247927 303653
rect 247788 303648 247927 303650
rect 247788 303592 247866 303648
rect 247922 303592 247927 303648
rect 247788 303590 247927 303592
rect 247788 303588 247794 303590
rect 247861 303587 247927 303590
rect 251357 303650 251423 303653
rect 259678 303650 259684 303652
rect 251357 303648 259684 303650
rect 251357 303592 251362 303648
rect 251418 303592 259684 303648
rect 251357 303590 259684 303592
rect 251357 303587 251423 303590
rect 259678 303588 259684 303590
rect 259748 303588 259754 303652
rect 209037 302970 209103 302973
rect 225045 302970 225111 302973
rect 209037 302968 225111 302970
rect 209037 302912 209042 302968
rect 209098 302912 225050 302968
rect 225106 302912 225111 302968
rect 209037 302910 225111 302912
rect 209037 302907 209103 302910
rect 225045 302907 225111 302910
rect 197905 302834 197971 302837
rect 226793 302834 226859 302837
rect 197905 302832 226859 302834
rect 197905 302776 197910 302832
rect 197966 302776 226798 302832
rect 226854 302776 226859 302832
rect 197905 302774 226859 302776
rect 197905 302771 197971 302774
rect 226793 302771 226859 302774
rect 246297 302834 246363 302837
rect 258390 302834 258396 302836
rect 246297 302832 258396 302834
rect 246297 302776 246302 302832
rect 246358 302776 258396 302832
rect 246297 302774 258396 302776
rect 246297 302771 246363 302774
rect 258390 302772 258396 302774
rect 258460 302772 258466 302836
rect 258809 302834 258875 302837
rect 272149 302834 272215 302837
rect 258809 302832 272215 302834
rect 258809 302776 258814 302832
rect 258870 302776 272154 302832
rect 272210 302776 272215 302832
rect 258809 302774 272215 302776
rect 258809 302771 258875 302774
rect 272149 302771 272215 302774
rect 153929 302562 153995 302565
rect 201033 302562 201099 302565
rect 153929 302560 201099 302562
rect 153929 302504 153934 302560
rect 153990 302504 201038 302560
rect 201094 302504 201099 302560
rect 153929 302502 201099 302504
rect 153929 302499 153995 302502
rect 201033 302499 201099 302502
rect 180149 302426 180215 302429
rect 200389 302426 200455 302429
rect 180149 302424 200455 302426
rect 180149 302368 180154 302424
rect 180210 302368 200394 302424
rect 200450 302368 200455 302424
rect 180149 302366 200455 302368
rect 180149 302363 180215 302366
rect 200389 302363 200455 302366
rect 189901 302290 189967 302293
rect 196801 302290 196867 302293
rect 189901 302288 196867 302290
rect 189901 302232 189906 302288
rect 189962 302232 196806 302288
rect 196862 302232 196867 302288
rect 189901 302230 196867 302232
rect 189901 302227 189967 302230
rect 196801 302227 196867 302230
rect 241789 302290 241855 302293
rect 242157 302290 242223 302293
rect 276289 302290 276355 302293
rect 241789 302288 276355 302290
rect 241789 302232 241794 302288
rect 241850 302232 242162 302288
rect 242218 302232 276294 302288
rect 276350 302232 276355 302288
rect 241789 302230 276355 302232
rect 241789 302227 241855 302230
rect 242157 302227 242223 302230
rect 276289 302227 276355 302230
rect 232497 301746 232563 301749
rect 246389 301746 246455 301749
rect 247217 301746 247283 301749
rect 247861 301746 247927 301749
rect 281625 301746 281691 301749
rect 232497 301744 238770 301746
rect 232497 301688 232502 301744
rect 232558 301688 238770 301744
rect 232497 301686 238770 301688
rect 232497 301683 232563 301686
rect 160737 301610 160803 301613
rect 227713 301610 227779 301613
rect 160737 301608 227779 301610
rect 160737 301552 160742 301608
rect 160798 301552 227718 301608
rect 227774 301552 227779 301608
rect 160737 301550 227779 301552
rect 160737 301547 160803 301550
rect 227713 301547 227779 301550
rect 192334 301412 192340 301476
rect 192404 301474 192410 301476
rect 207933 301474 207999 301477
rect 192404 301472 207999 301474
rect 192404 301416 207938 301472
rect 207994 301416 207999 301472
rect 192404 301414 207999 301416
rect 238710 301474 238770 301686
rect 246389 301744 246498 301746
rect 246389 301688 246394 301744
rect 246450 301688 246498 301744
rect 246389 301683 246498 301688
rect 247217 301744 281691 301746
rect 247217 301688 247222 301744
rect 247278 301688 247866 301744
rect 247922 301688 281630 301744
rect 281686 301688 281691 301744
rect 247217 301686 281691 301688
rect 247217 301683 247283 301686
rect 247861 301683 247927 301686
rect 281625 301683 281691 301686
rect 246438 301610 246498 301683
rect 254577 301612 254643 301613
rect 254526 301610 254532 301612
rect 246438 301550 254226 301610
rect 254486 301550 254532 301610
rect 254596 301608 254643 301612
rect 254638 301552 254643 301608
rect 254025 301474 254091 301477
rect 238710 301472 254091 301474
rect 238710 301416 254030 301472
rect 254086 301416 254091 301472
rect 238710 301414 254091 301416
rect 254166 301474 254226 301550
rect 254526 301548 254532 301550
rect 254596 301548 254643 301552
rect 254577 301547 254643 301548
rect 256693 301474 256759 301477
rect 254166 301472 256759 301474
rect 254166 301416 256698 301472
rect 256754 301416 256759 301472
rect 254166 301414 256759 301416
rect 192404 301412 192410 301414
rect 207933 301411 207999 301414
rect 254025 301411 254091 301414
rect 256693 301411 256759 301414
rect 43437 301338 43503 301341
rect 198365 301338 198431 301341
rect 43437 301336 198431 301338
rect 43437 301280 43442 301336
rect 43498 301280 198370 301336
rect 198426 301280 198431 301336
rect 43437 301278 198431 301280
rect 43437 301275 43503 301278
rect 198365 301275 198431 301278
rect 193438 301140 193444 301204
rect 193508 301202 193514 301204
rect 194225 301202 194291 301205
rect 255405 301202 255471 301205
rect 193508 301200 194291 301202
rect 193508 301144 194230 301200
rect 194286 301144 194291 301200
rect 193508 301142 194291 301144
rect 253460 301200 255471 301202
rect 253460 301144 255410 301200
rect 255466 301144 255471 301200
rect 253460 301142 255471 301144
rect 193508 301140 193514 301142
rect 194225 301139 194291 301142
rect 255405 301139 255471 301142
rect 193305 301068 193371 301069
rect 193254 301066 193260 301068
rect 193214 301006 193260 301066
rect 193324 301064 193371 301068
rect 193366 301008 193371 301064
rect 193254 301004 193260 301006
rect 193324 301004 193371 301008
rect 241646 301004 241652 301068
rect 241716 301066 241722 301068
rect 242065 301066 242131 301069
rect 241716 301064 242131 301066
rect 241716 301008 242070 301064
rect 242126 301008 242131 301064
rect 241716 301006 242131 301008
rect 241716 301004 241722 301006
rect 193305 301003 193371 301004
rect 242065 301003 242131 301006
rect 191598 300868 191604 300932
rect 191668 300930 191674 300932
rect 191668 300870 193660 300930
rect 191668 300868 191674 300870
rect 194542 300868 194548 300932
rect 194612 300930 194618 300932
rect 194685 300930 194751 300933
rect 194612 300928 194751 300930
rect 194612 300872 194690 300928
rect 194746 300872 194751 300928
rect 194612 300870 194751 300872
rect 194612 300868 194618 300870
rect 194685 300867 194751 300870
rect 197302 300868 197308 300932
rect 197372 300930 197378 300932
rect 209129 300930 209195 300933
rect 197372 300928 209195 300930
rect 197372 300872 209134 300928
rect 209190 300872 209195 300928
rect 197372 300870 209195 300872
rect 197372 300868 197378 300870
rect 209129 300867 209195 300870
rect 252461 300794 252527 300797
rect 255313 300794 255379 300797
rect 252461 300792 255379 300794
rect 252461 300736 252466 300792
rect 252522 300736 255318 300792
rect 255374 300736 255379 300792
rect 252461 300734 255379 300736
rect 252461 300731 252527 300734
rect 255313 300731 255379 300734
rect 255589 300386 255655 300389
rect 253460 300384 255655 300386
rect 253460 300328 255594 300384
rect 255650 300328 255655 300384
rect 253460 300326 255655 300328
rect 255589 300323 255655 300326
rect 250294 300188 250300 300252
rect 250364 300250 250370 300252
rect 252829 300250 252895 300253
rect 250364 300248 252895 300250
rect 250364 300192 252834 300248
rect 252890 300192 252895 300248
rect 250364 300190 252895 300192
rect 250364 300188 250370 300190
rect 252829 300187 252895 300190
rect 162301 300114 162367 300117
rect 197302 300114 197308 300116
rect 162301 300112 197308 300114
rect 162301 300056 162306 300112
rect 162362 300056 197308 300112
rect 162301 300054 197308 300056
rect 162301 300051 162367 300054
rect 197302 300052 197308 300054
rect 197372 300052 197378 300116
rect 255405 299978 255471 299981
rect 253460 299976 255471 299978
rect 253460 299920 255410 299976
rect 255466 299920 255471 299976
rect 253460 299918 255471 299920
rect 255405 299915 255471 299918
rect 191741 299842 191807 299845
rect 252829 299842 252895 299845
rect 191741 299840 193660 299842
rect 191741 299784 191746 299840
rect 191802 299784 193660 299840
rect 191741 299782 193660 299784
rect 252829 299840 252938 299842
rect 252829 299784 252834 299840
rect 252890 299784 252938 299840
rect 191741 299779 191807 299782
rect 252829 299779 252938 299784
rect 191465 299706 191531 299709
rect 180750 299704 191531 299706
rect 180750 299648 191470 299704
rect 191526 299648 191531 299704
rect 180750 299646 191531 299648
rect 26141 299570 26207 299573
rect 180750 299570 180810 299646
rect 191465 299643 191531 299646
rect 252878 299706 252938 299779
rect 255773 299706 255839 299709
rect 252878 299704 255839 299706
rect 252878 299648 255778 299704
rect 255834 299648 255839 299704
rect 252878 299646 255839 299648
rect 26141 299568 180810 299570
rect 26141 299512 26146 299568
rect 26202 299512 180810 299568
rect 252878 299540 252938 299646
rect 255773 299643 255839 299646
rect 255313 299570 255379 299573
rect 280521 299570 280587 299573
rect 255313 299568 280587 299570
rect 26141 299510 180810 299512
rect 255313 299512 255318 299568
rect 255374 299512 280526 299568
rect 280582 299512 280587 299568
rect 255313 299510 280587 299512
rect 26141 299507 26207 299510
rect 255313 299507 255379 299510
rect 280521 299507 280587 299510
rect 255681 299162 255747 299165
rect 253460 299160 255747 299162
rect 253460 299104 255686 299160
rect 255742 299104 255747 299160
rect 253460 299102 255747 299104
rect 255681 299099 255747 299102
rect 138749 299026 138815 299029
rect 193489 299026 193555 299029
rect 138749 299024 193555 299026
rect 138749 298968 138754 299024
rect 138810 298968 193494 299024
rect 193550 298968 193555 299024
rect 138749 298966 193555 298968
rect 138749 298963 138815 298966
rect 193489 298963 193555 298966
rect 45461 298754 45527 298757
rect 188470 298754 188476 298756
rect 45461 298752 188476 298754
rect 45461 298696 45466 298752
rect 45522 298696 188476 298752
rect 45461 298694 188476 298696
rect 45461 298691 45527 298694
rect 188470 298692 188476 298694
rect 188540 298692 188546 298756
rect 191005 298754 191071 298757
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 191005 298752 193660 298754
rect 191005 298696 191010 298752
rect 191066 298696 193660 298752
rect 191005 298694 193660 298696
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 191005 298691 191071 298694
rect 580165 298691 580231 298694
rect 254117 298618 254183 298621
rect 255313 298618 255379 298621
rect 253460 298616 255379 298618
rect 253460 298560 254122 298616
rect 254178 298560 255318 298616
rect 255374 298560 255379 298616
rect 583520 298604 584960 298694
rect 253460 298558 255379 298560
rect 254117 298555 254183 298558
rect 255313 298555 255379 298558
rect 255405 298210 255471 298213
rect 253460 298208 255471 298210
rect 253460 298152 255410 298208
rect 255466 298152 255471 298208
rect 253460 298150 255471 298152
rect 255405 298147 255471 298150
rect 253289 298074 253355 298077
rect 253246 298072 253355 298074
rect 253246 298016 253294 298072
rect 253350 298016 253355 298072
rect 253246 298011 253355 298016
rect 259637 298076 259703 298077
rect 259637 298072 259684 298076
rect 259748 298074 259754 298076
rect 259637 298016 259642 298072
rect 259637 298012 259684 298016
rect 259748 298014 259794 298074
rect 259748 298012 259754 298014
rect 259637 298011 259703 298012
rect 253246 297772 253306 298011
rect 191741 297666 191807 297669
rect 191741 297664 193844 297666
rect 191741 297608 191746 297664
rect 191802 297636 193844 297664
rect 191802 297608 193874 297636
rect 191741 297606 193874 297608
rect 191741 297603 191807 297606
rect 81801 297530 81867 297533
rect 91502 297530 91508 297532
rect 81801 297528 91508 297530
rect 81801 297472 81806 297528
rect 81862 297472 91508 297528
rect 81801 297470 91508 297472
rect 81801 297467 81867 297470
rect 91502 297468 91508 297470
rect 91572 297530 91578 297532
rect 100017 297530 100083 297533
rect 91572 297528 100083 297530
rect 91572 297472 100022 297528
rect 100078 297472 100083 297528
rect 91572 297470 100083 297472
rect 91572 297468 91578 297470
rect 100017 297467 100083 297470
rect 129641 297530 129707 297533
rect 193814 297532 193874 297606
rect 191598 297530 191604 297532
rect 129641 297528 191604 297530
rect 129641 297472 129646 297528
rect 129702 297472 191604 297528
rect 129641 297470 191604 297472
rect 129641 297467 129707 297470
rect 191598 297468 191604 297470
rect 191668 297468 191674 297532
rect 193806 297468 193812 297532
rect 193876 297468 193882 297532
rect 4061 297394 4127 297397
rect 193254 297394 193260 297396
rect 4061 297392 193260 297394
rect 4061 297336 4066 297392
rect 4122 297336 193260 297392
rect 4061 297334 193260 297336
rect 4061 297331 4127 297334
rect 193254 297332 193260 297334
rect 193324 297332 193330 297396
rect 255405 297394 255471 297397
rect 253460 297392 255471 297394
rect 253460 297336 255410 297392
rect 255466 297336 255471 297392
rect 253460 297334 255471 297336
rect 255405 297331 255471 297334
rect 255957 297122 256023 297125
rect 255957 297120 267750 297122
rect 255957 297064 255962 297120
rect 256018 297064 267750 297120
rect 255957 297062 267750 297064
rect 255957 297059 256023 297062
rect 267690 296986 267750 297062
rect 274817 296986 274883 296989
rect 253460 296926 258090 296986
rect 267690 296984 274883 296986
rect 267690 296928 274822 296984
rect 274878 296928 274883 296984
rect 267690 296926 274883 296928
rect 258030 296850 258090 296926
rect 274817 296923 274883 296926
rect 295425 296850 295491 296853
rect 258030 296848 295491 296850
rect 258030 296792 295430 296848
rect 295486 296792 295491 296848
rect 258030 296790 295491 296792
rect 295425 296787 295491 296790
rect 191557 296578 191623 296581
rect 256601 296578 256667 296581
rect 191557 296576 193660 296578
rect 191557 296520 191562 296576
rect 191618 296520 193660 296576
rect 191557 296518 193660 296520
rect 253460 296576 256667 296578
rect 253460 296520 256606 296576
rect 256662 296520 256667 296576
rect 253460 296518 256667 296520
rect 191557 296515 191623 296518
rect 256601 296515 256667 296518
rect 255865 296170 255931 296173
rect 253460 296168 255931 296170
rect 253460 296112 255870 296168
rect 255926 296112 255931 296168
rect 253460 296110 255931 296112
rect 255865 296107 255931 296110
rect 253430 295490 253490 295596
rect 254025 295490 254091 295493
rect 253430 295488 258090 295490
rect 189809 295354 189875 295357
rect 193630 295354 193690 295460
rect 253430 295432 254030 295488
rect 254086 295432 258090 295488
rect 253430 295430 258090 295432
rect 254025 295427 254091 295430
rect 189809 295352 193690 295354
rect 189809 295296 189814 295352
rect 189870 295296 193690 295352
rect 189809 295294 193690 295296
rect 258030 295354 258090 295430
rect 291469 295354 291535 295357
rect 258030 295352 291535 295354
rect 258030 295296 291474 295352
rect 291530 295296 291535 295352
rect 258030 295294 291535 295296
rect 189809 295291 189875 295294
rect 291469 295291 291535 295294
rect 255405 295218 255471 295221
rect 253460 295216 255471 295218
rect 253460 295160 255410 295216
rect 255466 295160 255471 295216
rect 253460 295158 255471 295160
rect 255405 295155 255471 295158
rect 266629 295218 266695 295221
rect 266997 295218 267063 295221
rect 291193 295218 291259 295221
rect 266629 295216 291259 295218
rect 266629 295160 266634 295216
rect 266690 295160 267002 295216
rect 267058 295160 291198 295216
rect 291254 295160 291259 295216
rect 266629 295158 291259 295160
rect 266629 295155 266695 295158
rect 266997 295155 267063 295158
rect 291193 295155 291259 295158
rect 258533 294810 258599 294813
rect 253460 294808 258599 294810
rect 253460 294752 258538 294808
rect 258594 294752 258599 294808
rect 253460 294750 258599 294752
rect 258533 294747 258599 294750
rect 151169 294538 151235 294541
rect 192334 294538 192340 294540
rect 151169 294536 192340 294538
rect 151169 294480 151174 294536
rect 151230 294480 192340 294536
rect 151169 294478 192340 294480
rect 151169 294475 151235 294478
rect 192334 294476 192340 294478
rect 192404 294476 192410 294540
rect 191782 294340 191788 294404
rect 191852 294402 191858 294404
rect 255497 294402 255563 294405
rect 191852 294342 193660 294402
rect 253460 294400 255563 294402
rect 253460 294344 255502 294400
rect 255558 294344 255563 294400
rect 253460 294342 255563 294344
rect 191852 294340 191858 294342
rect 255497 294339 255563 294342
rect 255405 293994 255471 293997
rect 253460 293992 255471 293994
rect 253460 293936 255410 293992
rect 255466 293936 255471 293992
rect 253460 293934 255471 293936
rect 255405 293931 255471 293934
rect 255681 293586 255747 293589
rect 253460 293584 255747 293586
rect 253460 293528 255686 293584
rect 255742 293528 255747 293584
rect 253460 293526 255747 293528
rect 255681 293523 255747 293526
rect 84101 293314 84167 293317
rect 92790 293314 92796 293316
rect 84101 293312 92796 293314
rect -960 293178 480 293268
rect 84101 293256 84106 293312
rect 84162 293256 92796 293312
rect 84101 293254 92796 293256
rect 84101 293251 84167 293254
rect 92790 293252 92796 293254
rect 92860 293252 92866 293316
rect 191189 293314 191255 293317
rect 191189 293312 193660 293314
rect 191189 293256 191194 293312
rect 191250 293284 193660 293312
rect 191250 293256 193690 293284
rect 191189 293254 193690 293256
rect 191189 293251 191255 293254
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 89529 293178 89595 293181
rect 98494 293178 98500 293180
rect 89529 293176 98500 293178
rect 89529 293120 89534 293176
rect 89590 293120 98500 293176
rect 89529 293118 98500 293120
rect 89529 293115 89595 293118
rect 98494 293116 98500 293118
rect 98564 293116 98570 293180
rect 141509 293178 141575 293181
rect 193438 293178 193444 293180
rect 141509 293176 193444 293178
rect 141509 293120 141514 293176
rect 141570 293120 193444 293176
rect 141509 293118 193444 293120
rect 141509 293115 141575 293118
rect 193438 293116 193444 293118
rect 193508 293116 193514 293180
rect 77293 292770 77359 292773
rect 77293 292768 84210 292770
rect 77293 292712 77298 292768
rect 77354 292712 84210 292768
rect 77293 292710 84210 292712
rect 77293 292707 77359 292710
rect 76005 292634 76071 292637
rect 83222 292634 83228 292636
rect 76005 292632 83228 292634
rect 76005 292576 76010 292632
rect 76066 292576 83228 292632
rect 76005 292574 83228 292576
rect 76005 292571 76071 292574
rect 83222 292572 83228 292574
rect 83292 292572 83298 292636
rect 84150 292634 84210 292710
rect 193438 292708 193444 292772
rect 193508 292770 193514 292772
rect 193630 292770 193690 293254
rect 255497 293178 255563 293181
rect 253460 293176 255563 293178
rect 253460 293120 255502 293176
rect 255558 293120 255563 293176
rect 253460 293118 255563 293120
rect 255497 293115 255563 293118
rect 258533 293178 258599 293181
rect 284293 293178 284359 293181
rect 258533 293176 284359 293178
rect 258533 293120 258538 293176
rect 258594 293120 284298 293176
rect 284354 293120 284359 293176
rect 258533 293118 284359 293120
rect 258533 293115 258599 293118
rect 284293 293115 284359 293118
rect 193508 292710 193690 292770
rect 193508 292708 193514 292710
rect 119337 292634 119403 292637
rect 253841 292634 253907 292637
rect 84150 292632 119403 292634
rect 84150 292576 119342 292632
rect 119398 292576 119403 292632
rect 252908 292632 253907 292634
rect 252908 292604 253846 292632
rect 84150 292574 119403 292576
rect 119337 292571 119403 292574
rect 252878 292576 253846 292604
rect 253902 292576 253907 292632
rect 252878 292574 253907 292576
rect 252878 292501 252938 292574
rect 253841 292571 253907 292574
rect 252829 292496 252938 292501
rect 263501 292500 263567 292501
rect 263501 292498 263548 292500
rect 252829 292440 252834 292496
rect 252890 292440 252938 292496
rect 252829 292438 252938 292440
rect 263456 292496 263548 292498
rect 263456 292440 263506 292496
rect 263456 292438 263548 292440
rect 252829 292435 252895 292438
rect 263501 292436 263548 292438
rect 263612 292436 263618 292500
rect 263501 292435 263567 292436
rect 186129 292362 186195 292365
rect 191782 292362 191788 292364
rect 186129 292360 191788 292362
rect 186129 292304 186134 292360
rect 186190 292304 191788 292360
rect 186129 292302 191788 292304
rect 186129 292299 186195 292302
rect 191782 292300 191788 292302
rect 191852 292300 191858 292364
rect 191281 292226 191347 292229
rect 191281 292224 193660 292226
rect 191281 292168 191286 292224
rect 191342 292168 193660 292224
rect 191281 292166 193660 292168
rect 191281 292163 191347 292166
rect 252921 292090 252987 292093
rect 253430 292090 253490 292196
rect 256141 292090 256207 292093
rect 252921 292088 253122 292090
rect 252921 292032 252926 292088
rect 252982 292032 253122 292088
rect 252921 292030 253122 292032
rect 253430 292088 256207 292090
rect 253430 292032 256146 292088
rect 256202 292032 256207 292088
rect 253430 292030 256207 292032
rect 252921 292027 252987 292030
rect 253062 291954 253122 292030
rect 256141 292027 256207 292030
rect 253062 291894 253490 291954
rect 83089 291818 83155 291821
rect 92974 291818 92980 291820
rect 83089 291816 92980 291818
rect 83089 291760 83094 291816
rect 83150 291760 92980 291816
rect 83089 291758 92980 291760
rect 83089 291755 83155 291758
rect 92974 291756 92980 291758
rect 93044 291818 93050 291820
rect 120809 291818 120875 291821
rect 93044 291816 120875 291818
rect 93044 291760 120814 291816
rect 120870 291760 120875 291816
rect 253430 291818 253490 291894
rect 253841 291818 253907 291821
rect 253430 291816 253907 291818
rect 253430 291788 253846 291816
rect 93044 291758 120875 291760
rect 253460 291760 253846 291788
rect 253902 291760 253907 291816
rect 253460 291758 253907 291760
rect 93044 291756 93050 291758
rect 120809 291755 120875 291758
rect 253841 291755 253907 291758
rect 256417 291410 256483 291413
rect 253460 291408 256483 291410
rect 253460 291352 256422 291408
rect 256478 291352 256483 291408
rect 253460 291350 256483 291352
rect 256417 291347 256483 291350
rect 256601 291410 256667 291413
rect 280429 291410 280495 291413
rect 256601 291408 280495 291410
rect 256601 291352 256606 291408
rect 256662 291352 280434 291408
rect 280490 291352 280495 291408
rect 256601 291350 280495 291352
rect 256601 291347 256667 291350
rect 280429 291347 280495 291350
rect 116577 291274 116643 291277
rect 186129 291274 186195 291277
rect 116577 291272 186195 291274
rect 116577 291216 116582 291272
rect 116638 291216 186134 291272
rect 186190 291216 186195 291272
rect 116577 291214 186195 291216
rect 116577 291211 116643 291214
rect 186129 291211 186195 291214
rect 256141 291274 256207 291277
rect 269205 291274 269271 291277
rect 256141 291272 269271 291274
rect 256141 291216 256146 291272
rect 256202 291216 269210 291272
rect 269266 291216 269271 291272
rect 256141 291214 269271 291216
rect 256141 291211 256207 291214
rect 269205 291211 269271 291214
rect 86534 291076 86540 291140
rect 86604 291138 86610 291140
rect 91277 291138 91343 291141
rect 86604 291136 91343 291138
rect 86604 291080 91282 291136
rect 91338 291080 91343 291136
rect 86604 291078 91343 291080
rect 86604 291076 86610 291078
rect 91277 291075 91343 291078
rect 191741 291138 191807 291141
rect 191741 291136 193660 291138
rect 191741 291080 191746 291136
rect 191802 291080 193660 291136
rect 191741 291078 193660 291080
rect 191741 291075 191807 291078
rect 184054 290940 184060 291004
rect 184124 291002 184130 291004
rect 192569 291002 192635 291005
rect 256877 291002 256943 291005
rect 184124 291000 192635 291002
rect 184124 290944 192574 291000
rect 192630 290944 192635 291000
rect 184124 290942 192635 290944
rect 253460 291000 256943 291002
rect 253460 290944 256882 291000
rect 256938 290944 256943 291000
rect 253460 290942 256943 290944
rect 184124 290940 184130 290942
rect 192569 290939 192635 290942
rect 256877 290939 256943 290942
rect 61745 290458 61811 290461
rect 174537 290458 174603 290461
rect 61745 290456 174603 290458
rect 61745 290400 61750 290456
rect 61806 290400 174542 290456
rect 174598 290400 174603 290456
rect 61745 290398 174603 290400
rect 61745 290395 61811 290398
rect 174537 290395 174603 290398
rect 253430 290322 253490 290564
rect 253430 290262 263610 290322
rect 191046 289988 191052 290052
rect 191116 290050 191122 290052
rect 191649 290050 191715 290053
rect 256509 290050 256575 290053
rect 191116 290048 193660 290050
rect 191116 289992 191654 290048
rect 191710 289992 193660 290048
rect 191116 289990 193660 289992
rect 253460 290048 256575 290050
rect 253460 289992 256514 290048
rect 256570 289992 256575 290048
rect 253460 289990 256575 289992
rect 191116 289988 191122 289990
rect 191649 289987 191715 289990
rect 256509 289987 256575 289990
rect 91502 289852 91508 289916
rect 91572 289914 91578 289916
rect 96613 289914 96679 289917
rect 91572 289912 96679 289914
rect 91572 289856 96618 289912
rect 96674 289856 96679 289912
rect 91572 289854 96679 289856
rect 263550 289914 263610 290262
rect 582557 289914 582623 289917
rect 263550 289912 582623 289914
rect 263550 289856 582562 289912
rect 582618 289856 582623 289912
rect 263550 289854 582623 289856
rect 91572 289852 91578 289854
rect 96613 289851 96679 289854
rect 582557 289851 582623 289854
rect 258390 289781 258396 289832
rect 88006 289716 88012 289780
rect 88076 289778 88082 289780
rect 89713 289778 89779 289781
rect 88076 289776 89779 289778
rect 88076 289720 89718 289776
rect 89774 289720 89779 289776
rect 88076 289718 89779 289720
rect 88076 289716 88082 289718
rect 89713 289715 89779 289718
rect 258349 289776 258396 289781
rect 258349 289720 258354 289776
rect 258460 289768 258466 289832
rect 258410 289720 258458 289768
rect 258349 289718 258458 289720
rect 258349 289715 258415 289718
rect 259494 289642 259500 289644
rect 253460 289582 259500 289642
rect 259494 289580 259500 289582
rect 259564 289580 259570 289644
rect 67541 289234 67607 289237
rect 124949 289234 125015 289237
rect 67541 289232 125015 289234
rect 67541 289176 67546 289232
rect 67602 289176 124954 289232
rect 125010 289176 125015 289232
rect 67541 289174 125015 289176
rect 67541 289171 67607 289174
rect 124949 289171 125015 289174
rect 63125 289098 63191 289101
rect 177246 289098 177252 289100
rect 63125 289096 177252 289098
rect 63125 289040 63130 289096
rect 63186 289040 177252 289096
rect 63125 289038 177252 289040
rect 63125 289035 63191 289038
rect 177246 289036 177252 289038
rect 177316 289036 177322 289100
rect 253430 289098 253490 289204
rect 253430 289038 263610 289098
rect 191649 288962 191715 288965
rect 192702 288962 192708 288964
rect 191649 288960 192708 288962
rect 191649 288904 191654 288960
rect 191710 288904 192708 288960
rect 191649 288902 192708 288904
rect 191649 288899 191715 288902
rect 192702 288900 192708 288902
rect 192772 288962 192778 288964
rect 192772 288902 193660 288962
rect 192772 288900 192778 288902
rect 255957 288826 256023 288829
rect 253460 288824 256023 288826
rect 253460 288768 255962 288824
rect 256018 288768 256023 288824
rect 253460 288766 256023 288768
rect 255957 288763 256023 288766
rect 263550 288690 263610 289038
rect 273529 288690 273595 288693
rect 263550 288688 273595 288690
rect 263550 288632 273534 288688
rect 273590 288632 273595 288688
rect 263550 288630 273595 288632
rect 273529 288627 273595 288630
rect 90950 288492 90956 288556
rect 91020 288554 91026 288556
rect 95233 288554 95299 288557
rect 91020 288552 95299 288554
rect 91020 288496 95238 288552
rect 95294 288496 95299 288552
rect 91020 288494 95299 288496
rect 91020 288492 91026 288494
rect 95233 288491 95299 288494
rect 177798 288492 177804 288556
rect 177868 288554 177874 288556
rect 180793 288554 180859 288557
rect 177868 288552 180859 288554
rect 177868 288496 180798 288552
rect 180854 288496 180859 288552
rect 177868 288494 180859 288496
rect 177868 288492 177874 288494
rect 180793 288491 180859 288494
rect 11697 288418 11763 288421
rect 70894 288418 70900 288420
rect 11697 288416 70900 288418
rect 11697 288360 11702 288416
rect 11758 288360 70900 288416
rect 11697 288358 70900 288360
rect 11697 288355 11763 288358
rect 70894 288356 70900 288358
rect 70964 288356 70970 288420
rect 191833 288418 191899 288421
rect 192518 288418 192524 288420
rect 191833 288416 192524 288418
rect 191833 288360 191838 288416
rect 191894 288360 192524 288416
rect 191833 288358 192524 288360
rect 191833 288355 191899 288358
rect 192518 288356 192524 288358
rect 192588 288356 192594 288420
rect 256601 288418 256667 288421
rect 253460 288416 256667 288418
rect 253460 288360 256606 288416
rect 256662 288360 256667 288416
rect 253460 288358 256667 288360
rect 256601 288355 256667 288358
rect 269113 288418 269179 288421
rect 272149 288418 272215 288421
rect 269113 288416 272215 288418
rect 269113 288360 269118 288416
rect 269174 288360 272154 288416
rect 272210 288360 272215 288416
rect 269113 288358 272215 288360
rect 269113 288355 269179 288358
rect 272149 288355 272215 288358
rect 255865 288010 255931 288013
rect 253460 288008 255931 288010
rect 253460 287952 255870 288008
rect 255926 287952 255931 288008
rect 253460 287950 255931 287952
rect 255865 287947 255931 287950
rect 191741 287874 191807 287877
rect 192334 287874 192340 287876
rect 191741 287872 192340 287874
rect 191741 287816 191746 287872
rect 191802 287816 192340 287872
rect 191741 287814 192340 287816
rect 191741 287811 191807 287814
rect 192334 287812 192340 287814
rect 192404 287874 192410 287876
rect 192404 287814 193660 287874
rect 192404 287812 192410 287814
rect 66662 287676 66668 287740
rect 66732 287738 66738 287740
rect 97257 287738 97323 287741
rect 66732 287736 97323 287738
rect 66732 287680 97262 287736
rect 97318 287680 97323 287736
rect 66732 287678 97323 287680
rect 66732 287676 66738 287678
rect 97257 287675 97323 287678
rect 65977 287602 66043 287605
rect 66161 287602 66227 287605
rect 255773 287602 255839 287605
rect 65977 287600 66227 287602
rect 65977 287544 65982 287600
rect 66038 287544 66166 287600
rect 66222 287544 66227 287600
rect 65977 287542 66227 287544
rect 253460 287600 255839 287602
rect 253460 287544 255778 287600
rect 255834 287544 255839 287600
rect 253460 287542 255839 287544
rect 65977 287539 66043 287542
rect 66161 287539 66227 287542
rect 255773 287539 255839 287542
rect 256601 287330 256667 287333
rect 269113 287330 269179 287333
rect 256601 287328 269179 287330
rect 256601 287272 256606 287328
rect 256662 287272 269118 287328
rect 269174 287272 269179 287328
rect 256601 287270 269179 287272
rect 256601 287267 256667 287270
rect 269113 287267 269179 287270
rect 66161 287194 66227 287197
rect 120717 287194 120783 287197
rect 66161 287192 120783 287194
rect 66161 287136 66166 287192
rect 66222 287136 120722 287192
rect 120778 287136 120783 287192
rect 66161 287134 120783 287136
rect 66161 287131 66227 287134
rect 120717 287131 120783 287134
rect 253430 286922 253490 287028
rect 256509 286922 256575 286925
rect 263685 286922 263751 286925
rect 253430 286920 263751 286922
rect 253430 286864 256514 286920
rect 256570 286864 263690 286920
rect 263746 286864 263751 286920
rect 253430 286862 263751 286864
rect 256509 286859 256575 286862
rect 263685 286859 263751 286862
rect 191097 286786 191163 286789
rect 191097 286784 193660 286786
rect 191097 286728 191102 286784
rect 191158 286728 193660 286784
rect 191097 286726 193660 286728
rect 191097 286723 191163 286726
rect 256601 286650 256667 286653
rect 253460 286648 256667 286650
rect 253460 286592 256606 286648
rect 256662 286592 256667 286648
rect 253460 286590 256667 286592
rect 256601 286587 256667 286590
rect 97257 286378 97323 286381
rect 188337 286378 188403 286381
rect 97257 286376 188403 286378
rect 97257 286320 97262 286376
rect 97318 286320 188342 286376
rect 188398 286320 188403 286376
rect 97257 286318 188403 286320
rect 97257 286315 97323 286318
rect 188337 286315 188403 286318
rect 65977 286242 66043 286245
rect 73797 286242 73863 286245
rect 256417 286242 256483 286245
rect 65977 286240 73863 286242
rect 65977 286184 65982 286240
rect 66038 286184 73802 286240
rect 73858 286184 73863 286240
rect 65977 286182 73863 286184
rect 253460 286240 256483 286242
rect 253460 286184 256422 286240
rect 256478 286184 256483 286240
rect 253460 286182 256483 286184
rect 65977 286179 66043 286182
rect 73797 286179 73863 286182
rect 256417 286179 256483 286182
rect 72918 286044 72924 286108
rect 72988 286106 72994 286108
rect 81525 286106 81591 286109
rect 82077 286106 82143 286109
rect 72988 286104 82143 286106
rect 72988 286048 81530 286104
rect 81586 286048 82082 286104
rect 82138 286048 82143 286104
rect 72988 286046 82143 286048
rect 72988 286044 72994 286046
rect 81525 286043 81591 286046
rect 82077 286043 82143 286046
rect 83181 286106 83247 286109
rect 84101 286106 84167 286109
rect 83181 286104 84167 286106
rect 83181 286048 83186 286104
rect 83242 286048 84106 286104
rect 84162 286048 84167 286104
rect 83181 286046 84167 286048
rect 83181 286043 83247 286046
rect 84101 286043 84167 286046
rect 90265 286106 90331 286109
rect 91001 286106 91067 286109
rect 90265 286104 91067 286106
rect 90265 286048 90270 286104
rect 90326 286048 91006 286104
rect 91062 286048 91067 286104
rect 90265 286046 91067 286048
rect 90265 286043 90331 286046
rect 91001 286043 91067 286046
rect 52177 285970 52243 285973
rect 74901 285970 74967 285973
rect 75177 285970 75243 285973
rect 52177 285968 75243 285970
rect 52177 285912 52182 285968
rect 52238 285912 74906 285968
rect 74962 285912 75182 285968
rect 75238 285912 75243 285968
rect 52177 285910 75243 285912
rect 52177 285907 52243 285910
rect 74901 285907 74967 285910
rect 75177 285907 75243 285910
rect 80973 285970 81039 285973
rect 95182 285970 95188 285972
rect 80973 285968 95188 285970
rect 80973 285912 80978 285968
rect 81034 285912 95188 285968
rect 80973 285910 95188 285912
rect 80973 285907 81039 285910
rect 95182 285908 95188 285910
rect 95252 285908 95258 285972
rect 266353 285970 266419 285973
rect 253430 285968 267750 285970
rect 253430 285912 266358 285968
rect 266414 285912 267750 285968
rect 253430 285910 267750 285912
rect 70853 285836 70919 285837
rect 70853 285834 70900 285836
rect 70808 285832 70900 285834
rect 70808 285776 70858 285832
rect 70808 285774 70900 285776
rect 70853 285772 70900 285774
rect 70964 285772 70970 285836
rect 253430 285804 253490 285910
rect 266353 285907 266419 285910
rect 70853 285771 70919 285772
rect 70393 285698 70459 285701
rect 70894 285698 70900 285700
rect 70393 285696 70900 285698
rect 70393 285640 70398 285696
rect 70454 285640 70900 285696
rect 70393 285638 70900 285640
rect 70393 285635 70459 285638
rect 70894 285636 70900 285638
rect 70964 285636 70970 285700
rect 73705 285698 73771 285701
rect 79317 285698 79383 285701
rect 73705 285696 79383 285698
rect 73705 285640 73710 285696
rect 73766 285640 79322 285696
rect 79378 285640 79383 285696
rect 73705 285638 79383 285640
rect 73705 285635 73771 285638
rect 79317 285635 79383 285638
rect 90817 285698 90883 285701
rect 93853 285698 93919 285701
rect 90817 285696 93919 285698
rect 90817 285640 90822 285696
rect 90878 285640 93858 285696
rect 93914 285640 93919 285696
rect 90817 285638 93919 285640
rect 90817 285635 90883 285638
rect 93853 285635 93919 285638
rect 96429 285698 96495 285701
rect 149053 285698 149119 285701
rect 96429 285696 149119 285698
rect 96429 285640 96434 285696
rect 96490 285640 149058 285696
rect 149114 285640 149119 285696
rect 96429 285638 149119 285640
rect 96429 285635 96495 285638
rect 149053 285635 149119 285638
rect 192569 285698 192635 285701
rect 193121 285698 193187 285701
rect 267690 285698 267750 285910
rect 268009 285698 268075 285701
rect 192569 285696 193660 285698
rect 192569 285640 192574 285696
rect 192630 285640 193126 285696
rect 193182 285640 193660 285696
rect 192569 285638 193660 285640
rect 267690 285696 268075 285698
rect 267690 285640 268014 285696
rect 268070 285640 268075 285696
rect 267690 285638 268075 285640
rect 192569 285635 192635 285638
rect 193121 285635 193187 285638
rect 268009 285635 268075 285638
rect 256601 285426 256667 285429
rect 253460 285424 256667 285426
rect 253460 285368 256606 285424
rect 256662 285368 256667 285424
rect 253460 285366 256667 285368
rect 256601 285363 256667 285366
rect 583520 285276 584960 285516
rect 93853 285018 93919 285021
rect 113909 285018 113975 285021
rect 93853 285016 113975 285018
rect 93853 284960 93858 285016
rect 93914 284960 113914 285016
rect 113970 284960 113975 285016
rect 258349 285020 258415 285021
rect 258349 285016 258396 285020
rect 258460 285018 258466 285020
rect 93853 284958 113975 284960
rect 93853 284955 93919 284958
rect 113909 284955 113975 284958
rect 70301 284882 70367 284885
rect 76414 284882 76420 284884
rect 70301 284880 76420 284882
rect 70301 284824 70306 284880
rect 70362 284824 76420 284880
rect 70301 284822 76420 284824
rect 70301 284819 70367 284822
rect 76414 284820 76420 284822
rect 76484 284882 76490 284884
rect 98729 284882 98795 284885
rect 76484 284880 98795 284882
rect 76484 284824 98734 284880
rect 98790 284824 98795 284880
rect 76484 284822 98795 284824
rect 253430 284882 253490 284988
rect 258349 284960 258354 285016
rect 258349 284956 258396 284960
rect 258460 284958 258506 285018
rect 258460 284956 258466 284958
rect 258349 284955 258415 284956
rect 260833 284882 260899 284885
rect 273529 284882 273595 284885
rect 253430 284880 273595 284882
rect 253430 284824 260838 284880
rect 260894 284824 273534 284880
rect 273590 284824 273595 284880
rect 253430 284822 273595 284824
rect 76484 284820 76490 284822
rect 98729 284819 98795 284822
rect 260833 284819 260899 284822
rect 273529 284819 273595 284822
rect 191741 284610 191807 284613
rect 191741 284608 193660 284610
rect 191741 284552 191746 284608
rect 191802 284552 193660 284608
rect 191741 284550 193660 284552
rect 191741 284547 191807 284550
rect 253430 284474 253490 284580
rect 266353 284474 266419 284477
rect 266629 284474 266695 284477
rect 253430 284472 266695 284474
rect 253430 284416 266358 284472
rect 266414 284416 266634 284472
rect 266690 284416 266695 284472
rect 253430 284414 266695 284416
rect 266353 284411 266419 284414
rect 266629 284411 266695 284414
rect 50981 284338 51047 284341
rect 69197 284338 69263 284341
rect 50981 284336 69263 284338
rect 50981 284280 50986 284336
rect 51042 284280 69202 284336
rect 69258 284280 69263 284336
rect 50981 284278 69263 284280
rect 50981 284275 51047 284278
rect 69197 284275 69263 284278
rect 256601 284066 256667 284069
rect 253460 284064 256667 284066
rect 253460 284008 256606 284064
rect 256662 284008 256667 284064
rect 253460 284006 256667 284008
rect 256601 284003 256667 284006
rect 86677 283796 86743 283797
rect 86677 283792 86724 283796
rect 86788 283794 86794 283796
rect 86677 283736 86682 283792
rect 86677 283732 86724 283736
rect 86788 283734 86834 283794
rect 86788 283732 86794 283734
rect 86677 283731 86743 283732
rect 71630 283596 71636 283660
rect 71700 283658 71706 283660
rect 71957 283658 72023 283661
rect 258165 283658 258231 283661
rect 71700 283656 72023 283658
rect 71700 283600 71962 283656
rect 72018 283600 72023 283656
rect 71700 283598 72023 283600
rect 253460 283656 258231 283658
rect 253460 283600 258170 283656
rect 258226 283600 258231 283656
rect 253460 283598 258231 283600
rect 71700 283596 71706 283598
rect 71957 283595 72023 283598
rect 258165 283595 258231 283598
rect 68686 283460 68692 283524
rect 68756 283522 68762 283524
rect 69289 283522 69355 283525
rect 89529 283524 89595 283525
rect 90081 283524 90147 283525
rect 89478 283522 89484 283524
rect 68756 283520 69355 283522
rect 68756 283464 69294 283520
rect 69350 283464 69355 283520
rect 68756 283462 69355 283464
rect 89438 283462 89484 283522
rect 89548 283520 89595 283524
rect 90030 283522 90036 283524
rect 89590 283464 89595 283520
rect 68756 283460 68762 283462
rect 69289 283459 69355 283462
rect 89478 283460 89484 283462
rect 89548 283460 89595 283464
rect 89990 283462 90036 283522
rect 90100 283520 90147 283524
rect 90142 283464 90147 283520
rect 90030 283460 90036 283462
rect 90100 283460 90147 283464
rect 93894 283460 93900 283524
rect 93964 283522 93970 283524
rect 94037 283522 94103 283525
rect 93964 283520 94103 283522
rect 93964 283464 94042 283520
rect 94098 283464 94103 283520
rect 93964 283462 94103 283464
rect 93964 283460 93970 283462
rect 89529 283459 89595 283460
rect 90081 283459 90147 283460
rect 94037 283459 94103 283462
rect 191741 283522 191807 283525
rect 259269 283522 259335 283525
rect 269389 283522 269455 283525
rect 191741 283520 194212 283522
rect 191741 283464 191746 283520
rect 191802 283492 194212 283520
rect 259269 283520 269455 283522
rect 191802 283464 194242 283492
rect 191741 283462 194242 283464
rect 191741 283459 191807 283462
rect 60549 283386 60615 283389
rect 100845 283386 100911 283389
rect 194182 283388 194242 283462
rect 259269 283464 259274 283520
rect 259330 283464 269394 283520
rect 269450 283464 269455 283520
rect 259269 283462 269455 283464
rect 259269 283459 259335 283462
rect 269389 283459 269455 283462
rect 60549 283384 100911 283386
rect 60549 283328 60554 283384
rect 60610 283328 100850 283384
rect 100906 283328 100911 283384
rect 60549 283326 100911 283328
rect 60549 283323 60615 283326
rect 100845 283323 100911 283326
rect 194174 283324 194180 283388
rect 194244 283324 194250 283388
rect 69105 283250 69171 283253
rect 83457 283252 83523 283253
rect 69238 283250 69244 283252
rect 69105 283248 69244 283250
rect 69105 283192 69110 283248
rect 69166 283192 69244 283248
rect 69105 283190 69244 283192
rect 69105 283187 69171 283190
rect 69238 283188 69244 283190
rect 69308 283188 69314 283252
rect 83406 283250 83412 283252
rect 83366 283190 83412 283250
rect 83476 283248 83523 283252
rect 83518 283192 83523 283248
rect 83406 283188 83412 283190
rect 83476 283188 83523 283192
rect 84694 283188 84700 283252
rect 84764 283250 84770 283252
rect 88149 283250 88215 283253
rect 84764 283248 88215 283250
rect 84764 283192 88154 283248
rect 88210 283192 88215 283248
rect 84764 283190 88215 283192
rect 84764 283188 84770 283190
rect 83457 283187 83523 283188
rect 88149 283187 88215 283190
rect 92381 283250 92447 283253
rect 256325 283250 256391 283253
rect 92381 283248 180810 283250
rect 92381 283192 92386 283248
rect 92442 283192 180810 283248
rect 92381 283190 180810 283192
rect 253460 283248 256391 283250
rect 253460 283192 256330 283248
rect 256386 283192 256391 283248
rect 253460 283190 256391 283192
rect 92381 283187 92447 283190
rect 71630 283052 71636 283116
rect 71700 283114 71706 283116
rect 72693 283114 72759 283117
rect 71700 283112 72759 283114
rect 71700 283056 72698 283112
rect 72754 283056 72759 283112
rect 71700 283054 72759 283056
rect 71700 283052 71706 283054
rect 72693 283051 72759 283054
rect 73286 283052 73292 283116
rect 73356 283114 73362 283116
rect 73705 283114 73771 283117
rect 73356 283112 73771 283114
rect 73356 283056 73710 283112
rect 73766 283056 73771 283112
rect 73356 283054 73771 283056
rect 73356 283052 73362 283054
rect 73705 283051 73771 283054
rect 66253 282978 66319 282981
rect 68001 282978 68067 282981
rect 72417 282980 72483 282981
rect 73521 282980 73587 282981
rect 66253 282976 68908 282978
rect 66253 282920 66258 282976
rect 66314 282920 68006 282976
rect 68062 282920 68908 282976
rect 66253 282918 68908 282920
rect 66253 282915 66319 282918
rect 68001 282915 68067 282918
rect 72366 282916 72372 282980
rect 72436 282978 72483 282980
rect 72436 282976 72528 282978
rect 72478 282920 72528 282976
rect 72436 282918 72528 282920
rect 72436 282916 72483 282918
rect 73470 282916 73476 282980
rect 73540 282978 73587 282980
rect 97901 282978 97967 282981
rect 100109 282978 100175 282981
rect 73540 282976 73632 282978
rect 73582 282920 73632 282976
rect 73540 282918 73632 282920
rect 97901 282976 100175 282978
rect 97901 282920 97906 282976
rect 97962 282920 100114 282976
rect 100170 282920 100175 282976
rect 97901 282918 100175 282920
rect 180750 282978 180810 283190
rect 256325 283187 256391 283190
rect 186405 282978 186471 282981
rect 187049 282978 187115 282981
rect 263501 282980 263567 282981
rect 263501 282978 263548 282980
rect 180750 282976 187115 282978
rect 180750 282920 186410 282976
rect 186466 282920 187054 282976
rect 187110 282920 187115 282976
rect 180750 282918 187115 282920
rect 263456 282976 263548 282978
rect 263456 282920 263506 282976
rect 263456 282918 263548 282920
rect 73540 282916 73587 282918
rect 72417 282915 72483 282916
rect 73521 282915 73587 282916
rect 97901 282915 97967 282918
rect 100109 282915 100175 282918
rect 186405 282915 186471 282918
rect 187049 282915 187115 282918
rect 263501 282916 263548 282918
rect 263612 282916 263618 282980
rect 263501 282915 263567 282916
rect 67633 282842 67699 282845
rect 69054 282842 69060 282844
rect 67633 282840 69060 282842
rect 67633 282784 67638 282840
rect 67694 282784 69060 282840
rect 67633 282782 69060 282784
rect 67633 282779 67699 282782
rect 69054 282780 69060 282782
rect 69124 282780 69130 282844
rect 100753 282706 100819 282709
rect 98716 282704 100819 282706
rect 98716 282648 100758 282704
rect 100814 282648 100819 282704
rect 98716 282646 100819 282648
rect 253430 282706 253490 282812
rect 253430 282646 258090 282706
rect 100753 282643 100819 282646
rect 190453 282434 190519 282437
rect 255497 282434 255563 282437
rect 190453 282432 193660 282434
rect 190453 282376 190458 282432
rect 190514 282376 193660 282432
rect 190453 282374 193660 282376
rect 253460 282432 255563 282434
rect 253460 282376 255502 282432
rect 255558 282376 255563 282432
rect 253460 282374 255563 282376
rect 190453 282371 190519 282374
rect 255497 282371 255563 282374
rect 67541 282162 67607 282165
rect 142889 282162 142955 282165
rect 152733 282162 152799 282165
rect 67541 282160 68908 282162
rect 67541 282104 67546 282160
rect 67602 282104 68908 282160
rect 67541 282102 68908 282104
rect 142889 282160 152799 282162
rect 142889 282104 142894 282160
rect 142950 282104 152738 282160
rect 152794 282104 152799 282160
rect 142889 282102 152799 282104
rect 67541 282099 67607 282102
rect 142889 282099 142955 282102
rect 152733 282099 152799 282102
rect 256601 282026 256667 282029
rect 253460 282024 256667 282026
rect 253460 281968 256606 282024
rect 256662 281968 256667 282024
rect 253460 281966 256667 281968
rect 256601 281963 256667 281966
rect 98686 281618 98746 281860
rect 258030 281754 258090 282646
rect 276197 281754 276263 281757
rect 258030 281752 276263 281754
rect 258030 281696 276202 281752
rect 276258 281696 276263 281752
rect 258030 281694 276263 281696
rect 276197 281691 276263 281694
rect 133321 281618 133387 281621
rect 98686 281616 133387 281618
rect 98686 281560 133326 281616
rect 133382 281560 133387 281616
rect 98686 281558 133387 281560
rect 133321 281555 133387 281558
rect 103421 281482 103487 281485
rect 116485 281482 116551 281485
rect 259269 281482 259335 281485
rect 103421 281480 116551 281482
rect 103421 281424 103426 281480
rect 103482 281424 116490 281480
rect 116546 281424 116551 281480
rect 103421 281422 116551 281424
rect 253460 281480 259335 281482
rect 253460 281424 259274 281480
rect 259330 281424 259335 281480
rect 253460 281422 259335 281424
rect 103421 281419 103487 281422
rect 116485 281419 116551 281422
rect 259269 281419 259335 281422
rect 272149 281482 272215 281485
rect 274725 281482 274791 281485
rect 272149 281480 274791 281482
rect 272149 281424 272154 281480
rect 272210 281424 274730 281480
rect 274786 281424 274791 281480
rect 272149 281422 274791 281424
rect 272149 281419 272215 281422
rect 274725 281419 274791 281422
rect 190545 281346 190611 281349
rect 191741 281346 191807 281349
rect 190545 281344 193660 281346
rect 68878 281213 68938 281316
rect 190545 281288 190550 281344
rect 190606 281288 191746 281344
rect 191802 281288 193660 281344
rect 190545 281286 193660 281288
rect 190545 281283 190611 281286
rect 191741 281283 191807 281286
rect 68829 281208 68938 281213
rect 68829 281152 68834 281208
rect 68890 281152 68938 281208
rect 68829 281150 68938 281152
rect 68829 281147 68895 281150
rect 101673 281074 101739 281077
rect 255497 281074 255563 281077
rect 98716 281072 101739 281074
rect 98716 281016 101678 281072
rect 101734 281016 101739 281072
rect 98716 281014 101739 281016
rect 253460 281072 255563 281074
rect 253460 281016 255502 281072
rect 255558 281016 255563 281072
rect 253460 281014 255563 281016
rect 101673 281011 101739 281014
rect 255497 281011 255563 281014
rect 169661 280938 169727 280941
rect 177297 280938 177363 280941
rect 169661 280936 177363 280938
rect 169661 280880 169666 280936
rect 169722 280880 177302 280936
rect 177358 280880 177363 280936
rect 169661 280878 177363 280880
rect 169661 280875 169727 280878
rect 177297 280875 177363 280878
rect 175273 280802 175339 280805
rect 189809 280802 189875 280805
rect 175273 280800 189875 280802
rect 175273 280744 175278 280800
rect 175334 280744 189814 280800
rect 189870 280744 189875 280800
rect 175273 280742 189875 280744
rect 175273 280739 175339 280742
rect 189809 280739 189875 280742
rect 67950 280468 67956 280532
rect 68020 280530 68026 280532
rect 253430 280530 253490 280636
rect 68020 280470 68908 280530
rect 253430 280470 258090 280530
rect 68020 280468 68026 280470
rect 258030 280394 258090 280470
rect 272149 280394 272215 280397
rect 258030 280392 272215 280394
rect 258030 280336 272154 280392
rect 272210 280336 272215 280392
rect 258030 280334 272215 280336
rect 272149 280331 272215 280334
rect 99373 280258 99439 280261
rect 103421 280258 103487 280261
rect 98716 280256 103487 280258
rect -960 279972 480 280212
rect 98716 280200 99378 280256
rect 99434 280200 103426 280256
rect 103482 280200 103487 280256
rect 98716 280198 103487 280200
rect 99373 280195 99439 280198
rect 103421 280195 103487 280198
rect 191465 280258 191531 280261
rect 255313 280258 255379 280261
rect 191465 280256 193660 280258
rect 191465 280200 191470 280256
rect 191526 280200 193660 280256
rect 191465 280198 193660 280200
rect 253460 280256 255379 280258
rect 253460 280200 255318 280256
rect 255374 280200 255379 280256
rect 253460 280198 255379 280200
rect 191465 280195 191531 280198
rect 255313 280195 255379 280198
rect 162209 280122 162275 280125
rect 166206 280122 166212 280124
rect 162209 280120 166212 280122
rect 162209 280064 162214 280120
rect 162270 280064 166212 280120
rect 162209 280062 166212 280064
rect 162209 280059 162275 280062
rect 166206 280060 166212 280062
rect 166276 280060 166282 280124
rect 255681 279850 255747 279853
rect 253460 279848 255747 279850
rect 253460 279792 255686 279848
rect 255742 279792 255747 279848
rect 253460 279790 255747 279792
rect 255681 279787 255747 279790
rect 67357 279714 67423 279717
rect 67357 279712 68908 279714
rect 67357 279656 67362 279712
rect 67418 279656 68908 279712
rect 67357 279654 68908 279656
rect 67357 279651 67423 279654
rect 255313 279442 255379 279445
rect 253460 279440 255379 279442
rect 66805 278898 66871 278901
rect 98686 278898 98746 279412
rect 253460 279384 255318 279440
rect 255374 279384 255379 279440
rect 253460 279382 255379 279384
rect 255313 279379 255379 279382
rect 190453 279170 190519 279173
rect 190453 279168 193660 279170
rect 190453 279112 190458 279168
rect 190514 279112 193660 279168
rect 190453 279110 193660 279112
rect 190453 279107 190519 279110
rect 255497 279034 255563 279037
rect 253460 279032 255563 279034
rect 253460 278976 255502 279032
rect 255558 278976 255563 279032
rect 253460 278974 255563 278976
rect 255497 278971 255563 278974
rect 162393 278898 162459 278901
rect 66805 278896 68908 278898
rect 66805 278840 66810 278896
rect 66866 278840 68908 278896
rect 66805 278838 68908 278840
rect 98686 278896 162459 278898
rect 98686 278840 162398 278896
rect 162454 278840 162459 278896
rect 98686 278838 162459 278840
rect 66805 278835 66871 278838
rect 162393 278835 162459 278838
rect 100753 278626 100819 278629
rect 98716 278624 100819 278626
rect 98716 278568 100758 278624
rect 100814 278568 100819 278624
rect 98716 278566 100819 278568
rect 100753 278563 100819 278566
rect 255497 278490 255563 278493
rect 253460 278488 255563 278490
rect 253460 278432 255502 278488
rect 255558 278432 255563 278488
rect 253460 278430 255563 278432
rect 255497 278427 255563 278430
rect 111742 278218 111748 278220
rect 103470 278158 111748 278218
rect 66805 278082 66871 278085
rect 103470 278082 103530 278158
rect 111742 278156 111748 278158
rect 111812 278218 111818 278220
rect 112805 278218 112871 278221
rect 111812 278216 112871 278218
rect 111812 278160 112810 278216
rect 112866 278160 112871 278216
rect 111812 278158 112871 278160
rect 111812 278156 111818 278158
rect 112805 278155 112871 278158
rect 255681 278218 255747 278221
rect 255681 278216 258090 278218
rect 255681 278160 255686 278216
rect 255742 278160 258090 278216
rect 255681 278158 258090 278160
rect 255681 278155 255747 278158
rect 66805 278080 68908 278082
rect 66805 278024 66810 278080
rect 66866 278024 68908 278080
rect 66805 278022 68908 278024
rect 98686 278022 103530 278082
rect 190453 278082 190519 278085
rect 257286 278082 257292 278084
rect 190453 278080 193660 278082
rect 190453 278024 190458 278080
rect 190514 278024 193660 278080
rect 190453 278022 193660 278024
rect 253460 278022 257292 278082
rect 66805 278019 66871 278022
rect 98686 277810 98746 278022
rect 190453 278019 190519 278022
rect 257286 278020 257292 278022
rect 257356 278020 257362 278084
rect 258030 278082 258090 278158
rect 259453 278082 259519 278085
rect 269297 278082 269363 278085
rect 258030 278080 269363 278082
rect 258030 278024 259458 278080
rect 259514 278024 269302 278080
rect 269358 278024 269363 278080
rect 258030 278022 269363 278024
rect 259453 278019 259519 278022
rect 269297 278019 269363 278022
rect 98532 277780 98746 277810
rect 98502 277750 98716 277780
rect 98502 277540 98562 277750
rect 98494 277476 98500 277540
rect 98564 277476 98570 277540
rect 253430 277538 253490 277644
rect 262213 277538 262279 277541
rect 253430 277536 262279 277538
rect 253430 277480 262218 277536
rect 262274 277480 262279 277536
rect 253430 277478 262279 277480
rect 262213 277475 262279 277478
rect 67633 277266 67699 277269
rect 255497 277266 255563 277269
rect 67633 277264 68908 277266
rect 67633 277208 67638 277264
rect 67694 277208 68908 277264
rect 67633 277206 68908 277208
rect 253460 277264 255563 277266
rect 253460 277208 255502 277264
rect 255558 277208 255563 277264
rect 253460 277206 255563 277208
rect 67633 277203 67699 277206
rect 255497 277203 255563 277206
rect 101254 276994 101260 276996
rect 98716 276934 101260 276994
rect 101254 276932 101260 276934
rect 101324 276932 101330 276996
rect 190453 276994 190519 276997
rect 190453 276992 193660 276994
rect 190453 276936 190458 276992
rect 190514 276936 193660 276992
rect 190453 276934 193660 276936
rect 190453 276931 190519 276934
rect 259545 276858 259611 276861
rect 253460 276856 259611 276858
rect 253460 276800 259550 276856
rect 259606 276800 259611 276856
rect 253460 276798 259611 276800
rect 259545 276795 259611 276798
rect 66805 276450 66871 276453
rect 255313 276450 255379 276453
rect 66805 276448 68908 276450
rect 66805 276392 66810 276448
rect 66866 276392 68908 276448
rect 66805 276390 68908 276392
rect 253460 276448 255379 276450
rect 253460 276392 255318 276448
rect 255374 276392 255379 276448
rect 253460 276390 255379 276392
rect 66805 276387 66871 276390
rect 255313 276387 255379 276390
rect 100753 276178 100819 276181
rect 98716 276176 100819 276178
rect 98716 276120 100758 276176
rect 100814 276120 100819 276176
rect 98716 276118 100819 276120
rect 100753 276115 100819 276118
rect 68553 276042 68619 276045
rect 69238 276042 69244 276044
rect 68553 276040 69244 276042
rect 68553 275984 68558 276040
rect 68614 275984 69244 276040
rect 68553 275982 69244 275984
rect 68553 275979 68619 275982
rect 69238 275980 69244 275982
rect 69308 275980 69314 276044
rect 271873 276042 271939 276045
rect 273253 276042 273319 276045
rect 253460 276040 273319 276042
rect 253460 275984 271878 276040
rect 271934 275984 273258 276040
rect 273314 275984 273319 276040
rect 253460 275982 273319 275984
rect 271873 275979 271939 275982
rect 273253 275979 273319 275982
rect 190453 275906 190519 275909
rect 190453 275904 193660 275906
rect 190453 275848 190458 275904
rect 190514 275848 193660 275904
rect 190453 275846 193660 275848
rect 190453 275843 190519 275846
rect 66805 275634 66871 275637
rect 66805 275632 68908 275634
rect 66805 275576 66810 275632
rect 66866 275576 68908 275632
rect 66805 275574 68908 275576
rect 66805 275571 66871 275574
rect 255497 275498 255563 275501
rect 253460 275496 255563 275498
rect 253460 275440 255502 275496
rect 255558 275440 255563 275496
rect 253460 275438 255563 275440
rect 255497 275435 255563 275438
rect 101254 275362 101260 275364
rect 98716 275302 101260 275362
rect 101254 275300 101260 275302
rect 101324 275300 101330 275364
rect 258574 275226 258580 275228
rect 258030 275166 258580 275226
rect 255313 275090 255379 275093
rect 253460 275088 255379 275090
rect 253460 275032 255318 275088
rect 255374 275032 255379 275088
rect 253460 275030 255379 275032
rect 255313 275027 255379 275030
rect 258030 274954 258090 275166
rect 258574 275164 258580 275166
rect 258644 275226 258650 275228
rect 270493 275226 270559 275229
rect 258644 275224 270559 275226
rect 258644 275168 270498 275224
rect 270554 275168 270559 275224
rect 258644 275166 270559 275168
rect 258644 275164 258650 275166
rect 270493 275163 270559 275166
rect 253430 274894 258090 274954
rect 66713 274818 66779 274821
rect 190545 274818 190611 274821
rect 66713 274816 68908 274818
rect 66713 274760 66718 274816
rect 66774 274760 68908 274816
rect 66713 274758 68908 274760
rect 190545 274816 193660 274818
rect 190545 274760 190550 274816
rect 190606 274760 193660 274816
rect 190545 274758 193660 274760
rect 66713 274755 66779 274758
rect 190545 274755 190611 274758
rect 253430 274652 253490 274894
rect 100753 274546 100819 274549
rect 98716 274544 100819 274546
rect 98716 274488 100758 274544
rect 100814 274488 100819 274544
rect 98716 274486 100819 274488
rect 100753 274483 100819 274486
rect 255497 274274 255563 274277
rect 253460 274272 255563 274274
rect 253460 274216 255502 274272
rect 255558 274216 255563 274272
rect 253460 274214 255563 274216
rect 255497 274211 255563 274214
rect 66805 274002 66871 274005
rect 66805 274000 68908 274002
rect 66805 273944 66810 274000
rect 66866 273944 68908 274000
rect 66805 273942 68908 273944
rect 66805 273939 66871 273942
rect 255313 273866 255379 273869
rect 270585 273866 270651 273869
rect 253460 273864 255379 273866
rect 253460 273808 255318 273864
rect 255374 273808 255379 273864
rect 253460 273806 255379 273808
rect 255313 273803 255379 273806
rect 267690 273864 270651 273866
rect 267690 273808 270590 273864
rect 270646 273808 270651 273864
rect 267690 273806 270651 273808
rect 100845 273730 100911 273733
rect 98716 273728 100911 273730
rect 98716 273672 100850 273728
rect 100906 273672 100911 273728
rect 98716 273670 100911 273672
rect 100845 273667 100911 273670
rect 190453 273730 190519 273733
rect 190453 273728 193660 273730
rect 190453 273672 190458 273728
rect 190514 273672 193660 273728
rect 190453 273670 193660 273672
rect 190453 273667 190519 273670
rect 263777 273594 263843 273597
rect 267690 273594 267750 273806
rect 270585 273803 270651 273806
rect 253430 273592 267750 273594
rect 253430 273536 263782 273592
rect 263838 273536 267750 273592
rect 253430 273534 267750 273536
rect 253430 273428 253490 273534
rect 263777 273531 263843 273534
rect 65701 273186 65767 273189
rect 66069 273186 66135 273189
rect 255313 273186 255379 273189
rect 277393 273186 277459 273189
rect 278681 273186 278747 273189
rect 65701 273184 68908 273186
rect 65701 273128 65706 273184
rect 65762 273128 66074 273184
rect 66130 273128 68908 273184
rect 65701 273126 68908 273128
rect 255313 273184 278747 273186
rect 255313 273128 255318 273184
rect 255374 273128 277398 273184
rect 277454 273128 278686 273184
rect 278742 273128 278747 273184
rect 255313 273126 278747 273128
rect 65701 273123 65767 273126
rect 66069 273123 66135 273126
rect 255313 273123 255379 273126
rect 277393 273123 277459 273126
rect 278681 273123 278747 273126
rect 100753 272914 100819 272917
rect 98716 272912 100819 272914
rect 98716 272856 100758 272912
rect 100814 272856 100819 272912
rect 98716 272854 100819 272856
rect 100753 272851 100819 272854
rect 253430 272778 253490 272884
rect 258073 272778 258139 272781
rect 260925 272778 260991 272781
rect 253430 272776 260991 272778
rect 253430 272720 258078 272776
rect 258134 272720 260930 272776
rect 260986 272720 260991 272776
rect 253430 272718 260991 272720
rect 258073 272715 258139 272718
rect 260925 272715 260991 272718
rect 190821 272642 190887 272645
rect 190821 272640 193660 272642
rect 190821 272584 190826 272640
rect 190882 272584 193660 272640
rect 190821 272582 193660 272584
rect 190821 272579 190887 272582
rect 255497 272506 255563 272509
rect 253460 272504 255563 272506
rect 253460 272448 255502 272504
rect 255558 272448 255563 272504
rect 253460 272446 255563 272448
rect 255497 272443 255563 272446
rect 66805 272370 66871 272373
rect 66805 272368 68908 272370
rect 66805 272312 66810 272368
rect 66866 272312 68908 272368
rect 66805 272310 68908 272312
rect 66805 272307 66871 272310
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 101397 272098 101463 272101
rect 255313 272098 255379 272101
rect 98716 272096 101463 272098
rect 98716 272040 101402 272096
rect 101458 272040 101463 272096
rect 98716 272038 101463 272040
rect 253460 272096 255379 272098
rect 253460 272040 255318 272096
rect 255374 272040 255379 272096
rect 583520 272084 584960 272174
rect 253460 272038 255379 272040
rect 101397 272035 101463 272038
rect 255313 272035 255379 272038
rect 262213 271826 262279 271829
rect 266445 271826 266511 271829
rect 262213 271824 266511 271826
rect 262213 271768 262218 271824
rect 262274 271768 266450 271824
rect 266506 271768 266511 271824
rect 262213 271766 266511 271768
rect 262213 271763 262279 271766
rect 266445 271763 266511 271766
rect 191649 271554 191715 271557
rect 253430 271554 253490 271660
rect 262213 271554 262279 271557
rect 191649 271552 193660 271554
rect 68878 271010 68938 271524
rect 191649 271496 191654 271552
rect 191710 271496 193660 271552
rect 191649 271494 193660 271496
rect 253430 271552 262279 271554
rect 253430 271496 262218 271552
rect 262274 271496 262279 271552
rect 253430 271494 262279 271496
rect 191649 271491 191715 271494
rect 262213 271491 262279 271494
rect 101121 271282 101187 271285
rect 255497 271282 255563 271285
rect 98716 271280 101187 271282
rect 98716 271224 101126 271280
rect 101182 271224 101187 271280
rect 98716 271222 101187 271224
rect 253460 271280 255563 271282
rect 253460 271224 255502 271280
rect 255558 271224 255563 271280
rect 253460 271222 255563 271224
rect 101121 271219 101187 271222
rect 255497 271219 255563 271222
rect 64830 270950 68938 271010
rect 54753 270738 54819 270741
rect 64830 270738 64890 270950
rect 255497 270874 255563 270877
rect 253460 270872 255563 270874
rect 253460 270816 255502 270872
rect 255558 270816 255563 270872
rect 253460 270814 255563 270816
rect 255497 270811 255563 270814
rect 54753 270736 64890 270738
rect 54753 270680 54758 270736
rect 54814 270680 64890 270736
rect 54753 270678 64890 270680
rect 66805 270738 66871 270741
rect 66805 270736 68908 270738
rect 66805 270680 66810 270736
rect 66866 270680 68908 270736
rect 66805 270678 68908 270680
rect 54753 270675 54819 270678
rect 66805 270675 66871 270678
rect 99966 270466 99972 270468
rect 98716 270406 99972 270466
rect 99966 270404 99972 270406
rect 100036 270466 100042 270468
rect 100753 270466 100819 270469
rect 100036 270464 100819 270466
rect 100036 270408 100758 270464
rect 100814 270408 100819 270464
rect 100036 270406 100819 270408
rect 100036 270404 100042 270406
rect 100753 270403 100819 270406
rect 190821 270466 190887 270469
rect 255497 270466 255563 270469
rect 190821 270464 193660 270466
rect 190821 270408 190826 270464
rect 190882 270408 193660 270464
rect 190821 270406 193660 270408
rect 253460 270464 255563 270466
rect 253460 270408 255502 270464
rect 255558 270408 255563 270464
rect 253460 270406 255563 270408
rect 190821 270403 190887 270406
rect 255497 270403 255563 270406
rect 66621 269922 66687 269925
rect 255313 269922 255379 269925
rect 66621 269920 68908 269922
rect 66621 269864 66626 269920
rect 66682 269864 68908 269920
rect 66621 269862 68908 269864
rect 253460 269920 255379 269922
rect 253460 269864 255318 269920
rect 255374 269864 255379 269920
rect 253460 269862 255379 269864
rect 66621 269859 66687 269862
rect 255313 269859 255379 269862
rect 265249 269786 265315 269789
rect 295333 269786 295399 269789
rect 265249 269784 295399 269786
rect 265249 269728 265254 269784
rect 265310 269728 295338 269784
rect 295394 269728 295399 269784
rect 265249 269726 295399 269728
rect 265249 269723 265315 269726
rect 295333 269723 295399 269726
rect 98686 269378 98746 269620
rect 113265 269378 113331 269381
rect 98686 269376 113331 269378
rect 98686 269320 113270 269376
rect 113326 269320 113331 269376
rect 98686 269318 113331 269320
rect 113265 269315 113331 269318
rect 191557 269378 191623 269381
rect 253430 269378 253490 269484
rect 265249 269378 265315 269381
rect 191557 269376 193660 269378
rect 191557 269320 191562 269376
rect 191618 269320 193660 269376
rect 191557 269318 193660 269320
rect 253430 269376 265315 269378
rect 253430 269320 265254 269376
rect 265310 269320 265315 269376
rect 253430 269318 265315 269320
rect 191557 269315 191623 269318
rect 265249 269315 265315 269318
rect 66161 269106 66227 269109
rect 256601 269106 256667 269109
rect 66161 269104 68908 269106
rect 66161 269048 66166 269104
rect 66222 269048 68908 269104
rect 66161 269046 68908 269048
rect 253460 269104 256667 269106
rect 253460 269048 256606 269104
rect 256662 269048 256667 269104
rect 253460 269046 256667 269048
rect 66161 269043 66227 269046
rect 256601 269043 256667 269046
rect 100937 268834 101003 268837
rect 98716 268832 101003 268834
rect 98716 268776 100942 268832
rect 100998 268776 101003 268832
rect 98716 268774 101003 268776
rect 100937 268771 101003 268774
rect 253430 268562 253490 268668
rect 292573 268562 292639 268565
rect 253430 268560 292639 268562
rect 253430 268504 292578 268560
rect 292634 268504 292639 268560
rect 253430 268502 292639 268504
rect 292573 268499 292639 268502
rect 66805 268290 66871 268293
rect 191649 268290 191715 268293
rect 66805 268288 68908 268290
rect 66805 268232 66810 268288
rect 66866 268232 68908 268288
rect 66805 268230 68908 268232
rect 191649 268288 193660 268290
rect 191649 268232 191654 268288
rect 191710 268232 193660 268288
rect 191649 268230 193660 268232
rect 66805 268227 66871 268230
rect 191649 268227 191715 268230
rect 253430 268154 253490 268260
rect 273345 268154 273411 268157
rect 277393 268154 277459 268157
rect 253430 268152 277459 268154
rect 253430 268096 273350 268152
rect 273406 268096 277398 268152
rect 277454 268096 277459 268152
rect 253430 268094 277459 268096
rect 273345 268091 273411 268094
rect 277393 268091 277459 268094
rect 100753 268018 100819 268021
rect 98164 268016 100819 268018
rect 98164 267988 100758 268016
rect 98134 267960 100758 267988
rect 100814 267960 100819 268016
rect 98134 267958 100819 267960
rect 98134 267884 98194 267958
rect 100753 267955 100819 267958
rect 98126 267820 98132 267884
rect 98196 267820 98202 267884
rect 255497 267882 255563 267885
rect 253460 267880 255563 267882
rect 253460 267824 255502 267880
rect 255558 267824 255563 267880
rect 253460 267822 255563 267824
rect 255497 267819 255563 267822
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 68878 266930 68938 267444
rect 253430 267202 253490 267444
rect 64830 266870 68938 266930
rect 49601 266522 49667 266525
rect 64830 266522 64890 266870
rect 66805 266658 66871 266661
rect 98686 266658 98746 267172
rect 117313 266658 117379 266661
rect 66805 266656 68908 266658
rect 66805 266600 66810 266656
rect 66866 266600 68908 266656
rect 66805 266598 68908 266600
rect 98686 266656 117379 266658
rect 98686 266600 117318 266656
rect 117374 266600 117379 266656
rect 98686 266598 117379 266600
rect 66805 266595 66871 266598
rect 117313 266595 117379 266598
rect 49601 266520 64890 266522
rect 49601 266464 49606 266520
rect 49662 266464 64890 266520
rect 49601 266462 64890 266464
rect 49601 266459 49667 266462
rect 100753 266386 100819 266389
rect 98716 266384 100819 266386
rect 98716 266328 100758 266384
rect 100814 266328 100819 266384
rect 98716 266326 100819 266328
rect 100753 266323 100819 266326
rect 151077 266386 151143 266389
rect 193630 266386 193690 267172
rect 253430 267142 258090 267202
rect 255313 266930 255379 266933
rect 253460 266928 255379 266930
rect 253460 266872 255318 266928
rect 255374 266872 255379 266928
rect 253460 266870 255379 266872
rect 255313 266867 255379 266870
rect 258030 266794 258090 267142
rect 270769 266794 270835 266797
rect 258030 266792 270835 266794
rect 258030 266736 270774 266792
rect 270830 266736 270835 266792
rect 258030 266734 270835 266736
rect 270769 266731 270835 266734
rect 261017 266522 261083 266525
rect 253460 266520 261083 266522
rect 253460 266464 261022 266520
rect 261078 266464 261083 266520
rect 253460 266462 261083 266464
rect 261017 266459 261083 266462
rect 151077 266384 193690 266386
rect 151077 266328 151082 266384
rect 151138 266328 193690 266384
rect 151077 266326 193690 266328
rect 151077 266323 151143 266326
rect 191649 266114 191715 266117
rect 255497 266114 255563 266117
rect 191649 266112 193660 266114
rect 191649 266056 191654 266112
rect 191710 266056 193660 266112
rect 191649 266054 193660 266056
rect 253460 266112 255563 266114
rect 253460 266056 255502 266112
rect 255558 266056 255563 266112
rect 253460 266054 255563 266056
rect 191649 266051 191715 266054
rect 255497 266051 255563 266054
rect 68878 265298 68938 265812
rect 255497 265706 255563 265709
rect 253460 265704 255563 265706
rect 253460 265648 255502 265704
rect 255558 265648 255563 265704
rect 253460 265646 255563 265648
rect 255497 265643 255563 265646
rect 100753 265570 100819 265573
rect 98716 265568 100819 265570
rect 98716 265512 100758 265568
rect 100814 265512 100819 265568
rect 98716 265510 100819 265512
rect 100753 265507 100819 265510
rect 148174 265508 148180 265572
rect 148244 265570 148250 265572
rect 163681 265570 163747 265573
rect 148244 265568 163747 265570
rect 148244 265512 163686 265568
rect 163742 265512 163747 265568
rect 148244 265510 163747 265512
rect 148244 265508 148250 265510
rect 163681 265507 163747 265510
rect 64830 265238 68938 265298
rect 54845 265026 54911 265029
rect 64830 265026 64890 265238
rect 253430 265162 253490 265268
rect 273345 265162 273411 265165
rect 253430 265160 273411 265162
rect 253430 265104 273350 265160
rect 273406 265104 273411 265160
rect 253430 265102 273411 265104
rect 273345 265099 273411 265102
rect 54845 265024 64890 265026
rect 54845 264968 54850 265024
rect 54906 264968 64890 265024
rect 54845 264966 64890 264968
rect 66529 265026 66595 265029
rect 190821 265026 190887 265029
rect 66529 265024 68908 265026
rect 66529 264968 66534 265024
rect 66590 264968 68908 265024
rect 66529 264966 68908 264968
rect 190821 265024 193660 265026
rect 190821 264968 190826 265024
rect 190882 264968 193660 265024
rect 190821 264966 193660 264968
rect 54845 264963 54911 264966
rect 66529 264963 66595 264966
rect 190821 264963 190887 264966
rect 255313 264890 255379 264893
rect 253460 264888 255379 264890
rect 253460 264832 255318 264888
rect 255374 264832 255379 264888
rect 253460 264830 255379 264832
rect 255313 264827 255379 264830
rect 100845 264754 100911 264757
rect 98716 264752 100911 264754
rect 98716 264696 100850 264752
rect 100906 264696 100911 264752
rect 98716 264694 100911 264696
rect 100845 264691 100911 264694
rect 260833 264482 260899 264485
rect 260966 264482 260972 264484
rect 260833 264480 260972 264482
rect 260833 264424 260838 264480
rect 260894 264424 260972 264480
rect 260833 264422 260972 264424
rect 260833 264419 260899 264422
rect 260966 264420 260972 264422
rect 261036 264420 261042 264484
rect 260966 264346 260972 264348
rect 253460 264286 260972 264346
rect 260966 264284 260972 264286
rect 261036 264284 261042 264348
rect 66805 264210 66871 264213
rect 66805 264208 68908 264210
rect 66805 264152 66810 264208
rect 66866 264152 68908 264208
rect 66805 264150 68908 264152
rect 66805 264147 66871 264150
rect 262254 264148 262260 264212
rect 262324 264210 262330 264212
rect 284334 264210 284340 264212
rect 262324 264150 284340 264210
rect 262324 264148 262330 264150
rect 284334 264148 284340 264150
rect 284404 264148 284410 264212
rect 191649 263938 191715 263941
rect 255497 263938 255563 263941
rect 191649 263936 193660 263938
rect 98686 263666 98746 263908
rect 191649 263880 191654 263936
rect 191710 263880 193660 263936
rect 191649 263878 193660 263880
rect 253460 263936 255563 263938
rect 253460 263880 255502 263936
rect 255558 263880 255563 263936
rect 253460 263878 255563 263880
rect 191649 263875 191715 263878
rect 255497 263875 255563 263878
rect 130653 263666 130719 263669
rect 98686 263664 130719 263666
rect 98686 263608 130658 263664
rect 130714 263608 130719 263664
rect 98686 263606 130719 263608
rect 130653 263603 130719 263606
rect 256417 263530 256483 263533
rect 253460 263528 256483 263530
rect 253460 263472 256422 263528
rect 256478 263472 256483 263528
rect 253460 263470 256483 263472
rect 256417 263467 256483 263470
rect 67081 263394 67147 263397
rect 67449 263394 67515 263397
rect 265801 263394 265867 263397
rect 269246 263394 269252 263396
rect 67081 263392 68908 263394
rect 67081 263336 67086 263392
rect 67142 263336 67454 263392
rect 67510 263336 68908 263392
rect 67081 263334 68908 263336
rect 265801 263392 269252 263394
rect 265801 263336 265806 263392
rect 265862 263336 269252 263392
rect 265801 263334 269252 263336
rect 67081 263331 67147 263334
rect 67449 263331 67515 263334
rect 265801 263331 265867 263334
rect 269246 263332 269252 263334
rect 269316 263332 269322 263396
rect 100753 263122 100819 263125
rect 256877 263122 256943 263125
rect 98716 263120 100819 263122
rect 98716 263064 100758 263120
rect 100814 263064 100819 263120
rect 98716 263062 100819 263064
rect 253460 263120 256943 263122
rect 253460 263064 256882 263120
rect 256938 263064 256943 263120
rect 253460 263062 256943 263064
rect 100753 263059 100819 263062
rect 256877 263059 256943 263062
rect 191649 262850 191715 262853
rect 263777 262850 263843 262853
rect 270534 262850 270540 262852
rect 191649 262848 193660 262850
rect 191649 262792 191654 262848
rect 191710 262792 193660 262848
rect 191649 262790 193660 262792
rect 263777 262848 270540 262850
rect 263777 262792 263782 262848
rect 263838 262792 270540 262848
rect 263777 262790 270540 262792
rect 191649 262787 191715 262790
rect 263777 262787 263843 262790
rect 270534 262788 270540 262790
rect 270604 262788 270610 262852
rect 263869 262714 263935 262717
rect 265750 262714 265756 262716
rect 253890 262712 265756 262714
rect 66529 262578 66595 262581
rect 253430 262578 253490 262684
rect 253890 262656 263874 262712
rect 263930 262656 265756 262712
rect 253890 262654 265756 262656
rect 253890 262578 253950 262654
rect 263869 262651 263935 262654
rect 265750 262652 265756 262654
rect 265820 262652 265826 262716
rect 66529 262576 68908 262578
rect 66529 262520 66534 262576
rect 66590 262520 68908 262576
rect 66529 262518 68908 262520
rect 253430 262518 253950 262578
rect 66529 262515 66595 262518
rect 100661 262306 100727 262309
rect 100937 262306 101003 262309
rect 263542 262306 263548 262308
rect 98716 262304 101003 262306
rect 98716 262248 100666 262304
rect 100722 262248 100942 262304
rect 100998 262248 101003 262304
rect 98716 262246 101003 262248
rect 253460 262246 263548 262306
rect 100661 262243 100727 262246
rect 100937 262243 101003 262246
rect 263542 262244 263548 262246
rect 263612 262244 263618 262308
rect 280245 262172 280311 262173
rect 280245 262168 280292 262172
rect 280356 262170 280362 262172
rect 280245 262112 280250 262168
rect 280245 262108 280292 262112
rect 280356 262110 280402 262170
rect 280356 262108 280362 262110
rect 280245 262107 280311 262108
rect 191649 261762 191715 261765
rect 191649 261760 193660 261762
rect 68878 261218 68938 261732
rect 191649 261704 191654 261760
rect 191710 261704 193660 261760
rect 191649 261702 193660 261704
rect 191649 261699 191715 261702
rect 253430 261626 253490 261868
rect 263174 261626 263180 261628
rect 253430 261566 263180 261626
rect 263174 261564 263180 261566
rect 263244 261564 263250 261628
rect 102225 261490 102291 261493
rect 98348 261488 102291 261490
rect 98348 261460 102230 261488
rect 98318 261432 102230 261460
rect 102286 261432 102291 261488
rect 98318 261430 102291 261432
rect 98177 261354 98243 261357
rect 98318 261354 98378 261430
rect 102225 261427 102291 261430
rect 256601 261354 256667 261357
rect 98177 261352 98378 261354
rect 98177 261296 98182 261352
rect 98238 261296 98378 261352
rect 98177 261294 98378 261296
rect 253460 261352 256667 261354
rect 253460 261296 256606 261352
rect 256662 261296 256667 261352
rect 253460 261294 256667 261296
rect 98177 261291 98243 261294
rect 256601 261291 256667 261294
rect 64830 261158 68938 261218
rect 61009 260946 61075 260949
rect 64830 260946 64890 261158
rect 61009 260944 64890 260946
rect 61009 260888 61014 260944
rect 61070 260888 64890 260944
rect 61009 260886 64890 260888
rect 66253 260946 66319 260949
rect 263777 260946 263843 260949
rect 66253 260944 68908 260946
rect 66253 260888 66258 260944
rect 66314 260888 68908 260944
rect 66253 260886 68908 260888
rect 253460 260944 263843 260946
rect 253460 260888 263782 260944
rect 263838 260888 263843 260944
rect 253460 260886 263843 260888
rect 61009 260883 61075 260886
rect 66253 260883 66319 260886
rect 263777 260883 263843 260886
rect 107009 260810 107075 260813
rect 109677 260810 109743 260813
rect 107009 260808 109743 260810
rect 107009 260752 107014 260808
rect 107070 260752 109682 260808
rect 109738 260752 109743 260808
rect 107009 260750 109743 260752
rect 107009 260747 107075 260750
rect 109677 260747 109743 260750
rect 269062 260748 269068 260812
rect 269132 260810 269138 260812
rect 273294 260810 273300 260812
rect 269132 260750 273300 260810
rect 269132 260748 269138 260750
rect 273294 260748 273300 260750
rect 273364 260748 273370 260812
rect 100845 260674 100911 260677
rect 98716 260672 100911 260674
rect 98716 260616 100850 260672
rect 100906 260616 100911 260672
rect 98716 260614 100911 260616
rect 100845 260611 100911 260614
rect 191649 260674 191715 260677
rect 191649 260672 193660 260674
rect 191649 260616 191654 260672
rect 191710 260616 193660 260672
rect 191649 260614 193660 260616
rect 191649 260611 191715 260614
rect 258390 260538 258396 260540
rect 253460 260478 258396 260538
rect 258390 260476 258396 260478
rect 258460 260476 258466 260540
rect 66529 260130 66595 260133
rect 256601 260130 256667 260133
rect 66529 260128 68908 260130
rect 66529 260072 66534 260128
rect 66590 260072 68908 260128
rect 66529 260070 68908 260072
rect 253460 260128 256667 260130
rect 253460 260072 256606 260128
rect 256662 260072 256667 260128
rect 253460 260070 256667 260072
rect 66529 260067 66595 260070
rect 256601 260067 256667 260070
rect 263225 260130 263291 260133
rect 263358 260130 263364 260132
rect 263225 260128 263364 260130
rect 263225 260072 263230 260128
rect 263286 260072 263364 260128
rect 263225 260070 263364 260072
rect 263225 260067 263291 260070
rect 263358 260068 263364 260070
rect 263428 260130 263434 260132
rect 265750 260130 265756 260132
rect 263428 260070 265756 260130
rect 263428 260068 263434 260070
rect 265750 260068 265756 260070
rect 265820 260068 265826 260132
rect 262254 259994 262260 259996
rect 253430 259934 262260 259994
rect 100753 259858 100819 259861
rect 98716 259856 100819 259858
rect 98716 259800 100758 259856
rect 100814 259800 100819 259856
rect 98716 259798 100819 259800
rect 100753 259795 100819 259798
rect 253430 259692 253490 259934
rect 262254 259932 262260 259934
rect 262324 259932 262330 259996
rect 171777 259586 171843 259589
rect 285673 259588 285739 259589
rect 285622 259586 285628 259588
rect 171777 259584 193660 259586
rect 171777 259528 171782 259584
rect 171838 259528 193660 259584
rect 171777 259526 193660 259528
rect 285582 259526 285628 259586
rect 285692 259584 285739 259588
rect 285734 259528 285739 259584
rect 171777 259523 171843 259526
rect 285622 259524 285628 259526
rect 285692 259524 285739 259528
rect 285673 259523 285739 259524
rect 265065 259450 265131 259453
rect 269062 259450 269068 259452
rect 265065 259448 269068 259450
rect 265065 259392 265070 259448
rect 265126 259392 269068 259448
rect 265065 259390 269068 259392
rect 265065 259387 265131 259390
rect 269062 259388 269068 259390
rect 269132 259388 269138 259452
rect 271873 259450 271939 259453
rect 273294 259450 273300 259452
rect 271873 259448 273300 259450
rect 271873 259392 271878 259448
rect 271934 259392 273300 259448
rect 271873 259390 273300 259392
rect 271873 259387 271939 259390
rect 273294 259388 273300 259390
rect 273364 259450 273370 259452
rect 274582 259450 274588 259452
rect 273364 259390 274588 259450
rect 273364 259388 273370 259390
rect 274582 259388 274588 259390
rect 274652 259388 274658 259452
rect 255957 259314 256023 259317
rect 253460 259312 256023 259314
rect 68185 258770 68251 258773
rect 68878 258770 68938 259284
rect 253460 259256 255962 259312
rect 256018 259256 256023 259312
rect 253460 259254 256023 259256
rect 255957 259251 256023 259254
rect 100017 259042 100083 259045
rect 98716 259040 100083 259042
rect 98716 258984 100022 259040
rect 100078 258984 100083 259040
rect 98716 258982 100083 258984
rect 100017 258979 100083 258982
rect 256601 258906 256667 258909
rect 253460 258904 256667 258906
rect 253460 258848 256606 258904
rect 256662 258848 256667 258904
rect 253460 258846 256667 258848
rect 256601 258843 256667 258846
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 68185 258768 68938 258770
rect 68185 258712 68190 258768
rect 68246 258712 68938 258768
rect 68185 258710 68938 258712
rect 154481 258770 154547 258773
rect 191230 258770 191236 258772
rect 154481 258768 191236 258770
rect 154481 258712 154486 258768
rect 154542 258712 191236 258768
rect 154481 258710 191236 258712
rect 68185 258707 68251 258710
rect 154481 258707 154547 258710
rect 191230 258708 191236 258710
rect 191300 258708 191306 258772
rect 583520 258756 584960 258846
rect 60457 258226 60523 258229
rect 68878 258226 68938 258468
rect 100753 258226 100819 258229
rect 60457 258224 68938 258226
rect 60457 258168 60462 258224
rect 60518 258168 68938 258224
rect 60457 258166 68938 258168
rect 98716 258224 100819 258226
rect 98716 258168 100758 258224
rect 100814 258168 100819 258224
rect 98716 258166 100819 258168
rect 60457 258163 60523 258166
rect 99238 258093 99298 258166
rect 100753 258163 100819 258166
rect 99238 258088 99347 258093
rect 99238 258032 99286 258088
rect 99342 258032 99347 258088
rect 99238 258030 99347 258032
rect 99281 258027 99347 258030
rect 190453 258090 190519 258093
rect 190453 258088 190562 258090
rect 190453 258032 190458 258088
rect 190514 258032 190562 258088
rect 190453 258027 190562 258032
rect 190502 257954 190562 258027
rect 193630 257954 193690 258468
rect 253430 258226 253490 258332
rect 267774 258226 267780 258228
rect 253430 258166 267780 258226
rect 267774 258164 267780 258166
rect 267844 258164 267850 258228
rect 255814 257954 255820 257956
rect 190502 257894 193690 257954
rect 253460 257894 255820 257954
rect 255814 257892 255820 257894
rect 255884 257954 255890 257956
rect 259678 257954 259684 257956
rect 255884 257894 259684 257954
rect 255884 257892 255890 257894
rect 259678 257892 259684 257894
rect 259748 257892 259754 257956
rect 66437 257682 66503 257685
rect 66437 257680 68908 257682
rect 66437 257624 66442 257680
rect 66498 257624 68908 257680
rect 66437 257622 68908 257624
rect 66437 257619 66503 257622
rect 254526 257546 254532 257548
rect 253460 257486 254532 257546
rect 254526 257484 254532 257486
rect 254596 257546 254602 257548
rect 258257 257546 258323 257549
rect 254596 257544 258323 257546
rect 254596 257488 258262 257544
rect 258318 257488 258323 257544
rect 254596 257486 258323 257488
rect 254596 257484 254602 257486
rect 258257 257483 258323 257486
rect 102041 257410 102107 257413
rect 98716 257408 102107 257410
rect 98716 257352 102046 257408
rect 102102 257352 102107 257408
rect 98716 257350 102107 257352
rect 102041 257347 102107 257350
rect 191649 257410 191715 257413
rect 267733 257412 267799 257413
rect 191649 257408 193660 257410
rect 191649 257352 191654 257408
rect 191710 257352 193660 257408
rect 191649 257350 193660 257352
rect 267733 257408 267780 257412
rect 267844 257410 267850 257412
rect 267733 257352 267738 257408
rect 191649 257347 191715 257350
rect 267733 257348 267780 257352
rect 267844 257350 267890 257410
rect 267844 257348 267850 257350
rect 267733 257347 267799 257348
rect 256325 257138 256391 257141
rect 253460 257136 256391 257138
rect 253460 257080 256330 257136
rect 256386 257080 256391 257136
rect 253460 257078 256391 257080
rect 256325 257075 256391 257078
rect 66529 256730 66595 256733
rect 66662 256730 66668 256732
rect 66529 256728 66668 256730
rect 66529 256672 66534 256728
rect 66590 256672 66668 256728
rect 66529 256670 66668 256672
rect 66529 256667 66595 256670
rect 66662 256668 66668 256670
rect 66732 256730 66738 256732
rect 68878 256730 68938 256836
rect 256601 256730 256667 256733
rect 66732 256670 68938 256730
rect 253460 256728 256667 256730
rect 253460 256672 256606 256728
rect 256662 256672 256667 256728
rect 253460 256670 256667 256672
rect 66732 256668 66738 256670
rect 256601 256667 256667 256670
rect 100753 256594 100819 256597
rect 98716 256592 100819 256594
rect 98716 256536 100758 256592
rect 100814 256536 100819 256592
rect 98716 256534 100819 256536
rect 100753 256531 100819 256534
rect 190637 256322 190703 256325
rect 256601 256322 256667 256325
rect 190637 256320 193660 256322
rect 190637 256264 190642 256320
rect 190698 256264 193660 256320
rect 190637 256262 193660 256264
rect 253460 256320 256667 256322
rect 253460 256264 256606 256320
rect 256662 256264 256667 256320
rect 253460 256262 256667 256264
rect 190637 256259 190703 256262
rect 256601 256259 256667 256262
rect 68878 255506 68938 256020
rect 100845 255778 100911 255781
rect 258165 255778 258231 255781
rect 98716 255776 100911 255778
rect 98716 255720 100850 255776
rect 100906 255720 100911 255776
rect 98716 255718 100911 255720
rect 253460 255776 258231 255778
rect 253460 255720 258170 255776
rect 258226 255720 258231 255776
rect 253460 255718 258231 255720
rect 100845 255715 100911 255718
rect 258165 255715 258231 255718
rect 68510 255446 68938 255506
rect 66110 255308 66116 255372
rect 66180 255370 66186 255372
rect 66253 255370 66319 255373
rect 68510 255370 68570 255446
rect 66180 255368 68570 255370
rect 66180 255312 66258 255368
rect 66314 255312 68570 255368
rect 66180 255310 68570 255312
rect 66180 255308 66186 255310
rect 66253 255307 66319 255310
rect 177246 255308 177252 255372
rect 177316 255370 177322 255372
rect 178953 255370 179019 255373
rect 256601 255370 256667 255373
rect 177316 255368 179019 255370
rect 177316 255312 178958 255368
rect 179014 255312 179019 255368
rect 177316 255310 179019 255312
rect 253460 255368 256667 255370
rect 253460 255312 256606 255368
rect 256662 255312 256667 255368
rect 253460 255310 256667 255312
rect 177316 255308 177322 255310
rect 178953 255307 179019 255310
rect 256601 255307 256667 255310
rect 276381 255372 276447 255373
rect 276381 255368 276428 255372
rect 276492 255370 276498 255372
rect 276381 255312 276386 255368
rect 276381 255308 276428 255312
rect 276492 255310 276538 255370
rect 276492 255308 276498 255310
rect 276381 255307 276447 255308
rect 66805 255234 66871 255237
rect 191649 255234 191715 255237
rect 269430 255234 269436 255236
rect 66805 255232 68908 255234
rect 66805 255176 66810 255232
rect 66866 255176 68908 255232
rect 66805 255174 68908 255176
rect 191649 255232 193660 255234
rect 191649 255176 191654 255232
rect 191710 255176 193660 255232
rect 191649 255174 193660 255176
rect 253430 255174 269436 255234
rect 66805 255171 66871 255174
rect 191649 255171 191715 255174
rect 100569 254962 100635 254965
rect 100753 254962 100819 254965
rect 98716 254960 100819 254962
rect 98716 254904 100574 254960
rect 100630 254904 100758 254960
rect 100814 254904 100819 254960
rect 253430 254932 253490 255174
rect 269430 255172 269436 255174
rect 269500 255234 269506 255236
rect 270534 255234 270540 255236
rect 269500 255174 270540 255234
rect 269500 255172 269506 255174
rect 270534 255172 270540 255174
rect 270604 255172 270610 255236
rect 98716 254902 100819 254904
rect 100569 254899 100635 254902
rect 100753 254899 100819 254902
rect 130653 254554 130719 254557
rect 184197 254554 184263 254557
rect 256601 254554 256667 254557
rect 130653 254552 184263 254554
rect 130653 254496 130658 254552
rect 130714 254496 184202 254552
rect 184258 254496 184263 254552
rect 130653 254494 184263 254496
rect 253460 254552 256667 254554
rect 253460 254496 256606 254552
rect 256662 254496 256667 254552
rect 253460 254494 256667 254496
rect 130653 254491 130719 254494
rect 184197 254491 184263 254494
rect 256601 254491 256667 254494
rect 66805 254418 66871 254421
rect 66805 254416 68908 254418
rect 66805 254360 66810 254416
rect 66866 254360 68908 254416
rect 66805 254358 68908 254360
rect 66805 254355 66871 254358
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect 100753 254146 100819 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect 98716 254144 100819 254146
rect 98716 254088 100758 254144
rect 100814 254088 100819 254144
rect 98716 254086 100819 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 100753 254083 100819 254086
rect 191557 254146 191623 254149
rect 259729 254146 259795 254149
rect 191557 254144 193660 254146
rect 191557 254088 191562 254144
rect 191618 254088 193660 254144
rect 191557 254086 193660 254088
rect 253460 254144 259795 254146
rect 253460 254088 259734 254144
rect 259790 254088 259795 254144
rect 253460 254086 259795 254088
rect 191557 254083 191623 254086
rect 259729 254083 259795 254086
rect 184974 253948 184980 254012
rect 185044 254010 185050 254012
rect 186037 254010 186103 254013
rect 185044 254008 186103 254010
rect 185044 253952 186042 254008
rect 186098 253952 186103 254008
rect 185044 253950 186103 253952
rect 185044 253948 185050 253950
rect 186037 253947 186103 253950
rect 252870 253948 252876 254012
rect 252940 253948 252946 254012
rect 252878 253738 252938 253948
rect 260925 253738 260991 253741
rect 252878 253736 260991 253738
rect 252878 253708 260930 253736
rect 252908 253680 260930 253708
rect 260986 253680 260991 253736
rect 252908 253678 260991 253680
rect 260925 253675 260991 253678
rect 66989 253602 67055 253605
rect 66989 253600 68908 253602
rect 66989 253544 66994 253600
rect 67050 253544 68908 253600
rect 66989 253542 68908 253544
rect 66989 253539 67055 253542
rect 100753 253330 100819 253333
rect 255773 253330 255839 253333
rect 98716 253328 100819 253330
rect 98716 253272 100758 253328
rect 100814 253272 100819 253328
rect 98716 253270 100819 253272
rect 253460 253328 255839 253330
rect 253460 253272 255778 253328
rect 255834 253272 255839 253328
rect 253460 253270 255839 253272
rect 100753 253267 100819 253270
rect 255773 253267 255839 253270
rect 285765 253194 285831 253197
rect 267690 253192 285831 253194
rect 267690 253136 285770 253192
rect 285826 253136 285831 253192
rect 267690 253134 285831 253136
rect 191649 253058 191715 253061
rect 191649 253056 193660 253058
rect 191649 253000 191654 253056
rect 191710 253000 193660 253056
rect 191649 252998 193660 253000
rect 191649 252995 191715 252998
rect 63033 252786 63099 252789
rect 64689 252786 64755 252789
rect 254117 252786 254183 252789
rect 63033 252784 68908 252786
rect 63033 252728 63038 252784
rect 63094 252728 64694 252784
rect 64750 252728 68908 252784
rect 63033 252726 68908 252728
rect 253460 252784 254183 252786
rect 253460 252728 254122 252784
rect 254178 252728 254183 252784
rect 253460 252726 254183 252728
rect 63033 252723 63099 252726
rect 64689 252723 64755 252726
rect 254117 252723 254183 252726
rect 266486 252650 266492 252652
rect 256558 252590 266492 252650
rect 100702 252514 100708 252516
rect 98716 252454 100708 252514
rect 100702 252452 100708 252454
rect 100772 252514 100778 252516
rect 100845 252514 100911 252517
rect 100772 252512 100911 252514
rect 100772 252456 100850 252512
rect 100906 252456 100911 252512
rect 100772 252454 100911 252456
rect 100772 252452 100778 252454
rect 100845 252451 100911 252454
rect 256417 252378 256483 252381
rect 253460 252376 256483 252378
rect 253460 252320 256422 252376
rect 256478 252320 256483 252376
rect 253460 252318 256483 252320
rect 256417 252315 256483 252318
rect 256558 252242 256618 252590
rect 266486 252588 266492 252590
rect 266556 252650 266562 252652
rect 267690 252650 267750 253134
rect 285765 253131 285831 253134
rect 266556 252590 267750 252650
rect 266556 252588 266562 252590
rect 253430 252182 256618 252242
rect 66621 251970 66687 251973
rect 191649 251970 191715 251973
rect 66621 251968 68908 251970
rect 66621 251912 66626 251968
rect 66682 251912 68908 251968
rect 66621 251910 68908 251912
rect 191649 251968 193660 251970
rect 191649 251912 191654 251968
rect 191710 251912 193660 251968
rect 253430 251940 253490 252182
rect 191649 251910 193660 251912
rect 66621 251907 66687 251910
rect 191649 251907 191715 251910
rect 34329 251834 34395 251837
rect 66529 251834 66595 251837
rect 34329 251832 66595 251834
rect 34329 251776 34334 251832
rect 34390 251776 66534 251832
rect 66590 251776 66595 251832
rect 34329 251774 66595 251776
rect 34329 251771 34395 251774
rect 66529 251771 66595 251774
rect 100753 251698 100819 251701
rect 98716 251696 100819 251698
rect 98716 251640 100758 251696
rect 100814 251640 100819 251696
rect 98716 251638 100819 251640
rect 100753 251635 100819 251638
rect 254669 251562 254735 251565
rect 256601 251562 256667 251565
rect 253460 251560 256667 251562
rect 253460 251504 254674 251560
rect 254730 251504 256606 251560
rect 256662 251504 256667 251560
rect 253460 251502 256667 251504
rect 254669 251499 254735 251502
rect 256601 251499 256667 251502
rect 69062 250612 69122 251124
rect 253430 251018 253490 251124
rect 253430 250958 263610 251018
rect 100753 250882 100819 250885
rect 98716 250880 100819 250882
rect 98716 250824 100758 250880
rect 100814 250824 100819 250880
rect 98716 250822 100819 250824
rect 100753 250819 100819 250822
rect 190637 250882 190703 250885
rect 190637 250880 193660 250882
rect 190637 250824 190642 250880
rect 190698 250824 193660 250880
rect 190637 250822 193660 250824
rect 190637 250819 190703 250822
rect 256601 250746 256667 250749
rect 253460 250744 256667 250746
rect 253460 250688 256606 250744
rect 256662 250688 256667 250744
rect 253460 250686 256667 250688
rect 256601 250683 256667 250686
rect 69054 250548 69060 250612
rect 69124 250548 69130 250612
rect 101254 250412 101260 250476
rect 101324 250474 101330 250476
rect 149789 250474 149855 250477
rect 101324 250472 149855 250474
rect 101324 250416 149794 250472
rect 149850 250416 149855 250472
rect 101324 250414 149855 250416
rect 101324 250412 101330 250414
rect 149789 250411 149855 250414
rect 66805 250338 66871 250341
rect 256601 250338 256667 250341
rect 66805 250336 68908 250338
rect 66805 250280 66810 250336
rect 66866 250280 68908 250336
rect 66805 250278 68908 250280
rect 253460 250336 256667 250338
rect 253460 250280 256606 250336
rect 256662 250280 256667 250336
rect 253460 250278 256667 250280
rect 66805 250275 66871 250278
rect 256601 250275 256667 250278
rect 263550 250202 263610 250958
rect 582649 250474 582715 250477
rect 277350 250472 582715 250474
rect 277350 250416 582654 250472
rect 582710 250416 582715 250472
rect 277350 250414 582715 250416
rect 274909 250202 274975 250205
rect 277350 250202 277410 250414
rect 582649 250411 582715 250414
rect 263550 250200 277410 250202
rect 263550 250144 274914 250200
rect 274970 250144 277410 250200
rect 263550 250142 277410 250144
rect 274909 250139 274975 250142
rect 100845 250066 100911 250069
rect 98716 250064 100911 250066
rect 98716 250008 100850 250064
rect 100906 250008 100911 250064
rect 98716 250006 100911 250008
rect 100845 250003 100911 250006
rect 190821 249794 190887 249797
rect 254669 249794 254735 249797
rect 190821 249792 193660 249794
rect 190821 249736 190826 249792
rect 190882 249736 193660 249792
rect 190821 249734 193660 249736
rect 253460 249792 254735 249794
rect 253460 249736 254674 249792
rect 254730 249736 254735 249792
rect 253460 249734 254735 249736
rect 190821 249731 190887 249734
rect 254669 249731 254735 249734
rect 67817 249522 67883 249525
rect 67817 249520 68908 249522
rect 67817 249464 67822 249520
rect 67878 249464 68908 249520
rect 67817 249462 68908 249464
rect 67817 249459 67883 249462
rect 256233 249386 256299 249389
rect 253460 249384 256299 249386
rect 253460 249328 256238 249384
rect 256294 249328 256299 249384
rect 253460 249326 256299 249328
rect 256233 249323 256299 249326
rect 98318 248845 98378 249220
rect 256601 248978 256667 248981
rect 253460 248976 256667 248978
rect 253460 248920 256606 248976
rect 256662 248920 256667 248976
rect 253460 248918 256667 248920
rect 256601 248915 256667 248918
rect 98269 248840 98378 248845
rect 98269 248784 98274 248840
rect 98330 248784 98378 248840
rect 98269 248782 98378 248784
rect 98269 248779 98335 248782
rect 66805 248706 66871 248709
rect 283097 248706 283163 248709
rect 66805 248704 68908 248706
rect 66805 248648 66810 248704
rect 66866 248648 68908 248704
rect 253430 248704 283163 248706
rect 66805 248646 68908 248648
rect 66805 248643 66871 248646
rect 100937 248434 101003 248437
rect 98716 248432 101003 248434
rect 98716 248376 100942 248432
rect 100998 248376 101003 248432
rect 98716 248374 101003 248376
rect 100937 248371 101003 248374
rect 170254 248372 170260 248436
rect 170324 248434 170330 248436
rect 193630 248434 193690 248676
rect 253430 248648 283102 248704
rect 283158 248648 283163 248704
rect 253430 248646 283163 248648
rect 253430 248540 253490 248646
rect 283097 248643 283163 248646
rect 170324 248374 193690 248434
rect 170324 248372 170330 248374
rect 253430 248026 253490 248132
rect 253430 247966 267750 248026
rect 66529 247890 66595 247893
rect 66529 247888 68908 247890
rect 66529 247832 66534 247888
rect 66590 247832 68908 247888
rect 66529 247830 68908 247832
rect 66529 247827 66595 247830
rect 258390 247754 258396 247756
rect 253460 247694 258396 247754
rect 258390 247692 258396 247694
rect 258460 247692 258466 247756
rect 100109 247618 100175 247621
rect 98716 247616 100175 247618
rect 98716 247560 100114 247616
rect 100170 247560 100175 247616
rect 98716 247558 100175 247560
rect 100109 247555 100175 247558
rect 173341 247618 173407 247621
rect 184054 247618 184060 247620
rect 173341 247616 184060 247618
rect 173341 247560 173346 247616
rect 173402 247560 184060 247616
rect 173341 247558 184060 247560
rect 173341 247555 173407 247558
rect 184054 247556 184060 247558
rect 184124 247556 184130 247620
rect 66662 247012 66668 247076
rect 66732 247074 66738 247076
rect 189717 247074 189783 247077
rect 193630 247074 193690 247588
rect 267690 247482 267750 247966
rect 287053 247482 287119 247485
rect 287329 247482 287395 247485
rect 267690 247480 287395 247482
rect 267690 247424 287058 247480
rect 287114 247424 287334 247480
rect 287390 247424 287395 247480
rect 267690 247422 287395 247424
rect 287053 247419 287119 247422
rect 287329 247419 287395 247422
rect 256509 247210 256575 247213
rect 253460 247208 256575 247210
rect 253460 247152 256514 247208
rect 256570 247152 256575 247208
rect 253460 247150 256575 247152
rect 256509 247147 256575 247150
rect 66732 247014 68908 247074
rect 189717 247072 193690 247074
rect 189717 247016 189722 247072
rect 189778 247016 193690 247072
rect 189717 247014 193690 247016
rect 66732 247012 66738 247014
rect 189717 247011 189783 247014
rect 100937 246802 101003 246805
rect 256601 246802 256667 246805
rect 98716 246800 101003 246802
rect 98716 246744 100942 246800
rect 100998 246744 101003 246800
rect 98716 246742 101003 246744
rect 253460 246800 256667 246802
rect 253460 246744 256606 246800
rect 256662 246744 256667 246800
rect 253460 246742 256667 246744
rect 100937 246739 101003 246742
rect 256601 246739 256667 246742
rect 67449 246258 67515 246261
rect 101397 246258 101463 246261
rect 170489 246258 170555 246261
rect 67449 246256 68908 246258
rect 67449 246200 67454 246256
rect 67510 246200 68908 246256
rect 67449 246198 68908 246200
rect 98686 246256 170555 246258
rect 98686 246200 101402 246256
rect 101458 246200 170494 246256
rect 170550 246200 170555 246256
rect 98686 246198 170555 246200
rect 67449 246195 67515 246198
rect 98686 245956 98746 246198
rect 101397 246195 101463 246198
rect 170489 246195 170555 246198
rect 189901 245714 189967 245717
rect 193630 245714 193690 246500
rect 253933 246394 253999 246397
rect 253460 246392 253999 246394
rect 253460 246336 253938 246392
rect 253994 246336 253999 246392
rect 253460 246334 253999 246336
rect 253933 246331 253999 246334
rect 256509 246258 256575 246261
rect 261201 246258 261267 246261
rect 266302 246258 266308 246260
rect 256509 246256 266308 246258
rect 256509 246200 256514 246256
rect 256570 246200 261206 246256
rect 261262 246200 266308 246256
rect 256509 246198 266308 246200
rect 256509 246195 256575 246198
rect 261201 246195 261267 246198
rect 266302 246196 266308 246198
rect 266372 246196 266378 246260
rect 252878 245853 252938 245956
rect 252878 245848 252987 245853
rect 252878 245792 252926 245848
rect 252982 245792 252987 245848
rect 252878 245790 252987 245792
rect 252921 245787 252987 245790
rect 189901 245712 193690 245714
rect 189901 245656 189906 245712
rect 189962 245656 193690 245712
rect 189901 245654 193690 245656
rect 189901 245651 189967 245654
rect 254025 245578 254091 245581
rect 276238 245578 276244 245580
rect 253460 245576 276244 245578
rect 253460 245520 254030 245576
rect 254086 245520 276244 245576
rect 253460 245518 276244 245520
rect 254025 245515 254091 245518
rect 276238 245516 276244 245518
rect 276308 245516 276314 245580
rect 582373 245578 582439 245581
rect 583520 245578 584960 245668
rect 582373 245576 584960 245578
rect 582373 245520 582378 245576
rect 582434 245520 584960 245576
rect 582373 245518 584960 245520
rect 582373 245515 582439 245518
rect 66805 245442 66871 245445
rect 66805 245440 68908 245442
rect 66805 245384 66810 245440
rect 66866 245384 68908 245440
rect 583520 245428 584960 245518
rect 66805 245382 68908 245384
rect 66805 245379 66871 245382
rect 100937 245170 101003 245173
rect 98716 245168 101003 245170
rect 98716 245112 100942 245168
rect 100998 245112 101003 245168
rect 98716 245110 101003 245112
rect 100937 245107 101003 245110
rect 104433 244898 104499 244901
rect 152549 244898 152615 244901
rect 104433 244896 152615 244898
rect 104433 244840 104438 244896
rect 104494 244840 152554 244896
rect 152610 244840 152615 244896
rect 104433 244838 152615 244840
rect 104433 244835 104499 244838
rect 152549 244835 152615 244838
rect 155309 244898 155375 244901
rect 181621 244898 181687 244901
rect 155309 244896 181687 244898
rect 155309 244840 155314 244896
rect 155370 244840 181626 244896
rect 181682 244840 181687 244896
rect 155309 244838 181687 244840
rect 155309 244835 155375 244838
rect 181621 244835 181687 244838
rect 69430 244356 69490 244596
rect 184054 244564 184060 244628
rect 184124 244626 184130 244628
rect 193630 244626 193690 245412
rect 252878 245037 252938 245140
rect 252829 245032 252938 245037
rect 252829 244976 252834 245032
rect 252890 244976 252938 245032
rect 252829 244974 252938 244976
rect 252829 244971 252895 244974
rect 255313 244762 255379 244765
rect 253460 244760 255379 244762
rect 253460 244704 255318 244760
rect 255374 244704 255379 244760
rect 253460 244702 255379 244704
rect 255313 244699 255379 244702
rect 184124 244566 193690 244626
rect 184124 244564 184130 244566
rect 184238 244428 184244 244492
rect 184308 244490 184314 244492
rect 252829 244490 252895 244493
rect 184308 244430 193690 244490
rect 184308 244428 184314 244430
rect 69422 244292 69428 244356
rect 69492 244292 69498 244356
rect 101029 244354 101095 244357
rect 98716 244352 101095 244354
rect 98716 244296 101034 244352
rect 101090 244296 101095 244352
rect 193630 244324 193690 244430
rect 252829 244488 255882 244490
rect 252829 244432 252834 244488
rect 252890 244432 255882 244488
rect 252829 244430 255882 244432
rect 252829 244427 252895 244430
rect 98716 244294 101095 244296
rect 101029 244291 101095 244294
rect 255681 244218 255747 244221
rect 253460 244216 255747 244218
rect 253460 244160 255686 244216
rect 255742 244160 255747 244216
rect 253460 244158 255747 244160
rect 255822 244218 255882 244430
rect 267958 244218 267964 244220
rect 255822 244158 267964 244218
rect 255681 244155 255747 244158
rect 267958 244156 267964 244158
rect 268028 244156 268034 244220
rect 66897 243810 66963 243813
rect 255773 243810 255839 243813
rect 66897 243808 68908 243810
rect 66897 243752 66902 243808
rect 66958 243752 68908 243808
rect 66897 243750 68908 243752
rect 253460 243808 255839 243810
rect 253460 243752 255778 243808
rect 255834 243752 255839 243808
rect 253460 243750 255839 243752
rect 66897 243747 66963 243750
rect 255773 243747 255839 243750
rect 253606 243612 253612 243676
rect 253676 243674 253682 243676
rect 260925 243674 260991 243677
rect 253676 243672 260991 243674
rect 253676 243616 260930 243672
rect 260986 243616 260991 243672
rect 253676 243614 260991 243616
rect 253676 243612 253682 243614
rect 260925 243611 260991 243614
rect 102726 243538 102732 243540
rect 98716 243478 102732 243538
rect 102726 243476 102732 243478
rect 102796 243476 102802 243540
rect 255497 243402 255563 243405
rect 253460 243400 255563 243402
rect 253460 243344 255502 243400
rect 255558 243344 255563 243400
rect 253460 243342 255563 243344
rect 255497 243339 255563 243342
rect 66713 242994 66779 242997
rect 189993 242994 190059 242997
rect 193630 242994 193690 243236
rect 253933 242994 253999 242997
rect 66713 242992 68908 242994
rect 66713 242936 66718 242992
rect 66774 242936 68908 242992
rect 66713 242934 68908 242936
rect 189993 242992 193690 242994
rect 189993 242936 189998 242992
rect 190054 242936 193690 242992
rect 189993 242934 193690 242936
rect 253460 242992 253999 242994
rect 253460 242936 253938 242992
rect 253994 242936 253999 242992
rect 253460 242934 253999 242936
rect 66713 242931 66779 242934
rect 189993 242931 190059 242934
rect 253933 242931 253999 242934
rect 193438 242796 193444 242860
rect 193508 242858 193514 242860
rect 193673 242858 193739 242861
rect 193508 242856 193739 242858
rect 193508 242800 193678 242856
rect 193734 242800 193739 242856
rect 193508 242798 193739 242800
rect 193508 242796 193514 242798
rect 193673 242795 193739 242798
rect 102225 242722 102291 242725
rect 98716 242720 102291 242722
rect 98716 242664 102230 242720
rect 102286 242664 102291 242720
rect 98716 242662 102291 242664
rect 102225 242659 102291 242662
rect 98729 242586 98795 242589
rect 112437 242586 112503 242589
rect 98729 242584 112503 242586
rect 98729 242528 98734 242584
rect 98790 242528 112442 242584
rect 112498 242528 112503 242584
rect 98729 242526 112503 242528
rect 98729 242523 98795 242526
rect 112437 242523 112503 242526
rect 252878 242453 252938 242556
rect 99097 242450 99163 242453
rect 129181 242450 129247 242453
rect 99097 242448 129247 242450
rect 99097 242392 99102 242448
rect 99158 242392 129186 242448
rect 129242 242392 129247 242448
rect 99097 242390 129247 242392
rect 99097 242387 99163 242390
rect 129181 242387 129247 242390
rect 252829 242448 252938 242453
rect 252829 242392 252834 242448
rect 252890 242392 252938 242448
rect 252829 242390 252938 242392
rect 255497 242450 255563 242453
rect 268285 242450 268351 242453
rect 255497 242448 268351 242450
rect 255497 242392 255502 242448
rect 255558 242392 268290 242448
rect 268346 242392 268351 242448
rect 255497 242390 268351 242392
rect 252829 242387 252895 242390
rect 255497 242387 255563 242390
rect 268285 242387 268351 242390
rect 261109 242314 261175 242317
rect 281574 242314 281580 242316
rect 261109 242312 281580 242314
rect 261109 242256 261114 242312
rect 261170 242256 281580 242312
rect 261109 242254 281580 242256
rect 261109 242251 261175 242254
rect 281574 242252 281580 242254
rect 281644 242252 281650 242316
rect 66805 242178 66871 242181
rect 255497 242178 255563 242181
rect 284385 242178 284451 242181
rect 66805 242176 68908 242178
rect 66805 242120 66810 242176
rect 66866 242120 68908 242176
rect 253460 242176 255563 242178
rect 66805 242118 68908 242120
rect 66805 242115 66871 242118
rect 104341 241906 104407 241909
rect 98716 241904 104407 241906
rect 98716 241848 104346 241904
rect 104402 241848 104407 241904
rect 98716 241846 104407 241848
rect 104341 241843 104407 241846
rect 70945 241772 71011 241773
rect 70894 241708 70900 241772
rect 70964 241770 71011 241772
rect 83825 241770 83891 241773
rect 86585 241772 86651 241773
rect 84510 241770 84516 241772
rect 70964 241768 71056 241770
rect 71006 241712 71056 241768
rect 70964 241710 71056 241712
rect 83825 241768 84516 241770
rect 83825 241712 83830 241768
rect 83886 241712 84516 241768
rect 83825 241710 84516 241712
rect 70964 241708 71011 241710
rect 70945 241707 71011 241708
rect 83825 241707 83891 241710
rect 84510 241708 84516 241710
rect 84580 241708 84586 241772
rect 86534 241708 86540 241772
rect 86604 241770 86651 241772
rect 90357 241770 90423 241773
rect 91553 241772 91619 241773
rect 90950 241770 90956 241772
rect 86604 241768 86696 241770
rect 86646 241712 86696 241768
rect 86604 241710 86696 241712
rect 90357 241768 90956 241770
rect 90357 241712 90362 241768
rect 90418 241712 90956 241768
rect 90357 241710 90956 241712
rect 86604 241708 86651 241710
rect 86585 241707 86651 241708
rect 90357 241707 90423 241710
rect 90950 241708 90956 241710
rect 91020 241708 91026 241772
rect 91502 241708 91508 241772
rect 91572 241770 91619 241772
rect 95877 241770 95943 241773
rect 98729 241770 98795 241773
rect 91572 241768 91664 241770
rect 91614 241712 91664 241768
rect 91572 241710 91664 241712
rect 95877 241768 98795 241770
rect 95877 241712 95882 241768
rect 95938 241712 98734 241768
rect 98790 241712 98795 241768
rect 95877 241710 98795 241712
rect 91572 241708 91619 241710
rect 91553 241707 91619 241708
rect 95877 241707 95943 241710
rect 98729 241707 98795 241710
rect 85849 241634 85915 241637
rect 88006 241634 88012 241636
rect 85849 241632 88012 241634
rect 85849 241576 85854 241632
rect 85910 241576 88012 241632
rect 85849 241574 88012 241576
rect 85849 241571 85915 241574
rect 88006 241572 88012 241574
rect 88076 241572 88082 241636
rect 186957 241634 187023 241637
rect 193630 241634 193690 242148
rect 253460 242120 255502 242176
rect 255558 242120 255563 242176
rect 253460 242118 255563 242120
rect 255497 242115 255563 242118
rect 258030 242176 284451 242178
rect 258030 242120 284390 242176
rect 284446 242120 284451 242176
rect 258030 242118 284451 242120
rect 193765 242042 193831 242045
rect 194501 242042 194567 242045
rect 195789 242044 195855 242045
rect 248505 242044 248571 242045
rect 195789 242042 195836 242044
rect 193765 242040 194567 242042
rect 193765 241984 193770 242040
rect 193826 241984 194506 242040
rect 194562 241984 194567 242040
rect 193765 241982 194567 241984
rect 195744 242040 195836 242042
rect 195744 241984 195794 242040
rect 195744 241982 195836 241984
rect 193765 241979 193831 241982
rect 194501 241979 194567 241982
rect 195789 241980 195836 241982
rect 195900 241980 195906 242044
rect 248454 241980 248460 242044
rect 248524 242042 248571 242044
rect 258030 242042 258090 242118
rect 284385 242115 284451 242118
rect 248524 242040 248616 242042
rect 248566 241984 248616 242040
rect 248524 241982 248616 241984
rect 253430 241982 258090 242042
rect 248524 241980 248571 241982
rect 195789 241979 195855 241980
rect 248505 241979 248571 241980
rect 253430 241740 253490 241982
rect 186957 241632 193690 241634
rect 186957 241576 186962 241632
rect 187018 241576 193690 241632
rect 186957 241574 193690 241576
rect 186957 241571 187023 241574
rect 67950 241436 67956 241500
rect 68020 241498 68026 241500
rect 68921 241498 68987 241501
rect 68020 241496 68987 241498
rect 68020 241440 68926 241496
rect 68982 241440 68987 241496
rect 68020 241438 68987 241440
rect 68020 241436 68026 241438
rect 68921 241435 68987 241438
rect 92335 241498 92401 241501
rect 255773 241498 255839 241501
rect 277158 241498 277164 241500
rect 92335 241496 277164 241498
rect 92335 241440 92340 241496
rect 92396 241440 255778 241496
rect 255834 241440 277164 241496
rect 92335 241438 277164 241440
rect 92335 241435 92401 241438
rect 255773 241435 255839 241438
rect 277158 241436 277164 241438
rect 277228 241436 277234 241500
rect 14457 241362 14523 241365
rect 93117 241362 93183 241365
rect 93439 241362 93505 241365
rect 14457 241360 93505 241362
rect 14457 241304 14462 241360
rect 14518 241304 93122 241360
rect 93178 241304 93444 241360
rect 93500 241304 93505 241360
rect 14457 241302 93505 241304
rect 14457 241299 14523 241302
rect 93117 241299 93183 241302
rect 93439 241299 93505 241302
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 68645 240818 68711 240821
rect 77937 240818 78003 240821
rect 68645 240816 78003 240818
rect 68645 240760 68650 240816
rect 68706 240760 77942 240816
rect 77998 240760 78003 240816
rect 68645 240758 78003 240760
rect 68645 240755 68711 240758
rect 77937 240755 78003 240758
rect 173709 240818 173775 240821
rect 182265 240818 182331 240821
rect 173709 240816 182331 240818
rect 173709 240760 173714 240816
rect 173770 240760 182270 240816
rect 182326 240760 182331 240816
rect 173709 240758 182331 240760
rect 173709 240755 173775 240758
rect 182265 240755 182331 240758
rect 184197 240818 184263 240821
rect 217961 240818 218027 240821
rect 184197 240816 218027 240818
rect 184197 240760 184202 240816
rect 184258 240760 217966 240816
rect 218022 240760 218027 240816
rect 184197 240758 218027 240760
rect 184197 240755 184263 240758
rect 217961 240755 218027 240758
rect 218697 240818 218763 240821
rect 256877 240818 256943 240821
rect 218697 240816 256943 240818
rect 218697 240760 218702 240816
rect 218758 240760 256882 240816
rect 256938 240760 256943 240816
rect 218697 240758 256943 240760
rect 218697 240755 218763 240758
rect 256877 240755 256943 240758
rect 257337 240274 257403 240277
rect 258390 240274 258396 240276
rect 257337 240272 258396 240274
rect 257337 240216 257342 240272
rect 257398 240216 258396 240272
rect 257337 240214 258396 240216
rect 257337 240211 257403 240214
rect 258390 240212 258396 240214
rect 258460 240212 258466 240276
rect 277158 240212 277164 240276
rect 277228 240274 277234 240276
rect 277485 240274 277551 240277
rect 277228 240272 277551 240274
rect 277228 240216 277490 240272
rect 277546 240216 277551 240272
rect 277228 240214 277551 240216
rect 277228 240212 277234 240214
rect 277485 240211 277551 240214
rect 68553 240138 68619 240141
rect 71405 240140 71471 240141
rect 68870 240138 68876 240140
rect 68553 240136 68876 240138
rect 68553 240080 68558 240136
rect 68614 240080 68876 240136
rect 68553 240078 68876 240080
rect 68553 240075 68619 240078
rect 68870 240076 68876 240078
rect 68940 240076 68946 240140
rect 71405 240136 71452 240140
rect 71516 240138 71522 240140
rect 71865 240138 71931 240141
rect 72969 240140 73035 240141
rect 72366 240138 72372 240140
rect 71405 240080 71410 240136
rect 71405 240076 71452 240080
rect 71516 240078 71562 240138
rect 71865 240136 72372 240138
rect 71865 240080 71870 240136
rect 71926 240080 72372 240136
rect 71865 240078 72372 240080
rect 71516 240076 71522 240078
rect 71405 240075 71471 240076
rect 71865 240075 71931 240078
rect 72366 240076 72372 240078
rect 72436 240076 72442 240140
rect 72918 240138 72924 240140
rect 72878 240078 72924 240138
rect 72988 240136 73035 240140
rect 73030 240080 73035 240136
rect 72918 240076 72924 240078
rect 72988 240076 73035 240080
rect 73286 240076 73292 240140
rect 73356 240138 73362 240140
rect 74349 240138 74415 240141
rect 90909 240140 90975 240141
rect 90909 240138 90956 240140
rect 73356 240136 74415 240138
rect 73356 240080 74354 240136
rect 74410 240080 74415 240136
rect 73356 240078 74415 240080
rect 90864 240136 90956 240138
rect 90864 240080 90914 240136
rect 90864 240078 90956 240080
rect 73356 240076 73362 240078
rect 72969 240075 73035 240076
rect 74349 240075 74415 240078
rect 90909 240076 90956 240078
rect 91020 240076 91026 240140
rect 97533 240138 97599 240141
rect 97758 240138 97764 240140
rect 97533 240136 97764 240138
rect 97533 240080 97538 240136
rect 97594 240080 97764 240136
rect 97533 240078 97764 240080
rect 90909 240075 90975 240076
rect 97533 240075 97599 240078
rect 97758 240076 97764 240078
rect 97828 240076 97834 240140
rect 168373 240138 168439 240141
rect 169109 240138 169175 240141
rect 247033 240138 247099 240141
rect 168373 240136 247099 240138
rect 168373 240080 168378 240136
rect 168434 240080 169114 240136
rect 169170 240080 247038 240136
rect 247094 240080 247099 240136
rect 168373 240078 247099 240080
rect 168373 240075 168439 240078
rect 169109 240075 169175 240078
rect 247033 240075 247099 240078
rect 251909 240138 251975 240141
rect 253933 240138 253999 240141
rect 251909 240136 253999 240138
rect 251909 240080 251914 240136
rect 251970 240080 253938 240136
rect 253994 240080 253999 240136
rect 251909 240078 253999 240080
rect 251909 240075 251975 240078
rect 253933 240075 253999 240078
rect 72233 240002 72299 240005
rect 72734 240002 72740 240004
rect 72233 240000 72740 240002
rect 72233 239944 72238 240000
rect 72294 239944 72740 240000
rect 72233 239942 72740 239944
rect 72233 239939 72299 239942
rect 72734 239940 72740 239942
rect 72804 239940 72810 240004
rect 82261 240002 82327 240005
rect 98269 240002 98335 240005
rect 82261 240000 98335 240002
rect 82261 239944 82266 240000
rect 82322 239944 98274 240000
rect 98330 239944 98335 240000
rect 82261 239942 98335 239944
rect 82261 239939 82327 239942
rect 98269 239939 98335 239942
rect 98729 240002 98795 240005
rect 103421 240002 103487 240005
rect 170949 240002 171015 240005
rect 180333 240002 180399 240005
rect 252277 240002 252343 240005
rect 98729 240000 171150 240002
rect 98729 239944 98734 240000
rect 98790 239944 103426 240000
rect 103482 239944 170954 240000
rect 171010 239944 171150 240000
rect 98729 239942 171150 239944
rect 98729 239939 98795 239942
rect 103421 239939 103487 239942
rect 170949 239939 171015 239942
rect 72550 239804 72556 239868
rect 72620 239866 72626 239868
rect 73521 239866 73587 239869
rect 72620 239864 73587 239866
rect 72620 239808 73526 239864
rect 73582 239808 73587 239864
rect 72620 239806 73587 239808
rect 72620 239804 72626 239806
rect 73521 239803 73587 239806
rect 87597 239866 87663 239869
rect 88006 239866 88012 239868
rect 87597 239864 88012 239866
rect 87597 239808 87602 239864
rect 87658 239808 88012 239864
rect 87597 239806 88012 239808
rect 87597 239803 87663 239806
rect 88006 239804 88012 239806
rect 88076 239804 88082 239868
rect 171090 239866 171150 239942
rect 180333 240000 252343 240002
rect 180333 239944 180338 240000
rect 180394 239944 252282 240000
rect 252338 239944 252343 240000
rect 180333 239942 252343 239944
rect 180333 239939 180399 239942
rect 252277 239939 252343 239942
rect 171090 239806 180810 239866
rect 180750 239730 180810 239806
rect 192334 239804 192340 239868
rect 192404 239866 192410 239868
rect 193121 239866 193187 239869
rect 192404 239864 193187 239866
rect 192404 239808 193126 239864
rect 193182 239808 193187 239864
rect 192404 239806 193187 239808
rect 192404 239804 192410 239806
rect 193121 239803 193187 239806
rect 195237 239730 195303 239733
rect 180750 239728 195303 239730
rect 180750 239672 195242 239728
rect 195298 239672 195303 239728
rect 180750 239670 195303 239672
rect 195237 239667 195303 239670
rect 56501 239458 56567 239461
rect 72877 239458 72943 239461
rect 56501 239456 72943 239458
rect 56501 239400 56506 239456
rect 56562 239400 72882 239456
rect 72938 239400 72943 239456
rect 56501 239398 72943 239400
rect 56501 239395 56567 239398
rect 72877 239395 72943 239398
rect 86861 239458 86927 239461
rect 96654 239458 96660 239460
rect 86861 239456 96660 239458
rect 86861 239400 86866 239456
rect 86922 239400 96660 239456
rect 86861 239398 96660 239400
rect 86861 239395 86927 239398
rect 96654 239396 96660 239398
rect 96724 239396 96730 239460
rect 246297 239458 246363 239461
rect 259678 239458 259684 239460
rect 246297 239456 259684 239458
rect 246297 239400 246302 239456
rect 246358 239400 259684 239456
rect 246297 239398 259684 239400
rect 246297 239395 246363 239398
rect 259678 239396 259684 239398
rect 259748 239396 259754 239460
rect 72785 239322 72851 239325
rect 168373 239322 168439 239325
rect 72785 239320 168439 239322
rect 72785 239264 72790 239320
rect 72846 239264 168378 239320
rect 168434 239264 168439 239320
rect 72785 239262 168439 239264
rect 72785 239259 72851 239262
rect 168373 239259 168439 239262
rect 70301 239186 70367 239189
rect 76557 239186 76623 239189
rect 70301 239184 76623 239186
rect 70301 239128 70306 239184
rect 70362 239128 76562 239184
rect 76618 239128 76623 239184
rect 70301 239126 76623 239128
rect 70301 239123 70367 239126
rect 76557 239123 76623 239126
rect 84101 238778 84167 238781
rect 84510 238778 84516 238780
rect 84101 238776 84516 238778
rect 84101 238720 84106 238776
rect 84162 238720 84516 238776
rect 84101 238718 84516 238720
rect 84101 238715 84167 238718
rect 84510 238716 84516 238718
rect 84580 238716 84586 238780
rect 96521 238778 96587 238781
rect 96654 238778 96660 238780
rect 96521 238776 96660 238778
rect 96521 238720 96526 238776
rect 96582 238720 96660 238776
rect 96521 238718 96660 238720
rect 96521 238715 96587 238718
rect 96654 238716 96660 238718
rect 96724 238716 96730 238780
rect 160921 238642 160987 238645
rect 265249 238642 265315 238645
rect 160921 238640 265315 238642
rect 160921 238584 160926 238640
rect 160982 238584 265254 238640
rect 265310 238584 265315 238640
rect 160921 238582 265315 238584
rect 160921 238579 160987 238582
rect 265249 238579 265315 238582
rect 75913 238506 75979 238509
rect 110597 238506 110663 238509
rect 75913 238504 110663 238506
rect 75913 238448 75918 238504
rect 75974 238448 110602 238504
rect 110658 238448 110663 238504
rect 75913 238446 110663 238448
rect 75913 238443 75979 238446
rect 110597 238443 110663 238446
rect 57513 238370 57579 238373
rect 77569 238370 77635 238373
rect 57513 238368 77635 238370
rect 57513 238312 57518 238368
rect 57574 238312 77574 238368
rect 77630 238312 77635 238368
rect 57513 238310 77635 238312
rect 57513 238307 57579 238310
rect 77569 238307 77635 238310
rect 67357 238234 67423 238237
rect 113817 238234 113883 238237
rect 67357 238232 113883 238234
rect 67357 238176 67362 238232
rect 67418 238176 113822 238232
rect 113878 238176 113883 238232
rect 67357 238174 113883 238176
rect 67357 238171 67423 238174
rect 113817 238171 113883 238174
rect 103421 238098 103487 238101
rect 187141 238098 187207 238101
rect 103421 238096 187207 238098
rect 103421 238040 103426 238096
rect 103482 238040 187146 238096
rect 187202 238040 187207 238096
rect 103421 238038 187207 238040
rect 103421 238035 103487 238038
rect 187141 238035 187207 238038
rect 191741 238098 191807 238101
rect 200614 238098 200620 238100
rect 191741 238096 200620 238098
rect 191741 238040 191746 238096
rect 191802 238040 200620 238096
rect 191741 238038 200620 238040
rect 191741 238035 191807 238038
rect 200614 238036 200620 238038
rect 200684 238036 200690 238100
rect 180057 237962 180123 237965
rect 197353 237962 197419 237965
rect 258349 237962 258415 237965
rect 180057 237960 258415 237962
rect 180057 237904 180062 237960
rect 180118 237904 197358 237960
rect 197414 237904 258354 237960
rect 258410 237904 258415 237960
rect 180057 237902 258415 237904
rect 180057 237899 180123 237902
rect 197353 237899 197419 237902
rect 258349 237899 258415 237902
rect 93710 237356 93716 237420
rect 93780 237418 93786 237420
rect 93945 237418 94011 237421
rect 93780 237416 94011 237418
rect 93780 237360 93950 237416
rect 94006 237360 94011 237416
rect 93780 237358 94011 237360
rect 93780 237356 93786 237358
rect 93945 237355 94011 237358
rect 160737 237418 160803 237421
rect 160921 237418 160987 237421
rect 160737 237416 160987 237418
rect 160737 237360 160742 237416
rect 160798 237360 160926 237416
rect 160982 237360 160987 237416
rect 160737 237358 160987 237360
rect 160737 237355 160803 237358
rect 160921 237355 160987 237358
rect 175181 237282 175247 237285
rect 262397 237282 262463 237285
rect 175181 237280 262463 237282
rect 175181 237224 175186 237280
rect 175242 237224 262402 237280
rect 262458 237224 262463 237280
rect 175181 237222 262463 237224
rect 175181 237219 175247 237222
rect 262397 237219 262463 237222
rect 94129 236738 94195 236741
rect 116577 236738 116643 236741
rect 122097 236738 122163 236741
rect 94129 236736 122163 236738
rect 94129 236680 94134 236736
rect 94190 236680 116582 236736
rect 116638 236680 122102 236736
rect 122158 236680 122163 236736
rect 94129 236678 122163 236680
rect 94129 236675 94195 236678
rect 116577 236675 116643 236678
rect 122097 236675 122163 236678
rect 15101 236602 15167 236605
rect 189993 236602 190059 236605
rect 15101 236600 190059 236602
rect 15101 236544 15106 236600
rect 15162 236544 189998 236600
rect 190054 236544 190059 236600
rect 15101 236542 190059 236544
rect 15101 236539 15167 236542
rect 189993 236539 190059 236542
rect 192569 236602 192635 236605
rect 208342 236602 208348 236604
rect 192569 236600 208348 236602
rect 192569 236544 192574 236600
rect 192630 236544 208348 236600
rect 192569 236542 208348 236544
rect 192569 236539 192635 236542
rect 208342 236540 208348 236542
rect 208412 236540 208418 236604
rect 222101 236602 222167 236605
rect 263869 236602 263935 236605
rect 222101 236600 263935 236602
rect 222101 236544 222106 236600
rect 222162 236544 263874 236600
rect 263930 236544 263935 236600
rect 222101 236542 263935 236544
rect 222101 236539 222167 236542
rect 263869 236539 263935 236542
rect 69606 235860 69612 235924
rect 69676 235922 69682 235924
rect 116761 235922 116827 235925
rect 69676 235920 116827 235922
rect 69676 235864 116766 235920
rect 116822 235864 116827 235920
rect 69676 235862 116827 235864
rect 69676 235860 69682 235862
rect 116761 235859 116827 235862
rect 159541 235922 159607 235925
rect 160001 235922 160067 235925
rect 258390 235922 258396 235924
rect 159541 235920 258396 235922
rect 159541 235864 159546 235920
rect 159602 235864 160006 235920
rect 160062 235864 258396 235920
rect 159541 235862 258396 235864
rect 159541 235859 159607 235862
rect 160001 235859 160067 235862
rect 258390 235860 258396 235862
rect 258460 235860 258466 235924
rect 181621 235378 181687 235381
rect 181621 235376 219450 235378
rect 181621 235320 181626 235376
rect 181682 235320 219450 235376
rect 181621 235318 219450 235320
rect 181621 235315 181687 235318
rect 28901 235242 28967 235245
rect 189901 235242 189967 235245
rect 28901 235240 189967 235242
rect 28901 235184 28906 235240
rect 28962 235184 189906 235240
rect 189962 235184 189967 235240
rect 28901 235182 189967 235184
rect 28901 235179 28967 235182
rect 189901 235179 189967 235182
rect 193806 235180 193812 235244
rect 193876 235242 193882 235244
rect 218145 235242 218211 235245
rect 193876 235240 218211 235242
rect 193876 235184 218150 235240
rect 218206 235184 218211 235240
rect 193876 235182 218211 235184
rect 219390 235242 219450 235318
rect 219525 235242 219591 235245
rect 248454 235242 248460 235244
rect 219390 235240 248460 235242
rect 219390 235184 219530 235240
rect 219586 235184 248460 235240
rect 219390 235182 248460 235184
rect 193876 235180 193882 235182
rect 218145 235179 218211 235182
rect 219525 235179 219591 235182
rect 248454 235180 248460 235182
rect 248524 235180 248530 235244
rect 84285 234562 84351 234565
rect 181529 234562 181595 234565
rect 84285 234560 181595 234562
rect 84285 234504 84290 234560
rect 84346 234504 181534 234560
rect 181590 234504 181595 234560
rect 84285 234502 181595 234504
rect 84285 234499 84351 234502
rect 181529 234499 181595 234502
rect 96705 234018 96771 234021
rect 97574 234018 97580 234020
rect 96705 234016 97580 234018
rect 96705 233960 96710 234016
rect 96766 233960 97580 234016
rect 96705 233958 97580 233960
rect 96705 233955 96771 233958
rect 97574 233956 97580 233958
rect 97644 233956 97650 234020
rect 97809 234018 97875 234021
rect 99966 234018 99972 234020
rect 97809 234016 99972 234018
rect 97809 233960 97814 234016
rect 97870 233960 99972 234016
rect 97809 233958 99972 233960
rect 97809 233955 97875 233958
rect 99966 233956 99972 233958
rect 100036 233956 100042 234020
rect 171133 234018 171199 234021
rect 227713 234018 227779 234021
rect 261109 234018 261175 234021
rect 171133 234016 261175 234018
rect 171133 233960 171138 234016
rect 171194 233960 227718 234016
rect 227774 233960 261114 234016
rect 261170 233960 261175 234016
rect 171133 233958 261175 233960
rect 171133 233955 171199 233958
rect 227713 233955 227779 233958
rect 261109 233955 261175 233958
rect 39941 233882 40007 233885
rect 188337 233882 188403 233885
rect 39941 233880 188403 233882
rect 39941 233824 39946 233880
rect 40002 233824 188342 233880
rect 188398 233824 188403 233880
rect 39941 233822 188403 233824
rect 39941 233819 40007 233822
rect 188337 233819 188403 233822
rect 192702 233820 192708 233884
rect 192772 233882 192778 233884
rect 202873 233882 202939 233885
rect 192772 233880 202939 233882
rect 192772 233824 202878 233880
rect 202934 233824 202939 233880
rect 192772 233822 202939 233824
rect 192772 233820 192778 233822
rect 202873 233819 202939 233822
rect 207054 233820 207060 233884
rect 207124 233882 207130 233884
rect 269389 233882 269455 233885
rect 207124 233880 269455 233882
rect 207124 233824 269394 233880
rect 269450 233824 269455 233880
rect 207124 233822 269455 233824
rect 207124 233820 207130 233822
rect 269389 233819 269455 233822
rect 60457 233202 60523 233205
rect 156689 233202 156755 233205
rect 60457 233200 156755 233202
rect 60457 233144 60462 233200
rect 60518 233144 156694 233200
rect 156750 233144 156755 233200
rect 60457 233142 156755 233144
rect 60457 233139 60523 233142
rect 156689 233139 156755 233142
rect 180701 233202 180767 233205
rect 215293 233202 215359 233205
rect 180701 233200 215359 233202
rect 180701 233144 180706 233200
rect 180762 233144 215298 233200
rect 215354 233144 215359 233200
rect 180701 233142 215359 233144
rect 180701 233139 180767 233142
rect 215293 233139 215359 233142
rect 189809 233066 189875 233069
rect 207054 233066 207060 233068
rect 189809 233064 207060 233066
rect 189809 233008 189814 233064
rect 189870 233008 207060 233064
rect 189809 233006 207060 233008
rect 189809 233003 189875 233006
rect 207054 233004 207060 233006
rect 207124 233004 207130 233068
rect 247677 232658 247743 232661
rect 270769 232658 270835 232661
rect 247677 232656 270835 232658
rect 247677 232600 247682 232656
rect 247738 232600 270774 232656
rect 270830 232600 270835 232656
rect 247677 232598 270835 232600
rect 247677 232595 247743 232598
rect 270769 232595 270835 232598
rect 92473 232522 92539 232525
rect 111241 232522 111307 232525
rect 92473 232520 111307 232522
rect 92473 232464 92478 232520
rect 92534 232464 111246 232520
rect 111302 232464 111307 232520
rect 92473 232462 111307 232464
rect 92473 232459 92539 232462
rect 111241 232459 111307 232462
rect 215201 232522 215267 232525
rect 255405 232522 255471 232525
rect 215201 232520 255471 232522
rect 215201 232464 215206 232520
rect 215262 232464 255410 232520
rect 255466 232464 255471 232520
rect 215201 232462 255471 232464
rect 215201 232459 215267 232462
rect 255405 232459 255471 232462
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 191230 231780 191236 231844
rect 191300 231842 191306 231844
rect 222837 231842 222903 231845
rect 223481 231842 223547 231845
rect 191300 231840 223547 231842
rect 191300 231784 222842 231840
rect 222898 231784 223486 231840
rect 223542 231784 223547 231840
rect 191300 231782 223547 231784
rect 191300 231780 191306 231782
rect 222837 231779 222903 231782
rect 223481 231779 223547 231782
rect 68921 231162 68987 231165
rect 128353 231162 128419 231165
rect 68921 231160 128419 231162
rect 68921 231104 68926 231160
rect 68982 231104 128358 231160
rect 128414 231104 128419 231160
rect 68921 231102 128419 231104
rect 68921 231099 68987 231102
rect 128353 231099 128419 231102
rect 186998 231100 187004 231164
rect 187068 231162 187074 231164
rect 276422 231162 276428 231164
rect 187068 231102 276428 231162
rect 187068 231100 187074 231102
rect 276422 231100 276428 231102
rect 276492 231100 276498 231164
rect 178953 230482 179019 230485
rect 262489 230482 262555 230485
rect 178953 230480 262555 230482
rect 178953 230424 178958 230480
rect 179014 230424 262494 230480
rect 262550 230424 262555 230480
rect 178953 230422 262555 230424
rect 178953 230419 179019 230422
rect 262489 230419 262555 230422
rect 152549 229802 152615 229805
rect 180057 229802 180123 229805
rect 152549 229800 180123 229802
rect 152549 229744 152554 229800
rect 152610 229744 180062 229800
rect 180118 229744 180123 229800
rect 152549 229742 180123 229744
rect 152549 229739 152615 229742
rect 180057 229739 180123 229742
rect 169569 228986 169635 228989
rect 263542 228986 263548 228988
rect 169569 228984 263548 228986
rect 169569 228928 169574 228984
rect 169630 228928 263548 228984
rect 169569 228926 263548 228928
rect 169569 228923 169635 228926
rect 263542 228924 263548 228926
rect 263612 228924 263618 228988
rect 152549 228306 152615 228309
rect 162209 228306 162275 228309
rect 152549 228304 162275 228306
rect 152549 228248 152554 228304
rect 152610 228248 162214 228304
rect 162270 228248 162275 228304
rect 152549 228246 162275 228248
rect 152549 228243 152615 228246
rect 162209 228243 162275 228246
rect -960 227884 480 228124
rect 69054 227564 69060 227628
rect 69124 227626 69130 227628
rect 144269 227626 144335 227629
rect 69124 227624 144335 227626
rect 69124 227568 144274 227624
rect 144330 227568 144335 227624
rect 69124 227566 144335 227568
rect 69124 227564 69130 227566
rect 144269 227563 144335 227566
rect 213821 227626 213887 227629
rect 267774 227626 267780 227628
rect 213821 227624 267780 227626
rect 213821 227568 213826 227624
rect 213882 227568 267780 227624
rect 213821 227566 267780 227568
rect 213821 227563 213887 227566
rect 267774 227564 267780 227566
rect 267844 227564 267850 227628
rect 90817 227082 90883 227085
rect 93894 227082 93900 227084
rect 90817 227080 93900 227082
rect 90817 227024 90822 227080
rect 90878 227024 93900 227080
rect 90817 227022 93900 227024
rect 90817 227019 90883 227022
rect 93894 227020 93900 227022
rect 93964 227020 93970 227084
rect 55121 226946 55187 226949
rect 69054 226946 69060 226948
rect 55121 226944 69060 226946
rect 55121 226888 55126 226944
rect 55182 226888 69060 226944
rect 55121 226886 69060 226888
rect 55121 226883 55187 226886
rect 69054 226884 69060 226886
rect 69124 226884 69130 226948
rect 131849 226946 131915 226949
rect 214557 226946 214623 226949
rect 131849 226944 214623 226946
rect 131849 226888 131854 226944
rect 131910 226888 214562 226944
rect 214618 226888 214623 226944
rect 131849 226886 214623 226888
rect 131849 226883 131915 226886
rect 214557 226883 214623 226886
rect 86861 226402 86927 226405
rect 90030 226402 90036 226404
rect 86861 226400 90036 226402
rect 86861 226344 86866 226400
rect 86922 226344 90036 226400
rect 86861 226342 90036 226344
rect 86861 226339 86927 226342
rect 90030 226340 90036 226342
rect 90100 226340 90106 226404
rect 115197 226266 115263 226269
rect 246297 226266 246363 226269
rect 115197 226264 246363 226266
rect 115197 226208 115202 226264
rect 115258 226208 246302 226264
rect 246358 226208 246363 226264
rect 115197 226206 246363 226208
rect 115197 226203 115263 226206
rect 246297 226203 246363 226206
rect 104249 225586 104315 225589
rect 114553 225586 114619 225589
rect 104249 225584 114619 225586
rect 104249 225528 104254 225584
rect 104310 225528 114558 225584
rect 114614 225528 114619 225584
rect 104249 225526 114619 225528
rect 104249 225523 104315 225526
rect 114553 225523 114619 225526
rect 230381 225586 230447 225589
rect 265750 225586 265756 225588
rect 230381 225584 265756 225586
rect 230381 225528 230386 225584
rect 230442 225528 265756 225584
rect 230381 225526 265756 225528
rect 230381 225523 230447 225526
rect 265750 225524 265756 225526
rect 265820 225524 265826 225588
rect 245653 225042 245719 225045
rect 246297 225042 246363 225045
rect 245653 225040 246363 225042
rect 245653 224984 245658 225040
rect 245714 224984 246302 225040
rect 246358 224984 246363 225040
rect 245653 224982 246363 224984
rect 245653 224979 245719 224982
rect 246297 224979 246363 224982
rect 66662 224844 66668 224908
rect 66732 224906 66738 224908
rect 272149 224906 272215 224909
rect 66732 224904 272215 224906
rect 66732 224848 272154 224904
rect 272210 224848 272215 224904
rect 66732 224846 272215 224848
rect 66732 224844 66738 224846
rect 272149 224843 272215 224846
rect 102726 224708 102732 224772
rect 102796 224770 102802 224772
rect 177798 224770 177804 224772
rect 102796 224710 177804 224770
rect 102796 224708 102802 224710
rect 177798 224708 177804 224710
rect 177868 224770 177874 224772
rect 218697 224770 218763 224773
rect 177868 224768 218763 224770
rect 177868 224712 218702 224768
rect 218758 224712 218763 224768
rect 177868 224710 218763 224712
rect 177868 224708 177874 224710
rect 218697 224707 218763 224710
rect 149789 223546 149855 223549
rect 229093 223546 229159 223549
rect 230381 223546 230447 223549
rect 149789 223544 230447 223546
rect 149789 223488 149794 223544
rect 149850 223488 229098 223544
rect 229154 223488 230386 223544
rect 230442 223488 230447 223544
rect 149789 223486 230447 223488
rect 149789 223483 149855 223486
rect 229093 223483 229159 223486
rect 230381 223483 230447 223486
rect 186129 222866 186195 222869
rect 206277 222866 206343 222869
rect 186129 222864 206343 222866
rect 186129 222808 186134 222864
rect 186190 222808 206282 222864
rect 206338 222808 206343 222864
rect 186129 222806 206343 222808
rect 186129 222803 186195 222806
rect 206277 222803 206343 222806
rect 232497 222866 232563 222869
rect 258257 222866 258323 222869
rect 232497 222864 258323 222866
rect 232497 222808 232502 222864
rect 232558 222808 258262 222864
rect 258318 222808 258323 222864
rect 232497 222806 258323 222808
rect 232497 222803 232563 222806
rect 258257 222803 258323 222806
rect 214557 222186 214623 222189
rect 268377 222186 268443 222189
rect 214557 222184 268443 222186
rect 214557 222128 214562 222184
rect 214618 222128 268382 222184
rect 268438 222128 268443 222184
rect 214557 222126 268443 222128
rect 214557 222123 214623 222126
rect 268377 222123 268443 222126
rect 5441 221506 5507 221509
rect 194542 221506 194548 221508
rect 5441 221504 194548 221506
rect 5441 221448 5446 221504
rect 5502 221448 194548 221504
rect 5441 221446 194548 221448
rect 5441 221443 5507 221446
rect 194542 221444 194548 221446
rect 194612 221444 194618 221508
rect 88241 220962 88307 220965
rect 95182 220962 95188 220964
rect 88241 220960 95188 220962
rect 88241 220904 88246 220960
rect 88302 220904 95188 220960
rect 88241 220902 95188 220904
rect 88241 220899 88307 220902
rect 95182 220900 95188 220902
rect 95252 220900 95258 220964
rect 133321 220826 133387 220829
rect 227805 220826 227871 220829
rect 133321 220824 227871 220826
rect 133321 220768 133326 220824
rect 133382 220768 227810 220824
rect 227866 220768 227871 220824
rect 133321 220766 227871 220768
rect 133321 220763 133387 220766
rect 227805 220763 227871 220766
rect 74809 220146 74875 220149
rect 176009 220146 176075 220149
rect 74809 220144 176075 220146
rect 74809 220088 74814 220144
rect 74870 220088 176014 220144
rect 176070 220088 176075 220144
rect 74809 220086 176075 220088
rect 74809 220083 74875 220086
rect 176009 220083 176075 220086
rect 180057 220146 180123 220149
rect 240133 220146 240199 220149
rect 270534 220146 270540 220148
rect 180057 220144 270540 220146
rect 180057 220088 180062 220144
rect 180118 220088 240138 220144
rect 240194 220088 270540 220144
rect 180057 220086 270540 220088
rect 180057 220083 180123 220086
rect 240133 220083 240199 220086
rect 270534 220084 270540 220086
rect 270604 220084 270610 220148
rect 111149 219330 111215 219333
rect 269062 219330 269068 219332
rect 111149 219328 269068 219330
rect 111149 219272 111154 219328
rect 111210 219272 269068 219328
rect 111149 219270 269068 219272
rect 111149 219267 111215 219270
rect 269062 219268 269068 219270
rect 269132 219268 269138 219332
rect 580257 219058 580323 219061
rect 583520 219058 584960 219148
rect 580257 219056 584960 219058
rect 580257 219000 580262 219056
rect 580318 219000 584960 219056
rect 580257 218998 584960 219000
rect 580257 218995 580323 218998
rect 583520 218908 584960 218998
rect 20621 218650 20687 218653
rect 184238 218650 184244 218652
rect 20621 218648 184244 218650
rect 20621 218592 20626 218648
rect 20682 218592 184244 218648
rect 20621 218590 184244 218592
rect 20621 218587 20687 218590
rect 184238 218588 184244 218590
rect 184308 218588 184314 218652
rect 269062 218044 269068 218108
rect 269132 218106 269138 218108
rect 269205 218106 269271 218109
rect 269132 218104 269271 218106
rect 269132 218048 269210 218104
rect 269266 218048 269271 218104
rect 269132 218046 269271 218048
rect 269132 218044 269138 218046
rect 269205 218043 269271 218046
rect 235993 217970 236059 217973
rect 237281 217970 237347 217973
rect 261201 217970 261267 217973
rect 235993 217968 261267 217970
rect 235993 217912 235998 217968
rect 236054 217912 237286 217968
rect 237342 217912 261206 217968
rect 261262 217912 261267 217968
rect 235993 217910 261267 217912
rect 235993 217907 236059 217910
rect 237281 217907 237347 217910
rect 261201 217907 261267 217910
rect 197118 217364 197124 217428
rect 197188 217426 197194 217428
rect 220813 217426 220879 217429
rect 197188 217424 220879 217426
rect 197188 217368 220818 217424
rect 220874 217368 220879 217424
rect 197188 217366 220879 217368
rect 197188 217364 197194 217366
rect 220813 217363 220879 217366
rect 33041 217290 33107 217293
rect 189717 217290 189783 217293
rect 33041 217288 189783 217290
rect 33041 217232 33046 217288
rect 33102 217232 189722 217288
rect 189778 217232 189783 217288
rect 33041 217230 189783 217232
rect 33041 217227 33107 217230
rect 189717 217227 189783 217230
rect 210417 217290 210483 217293
rect 254025 217290 254091 217293
rect 210417 217288 254091 217290
rect 210417 217232 210422 217288
rect 210478 217232 254030 217288
rect 254086 217232 254091 217288
rect 210417 217230 254091 217232
rect 210417 217227 210483 217230
rect 254025 217227 254091 217230
rect 262121 217290 262187 217293
rect 276289 217290 276355 217293
rect 262121 217288 276355 217290
rect 262121 217232 262126 217288
rect 262182 217232 276294 217288
rect 276350 217232 276355 217288
rect 262121 217230 276355 217232
rect 262121 217227 262187 217230
rect 276289 217227 276355 217230
rect 156597 216610 156663 216613
rect 274909 216610 274975 216613
rect 156597 216608 274975 216610
rect 156597 216552 156602 216608
rect 156658 216552 274914 216608
rect 274970 216552 274975 216608
rect 156597 216550 274975 216552
rect 156597 216547 156663 216550
rect 274909 216547 274975 216550
rect 70301 215250 70367 215253
rect 70301 215248 180810 215250
rect 70301 215192 70306 215248
rect 70362 215192 180810 215248
rect 70301 215190 180810 215192
rect 70301 215187 70367 215190
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 69657 214842 69723 214845
rect 70301 214842 70367 214845
rect 69657 214840 70367 214842
rect 69657 214784 69662 214840
rect 69718 214784 70306 214840
rect 70362 214784 70367 214840
rect 69657 214782 70367 214784
rect 69657 214779 69723 214782
rect 70301 214779 70367 214782
rect 180750 214706 180810 215190
rect 182265 214706 182331 214709
rect 202086 214706 202092 214708
rect 180750 214704 202092 214706
rect 180750 214648 182270 214704
rect 182326 214648 202092 214704
rect 180750 214646 202092 214648
rect 182265 214643 182331 214646
rect 202086 214644 202092 214646
rect 202156 214706 202162 214708
rect 260966 214706 260972 214708
rect 202156 214646 260972 214706
rect 202156 214644 202162 214646
rect 260966 214644 260972 214646
rect 261036 214644 261042 214708
rect 202229 214570 202295 214573
rect 273294 214570 273300 214572
rect 202229 214568 273300 214570
rect 202229 214512 202234 214568
rect 202290 214512 273300 214568
rect 202229 214510 273300 214512
rect 202229 214507 202295 214510
rect 273294 214508 273300 214510
rect 273364 214508 273370 214572
rect 72734 213828 72740 213892
rect 72804 213890 72810 213892
rect 271965 213890 272031 213893
rect 72804 213888 272031 213890
rect 72804 213832 271970 213888
rect 272026 213832 272031 213888
rect 72804 213830 272031 213832
rect 72804 213828 72810 213830
rect 271965 213827 272031 213830
rect 71446 211788 71452 211852
rect 71516 211850 71522 211852
rect 254117 211850 254183 211853
rect 71516 211848 254183 211850
rect 71516 211792 254122 211848
rect 254178 211792 254183 211848
rect 71516 211790 254183 211792
rect 71516 211788 71522 211790
rect 254117 211787 254183 211790
rect 97758 210292 97764 210356
rect 97828 210354 97834 210356
rect 106365 210354 106431 210357
rect 97828 210352 106431 210354
rect 97828 210296 106370 210352
rect 106426 210296 106431 210352
rect 97828 210294 106431 210296
rect 97828 210292 97834 210294
rect 106365 210291 106431 210294
rect 106365 209810 106431 209813
rect 270493 209810 270559 209813
rect 106365 209808 270559 209810
rect 106365 209752 106370 209808
rect 106426 209752 270498 209808
rect 270554 209752 270559 209808
rect 106365 209750 270559 209752
rect 106365 209747 106431 209750
rect 270493 209747 270559 209750
rect 204989 208994 205055 208997
rect 210366 208994 210372 208996
rect 204989 208992 210372 208994
rect 204989 208936 204994 208992
rect 205050 208936 210372 208992
rect 204989 208934 210372 208936
rect 204989 208931 205055 208934
rect 210366 208932 210372 208934
rect 210436 208994 210442 208996
rect 253841 208994 253907 208997
rect 210436 208992 253907 208994
rect 210436 208936 253846 208992
rect 253902 208936 253907 208992
rect 210436 208934 253907 208936
rect 210436 208932 210442 208934
rect 253841 208931 253907 208934
rect 97206 205668 97212 205732
rect 97276 205730 97282 205732
rect 201401 205730 201467 205733
rect 97276 205728 201467 205730
rect 97276 205672 201406 205728
rect 201462 205672 201467 205728
rect 97276 205670 201467 205672
rect 97276 205668 97282 205670
rect 201401 205667 201467 205670
rect 580349 205730 580415 205733
rect 583520 205730 584960 205820
rect 580349 205728 584960 205730
rect 580349 205672 580354 205728
rect 580410 205672 584960 205728
rect 580349 205670 584960 205672
rect 580349 205667 580415 205670
rect 583520 205580 584960 205670
rect 255957 204914 256023 204917
rect 266486 204914 266492 204916
rect 255957 204912 266492 204914
rect 255957 204856 255962 204912
rect 256018 204856 266492 204912
rect 255957 204854 266492 204856
rect 255957 204851 256023 204854
rect 266486 204852 266492 204854
rect 266556 204852 266562 204916
rect 6821 203554 6887 203557
rect 184974 203554 184980 203556
rect 6821 203552 184980 203554
rect 6821 203496 6826 203552
rect 6882 203496 184980 203552
rect 6821 203494 184980 203496
rect 6821 203491 6887 203494
rect 184974 203492 184980 203494
rect 185044 203492 185050 203556
rect 195830 202268 195836 202332
rect 195900 202330 195906 202332
rect 209037 202330 209103 202333
rect 195900 202328 209103 202330
rect 195900 202272 209042 202328
rect 209098 202272 209103 202328
rect 195900 202270 209103 202272
rect 195900 202268 195906 202270
rect 209037 202267 209103 202270
rect 171041 202194 171107 202197
rect 253054 202194 253060 202196
rect 171041 202192 253060 202194
rect 171041 202136 171046 202192
rect 171102 202136 253060 202192
rect 171041 202134 253060 202136
rect 171041 202131 171107 202134
rect 253054 202132 253060 202134
rect 253124 202132 253130 202196
rect -960 201922 480 202012
rect 3233 201922 3299 201925
rect -960 201920 3299 201922
rect -960 201864 3238 201920
rect 3294 201864 3299 201920
rect -960 201862 3299 201864
rect -960 201772 480 201862
rect 3233 201859 3299 201862
rect 173249 199338 173315 199341
rect 186814 199338 186820 199340
rect 173249 199336 186820 199338
rect 173249 199280 173254 199336
rect 173310 199280 186820 199336
rect 173249 199278 186820 199280
rect 173249 199275 173315 199278
rect 186814 199276 186820 199278
rect 186884 199276 186890 199340
rect 61837 196618 61903 196621
rect 186998 196618 187004 196620
rect 61837 196616 187004 196618
rect 61837 196560 61842 196616
rect 61898 196560 187004 196616
rect 61837 196558 187004 196560
rect 61837 196555 61903 196558
rect 186998 196556 187004 196558
rect 187068 196556 187074 196620
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 86534 190980 86540 191044
rect 86604 191042 86610 191044
rect 118785 191042 118851 191045
rect 86604 191040 118851 191042
rect 86604 190984 118790 191040
rect 118846 190984 118851 191040
rect 86604 190982 118851 190984
rect 86604 190980 86610 190982
rect 118785 190979 118851 190982
rect 211797 189138 211863 189141
rect 215334 189138 215340 189140
rect 211797 189136 215340 189138
rect 211797 189080 211802 189136
rect 211858 189080 215340 189136
rect 211797 189078 215340 189080
rect 211797 189075 211863 189078
rect 215334 189076 215340 189078
rect 215404 189076 215410 189140
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 24761 186962 24827 186965
rect 184054 186962 184060 186964
rect 24761 186960 184060 186962
rect 24761 186904 24766 186960
rect 24822 186904 184060 186960
rect 24761 186902 184060 186904
rect 24761 186899 24827 186902
rect 184054 186900 184060 186902
rect 184124 186900 184130 186964
rect 211797 186962 211863 186965
rect 262254 186962 262260 186964
rect 211797 186960 262260 186962
rect 211797 186904 211802 186960
rect 211858 186904 262260 186960
rect 211797 186902 262260 186904
rect 211797 186899 211863 186902
rect 262254 186900 262260 186902
rect 262324 186900 262330 186964
rect 104249 182882 104315 182885
rect 148174 182882 148180 182884
rect 104249 182880 148180 182882
rect 104249 182824 104254 182880
rect 104310 182824 148180 182880
rect 104249 182822 148180 182824
rect 104249 182819 104315 182822
rect 148174 182820 148180 182822
rect 148244 182820 148250 182884
rect 69606 180780 69612 180844
rect 69676 180842 69682 180844
rect 160737 180842 160803 180845
rect 69676 180840 160803 180842
rect 69676 180784 160742 180840
rect 160798 180784 160803 180840
rect 69676 180782 160803 180784
rect 69676 180780 69682 180782
rect 160737 180779 160803 180782
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 197261 175946 197327 175949
rect 211654 175946 211660 175948
rect 197261 175944 211660 175946
rect 197261 175888 197266 175944
rect 197322 175888 211660 175944
rect 197261 175886 211660 175888
rect 197261 175883 197327 175886
rect 211654 175884 211660 175886
rect 211724 175884 211730 175948
rect 255313 175810 255379 175813
rect 256049 175810 256115 175813
rect 255313 175808 256115 175810
rect 255313 175752 255318 175808
rect 255374 175752 256054 175808
rect 256110 175752 256115 175808
rect 255313 175750 256115 175752
rect 255313 175747 255379 175750
rect 256049 175747 256115 175750
rect 89069 175402 89135 175405
rect 89478 175402 89484 175404
rect 89069 175400 89484 175402
rect 89069 175344 89074 175400
rect 89130 175344 89484 175400
rect 89069 175342 89484 175344
rect 89069 175339 89135 175342
rect 89478 175340 89484 175342
rect 89548 175402 89554 175404
rect 214005 175402 214071 175405
rect 255313 175402 255379 175405
rect 89548 175400 255379 175402
rect 89548 175344 214010 175400
rect 214066 175344 255318 175400
rect 255374 175344 255379 175400
rect 89548 175342 255379 175344
rect 89548 175340 89554 175342
rect 214005 175339 214071 175342
rect 255313 175339 255379 175342
rect 78673 175266 78739 175269
rect 79317 175266 79383 175269
rect 172421 175266 172487 175269
rect 78673 175264 172487 175266
rect 78673 175208 78678 175264
rect 78734 175208 79322 175264
rect 79378 175208 172426 175264
rect 172482 175208 172487 175264
rect 78673 175206 172487 175208
rect 78673 175203 78739 175206
rect 79317 175203 79383 175206
rect 172421 175203 172487 175206
rect 172421 174586 172487 174589
rect 205633 174586 205699 174589
rect 172421 174584 205699 174586
rect 172421 174528 172426 174584
rect 172482 174528 205638 174584
rect 205694 174528 205699 174584
rect 172421 174526 205699 174528
rect 172421 174523 172487 174526
rect 205633 174523 205699 174526
rect 86217 171186 86283 171189
rect 214557 171186 214623 171189
rect 86217 171184 214623 171186
rect 86217 171128 86222 171184
rect 86278 171128 214562 171184
rect 214618 171128 214623 171184
rect 86217 171126 214623 171128
rect 86217 171123 86283 171126
rect 214557 171123 214623 171126
rect 90950 169764 90956 169828
rect 91020 169826 91026 169828
rect 219525 169826 219591 169829
rect 220261 169826 220327 169829
rect 91020 169824 220327 169826
rect 91020 169768 219530 169824
rect 219586 169768 220266 169824
rect 220322 169768 220327 169824
rect 91020 169766 220327 169768
rect 91020 169764 91026 169766
rect 219525 169763 219591 169766
rect 220261 169763 220327 169766
rect 86718 169084 86724 169148
rect 86788 169146 86794 169148
rect 210417 169146 210483 169149
rect 86788 169144 210483 169146
rect 86788 169088 210422 169144
rect 210478 169088 210483 169144
rect 86788 169086 210483 169088
rect 86788 169084 86794 169086
rect 210417 169083 210483 169086
rect 83457 169012 83523 169013
rect 83406 169010 83412 169012
rect 83330 168950 83412 169010
rect 83476 169010 83523 169012
rect 219433 169010 219499 169013
rect 220353 169010 220419 169013
rect 83476 169008 220419 169010
rect 83518 168952 219438 169008
rect 219494 168952 220358 169008
rect 220414 168952 220419 169008
rect 83406 168948 83412 168950
rect 83476 168950 220419 168952
rect 83476 168948 83523 168950
rect 83457 168947 83523 168948
rect 219433 168947 219499 168950
rect 220353 168947 220419 168950
rect 86309 168466 86375 168469
rect 86718 168466 86724 168468
rect 86309 168464 86724 168466
rect 86309 168408 86314 168464
rect 86370 168408 86724 168464
rect 86309 168406 86724 168408
rect 86309 168403 86375 168406
rect 86718 168404 86724 168406
rect 86788 168404 86794 168468
rect 91001 167786 91067 167789
rect 96654 167786 96660 167788
rect 91001 167784 96660 167786
rect 91001 167728 91006 167784
rect 91062 167728 96660 167784
rect 91001 167726 96660 167728
rect 91001 167723 91067 167726
rect 96654 167724 96660 167726
rect 96724 167724 96730 167788
rect 114461 167786 114527 167789
rect 181437 167786 181503 167789
rect 114461 167784 181503 167786
rect 114461 167728 114466 167784
rect 114522 167728 181442 167784
rect 181498 167728 181503 167784
rect 114461 167726 181503 167728
rect 114461 167723 114527 167726
rect 181437 167723 181503 167726
rect 209037 167786 209103 167789
rect 222326 167786 222332 167788
rect 209037 167784 222332 167786
rect 209037 167728 209042 167784
rect 209098 167728 222332 167784
rect 209037 167726 222332 167728
rect 209037 167723 209103 167726
rect 222326 167724 222332 167726
rect 222396 167724 222402 167788
rect 78857 167650 78923 167653
rect 161289 167650 161355 167653
rect 197997 167650 198063 167653
rect 78857 167648 198063 167650
rect 78857 167592 78862 167648
rect 78918 167592 161294 167648
rect 161350 167592 198002 167648
rect 198058 167592 198063 167648
rect 78857 167590 198063 167592
rect 78857 167587 78923 167590
rect 161289 167587 161355 167590
rect 197997 167587 198063 167590
rect 201401 167650 201467 167653
rect 227662 167650 227668 167652
rect 201401 167648 227668 167650
rect 201401 167592 201406 167648
rect 201462 167592 227668 167648
rect 201401 167590 227668 167592
rect 201401 167587 201467 167590
rect 227662 167588 227668 167590
rect 227732 167588 227738 167652
rect 188429 166426 188495 166429
rect 253197 166426 253263 166429
rect 188429 166424 253263 166426
rect 188429 166368 188434 166424
rect 188490 166368 253202 166424
rect 253258 166368 253263 166424
rect 188429 166366 253263 166368
rect 188429 166363 188495 166366
rect 253197 166363 253263 166366
rect 92657 166290 92723 166293
rect 193213 166290 193279 166293
rect 223665 166290 223731 166293
rect 92657 166288 223731 166290
rect 92657 166232 92662 166288
rect 92718 166232 193218 166288
rect 193274 166232 223670 166288
rect 223726 166232 223731 166288
rect 92657 166230 223731 166232
rect 92657 166227 92723 166230
rect 193213 166227 193279 166230
rect 223665 166227 223731 166230
rect 582925 165882 582991 165885
rect 583520 165882 584960 165972
rect 582925 165880 584960 165882
rect 582925 165824 582930 165880
rect 582986 165824 584960 165880
rect 582925 165822 584960 165824
rect 582925 165819 582991 165822
rect 583520 165732 584960 165822
rect 67725 165610 67791 165613
rect 68686 165610 68692 165612
rect 67725 165608 68692 165610
rect 67725 165552 67730 165608
rect 67786 165552 68692 165608
rect 67725 165550 68692 165552
rect 67725 165547 67791 165550
rect 68686 165548 68692 165550
rect 68756 165548 68762 165612
rect 67725 164386 67791 164389
rect 191925 164386 191991 164389
rect 67725 164384 191991 164386
rect 67725 164328 67730 164384
rect 67786 164328 191930 164384
rect 191986 164328 191991 164384
rect 67725 164326 191991 164328
rect 67725 164323 67791 164326
rect 191925 164323 191991 164326
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 102869 162890 102935 162893
rect 227805 162890 227871 162893
rect 102869 162888 227871 162890
rect 102869 162832 102874 162888
rect 102930 162832 227810 162888
rect 227866 162832 227871 162888
rect 102869 162830 227871 162832
rect 102869 162827 102935 162830
rect 227805 162827 227871 162830
rect 74533 162074 74599 162077
rect 169569 162074 169635 162077
rect 187049 162074 187115 162077
rect 74533 162072 187115 162074
rect 74533 162016 74538 162072
rect 74594 162016 169574 162072
rect 169630 162016 187054 162072
rect 187110 162016 187115 162072
rect 74533 162014 187115 162016
rect 74533 162011 74599 162014
rect 169569 162011 169635 162014
rect 187049 162011 187115 162014
rect 93526 161468 93532 161532
rect 93596 161530 93602 161532
rect 222193 161530 222259 161533
rect 93596 161528 222259 161530
rect 93596 161472 222198 161528
rect 222254 161472 222259 161528
rect 93596 161470 222259 161472
rect 93596 161468 93602 161470
rect 222193 161467 222259 161470
rect 68134 160788 68140 160852
rect 68204 160850 68210 160852
rect 183461 160850 183527 160853
rect 68204 160848 183527 160850
rect 68204 160792 183466 160848
rect 183522 160792 183527 160848
rect 68204 160790 183527 160792
rect 68204 160788 68210 160790
rect 183461 160787 183527 160790
rect 54937 160714 55003 160717
rect 191046 160714 191052 160716
rect 54937 160712 191052 160714
rect 54937 160656 54942 160712
rect 54998 160656 191052 160712
rect 54937 160654 191052 160656
rect 54937 160651 55003 160654
rect 191046 160652 191052 160654
rect 191116 160652 191122 160716
rect 127801 158810 127867 158813
rect 229093 158810 229159 158813
rect 127801 158808 229159 158810
rect 127801 158752 127806 158808
rect 127862 158752 229098 158808
rect 229154 158752 229159 158808
rect 127801 158750 229159 158752
rect 127801 158747 127867 158750
rect 229093 158747 229159 158750
rect 194358 157932 194364 157996
rect 194428 157994 194434 157996
rect 234613 157994 234679 157997
rect 194428 157992 234679 157994
rect 194428 157936 234618 157992
rect 234674 157936 234679 157992
rect 194428 157934 234679 157936
rect 194428 157932 194434 157934
rect 234613 157931 234679 157934
rect 79961 157450 80027 157453
rect 208393 157450 208459 157453
rect 208577 157450 208643 157453
rect 79961 157448 208643 157450
rect 79961 157392 79966 157448
rect 80022 157392 208398 157448
rect 208454 157392 208582 157448
rect 208638 157392 208643 157448
rect 79961 157390 208643 157392
rect 79961 157387 80027 157390
rect 208393 157387 208459 157390
rect 208577 157387 208643 157390
rect 10961 156634 11027 156637
rect 186957 156634 187023 156637
rect 10961 156632 187023 156634
rect 10961 156576 10966 156632
rect 11022 156576 186962 156632
rect 187018 156576 187023 156632
rect 10961 156574 187023 156576
rect 10961 156571 11027 156574
rect 186957 156571 187023 156574
rect 148501 156090 148567 156093
rect 227713 156090 227779 156093
rect 148501 156088 227779 156090
rect 148501 156032 148506 156088
rect 148562 156032 227718 156088
rect 227774 156032 227779 156088
rect 148501 156030 227779 156032
rect 148501 156027 148567 156030
rect 227713 156027 227779 156030
rect 160737 155274 160803 155277
rect 188613 155274 188679 155277
rect 160737 155272 188679 155274
rect 160737 155216 160742 155272
rect 160798 155216 188618 155272
rect 188674 155216 188679 155272
rect 160737 155214 188679 155216
rect 160737 155211 160803 155214
rect 188613 155211 188679 155214
rect 190361 155274 190427 155277
rect 201585 155274 201651 155277
rect 190361 155272 201651 155274
rect 190361 155216 190366 155272
rect 190422 155216 201590 155272
rect 201646 155216 201651 155272
rect 190361 155214 201651 155216
rect 190361 155211 190427 155214
rect 201585 155211 201651 155214
rect 88333 154594 88399 154597
rect 218237 154594 218303 154597
rect 88333 154592 218303 154594
rect 88333 154536 88338 154592
rect 88394 154536 218242 154592
rect 218298 154536 218303 154592
rect 88333 154534 218303 154536
rect 88333 154531 88399 154534
rect 218237 154531 218303 154534
rect 220261 154594 220327 154597
rect 582833 154594 582899 154597
rect 220261 154592 582899 154594
rect 220261 154536 220266 154592
rect 220322 154536 582838 154592
rect 582894 154536 582899 154592
rect 220261 154534 582899 154536
rect 220261 154531 220327 154534
rect 582833 154531 582899 154534
rect 81433 153778 81499 153781
rect 177389 153778 177455 153781
rect 204989 153778 205055 153781
rect 81433 153776 205055 153778
rect 81433 153720 81438 153776
rect 81494 153720 177394 153776
rect 177450 153720 204994 153776
rect 205050 153720 205055 153776
rect 81433 153718 205055 153720
rect 81433 153715 81499 153718
rect 177389 153715 177455 153718
rect 204989 153715 205055 153718
rect 208485 153778 208551 153781
rect 281717 153778 281783 153781
rect 208485 153776 281783 153778
rect 208485 153720 208490 153776
rect 208546 153720 281722 153776
rect 281778 153720 281783 153776
rect 208485 153718 281783 153720
rect 208485 153715 208551 153718
rect 281717 153715 281783 153718
rect 155401 153234 155467 153237
rect 240133 153234 240199 153237
rect 155401 153232 240199 153234
rect 155401 153176 155406 153232
rect 155462 153176 240138 153232
rect 240194 153176 240199 153232
rect 155401 153174 240199 153176
rect 155401 153171 155467 153174
rect 240133 153171 240199 153174
rect 70485 153098 70551 153101
rect 71630 153098 71636 153100
rect 70485 153096 71636 153098
rect 70485 153040 70490 153096
rect 70546 153040 71636 153096
rect 70485 153038 71636 153040
rect 70485 153035 70551 153038
rect 71630 153036 71636 153038
rect 71700 153036 71706 153100
rect 218053 153098 218119 153101
rect 218237 153098 218303 153101
rect 267825 153098 267891 153101
rect 218053 153096 267891 153098
rect 218053 153040 218058 153096
rect 218114 153040 218242 153096
rect 218298 153040 267830 153096
rect 267886 153040 267891 153096
rect 218053 153038 267891 153040
rect 218053 153035 218119 153038
rect 218237 153035 218303 153038
rect 267825 153035 267891 153038
rect 582649 152690 582715 152693
rect 583520 152690 584960 152780
rect 582649 152688 584960 152690
rect 582649 152632 582654 152688
rect 582710 152632 584960 152688
rect 582649 152630 584960 152632
rect 582649 152627 582715 152630
rect 583520 152540 584960 152630
rect 71630 152084 71636 152148
rect 71700 152146 71706 152148
rect 196065 152146 196131 152149
rect 71700 152144 196131 152146
rect 71700 152088 196070 152144
rect 196126 152088 196131 152144
rect 71700 152086 196131 152088
rect 71700 152084 71706 152086
rect 196065 152083 196131 152086
rect 195881 152010 195947 152013
rect 281441 152010 281507 152013
rect 195881 152008 281507 152010
rect 195881 151952 195886 152008
rect 195942 151952 281446 152008
rect 281502 151952 281507 152008
rect 195881 151950 281507 151952
rect 195881 151947 195947 151950
rect 281441 151947 281507 151950
rect 80237 151874 80303 151877
rect 208485 151874 208551 151877
rect 80237 151872 208551 151874
rect 80237 151816 80242 151872
rect 80298 151816 208490 151872
rect 208546 151816 208551 151872
rect 80237 151814 208551 151816
rect 80237 151811 80303 151814
rect 208485 151811 208551 151814
rect 64505 151058 64571 151061
rect 161473 151058 161539 151061
rect 64505 151056 161539 151058
rect 64505 151000 64510 151056
rect 64566 151000 161478 151056
rect 161534 151000 161539 151056
rect 64505 150998 161539 151000
rect 64505 150995 64571 150998
rect 161473 150995 161539 150998
rect 160829 150650 160895 150653
rect 259453 150650 259519 150653
rect 160829 150648 259519 150650
rect 160829 150592 160834 150648
rect 160890 150592 259458 150648
rect 259514 150592 259519 150648
rect 160829 150590 259519 150592
rect 160829 150587 160895 150590
rect 259453 150587 259519 150590
rect 104801 150514 104867 150517
rect 227989 150514 228055 150517
rect 104801 150512 228055 150514
rect 104801 150456 104806 150512
rect 104862 150456 227994 150512
rect 228050 150456 228055 150512
rect 104801 150454 228055 150456
rect 104801 150451 104867 150454
rect 227989 150451 228055 150454
rect -960 149834 480 149924
rect 3141 149834 3207 149837
rect -960 149832 3207 149834
rect -960 149776 3146 149832
rect 3202 149776 3207 149832
rect -960 149774 3207 149776
rect -960 149684 480 149774
rect 3141 149771 3207 149774
rect 197997 149834 198063 149837
rect 207105 149834 207171 149837
rect 197997 149832 207171 149834
rect 197997 149776 198002 149832
rect 198058 149776 207110 149832
rect 207166 149776 207171 149832
rect 197997 149774 207171 149776
rect 197997 149771 198063 149774
rect 207105 149771 207171 149774
rect 116669 149698 116735 149701
rect 213821 149698 213887 149701
rect 224902 149698 224908 149700
rect 116669 149696 224908 149698
rect 116669 149640 116674 149696
rect 116730 149640 213826 149696
rect 213882 149640 224908 149696
rect 116669 149638 224908 149640
rect 116669 149635 116735 149638
rect 213821 149635 213887 149638
rect 224902 149636 224908 149638
rect 224972 149636 224978 149700
rect 177389 149154 177455 149157
rect 220997 149154 221063 149157
rect 222009 149154 222075 149157
rect 177389 149152 222075 149154
rect 177389 149096 177394 149152
rect 177450 149096 221002 149152
rect 221058 149096 222014 149152
rect 222070 149096 222075 149152
rect 177389 149094 222075 149096
rect 177389 149091 177455 149094
rect 220997 149091 221063 149094
rect 222009 149091 222075 149094
rect 198825 148474 198891 148477
rect 213177 148474 213243 148477
rect 198825 148472 213243 148474
rect 198825 148416 198830 148472
rect 198886 148416 213182 148472
rect 213238 148416 213243 148472
rect 198825 148414 213243 148416
rect 198825 148411 198891 148414
rect 213177 148411 213243 148414
rect 231761 148474 231827 148477
rect 285622 148474 285628 148476
rect 231761 148472 285628 148474
rect 231761 148416 231766 148472
rect 231822 148416 285628 148472
rect 231761 148414 285628 148416
rect 231761 148411 231827 148414
rect 285622 148412 285628 148414
rect 285692 148412 285698 148476
rect 215201 148338 215267 148341
rect 317413 148338 317479 148341
rect 215201 148336 317479 148338
rect 215201 148280 215206 148336
rect 215262 148280 317418 148336
rect 317474 148280 317479 148336
rect 215201 148278 317479 148280
rect 215201 148275 215267 148278
rect 317413 148275 317479 148278
rect 194685 147930 194751 147933
rect 247677 147930 247743 147933
rect 194685 147928 247743 147930
rect 194685 147872 194690 147928
rect 194746 147872 247682 147928
rect 247738 147872 247743 147928
rect 194685 147870 247743 147872
rect 194685 147867 194751 147870
rect 247677 147867 247743 147870
rect 73337 147794 73403 147797
rect 200297 147794 200363 147797
rect 201401 147794 201467 147797
rect 73337 147792 201467 147794
rect 73337 147736 73342 147792
rect 73398 147736 200302 147792
rect 200358 147736 201406 147792
rect 201462 147736 201467 147792
rect 73337 147734 201467 147736
rect 73337 147731 73403 147734
rect 200297 147731 200363 147734
rect 201401 147731 201467 147734
rect 212349 147794 212415 147797
rect 215201 147794 215267 147797
rect 212349 147792 215267 147794
rect 212349 147736 212354 147792
rect 212410 147736 215206 147792
rect 215262 147736 215267 147792
rect 212349 147734 215267 147736
rect 212349 147731 212415 147734
rect 215201 147731 215267 147734
rect 204345 147658 204411 147661
rect 211797 147658 211863 147661
rect 204345 147656 211863 147658
rect 204345 147600 204350 147656
rect 204406 147600 211802 147656
rect 211858 147600 211863 147656
rect 204345 147598 211863 147600
rect 204345 147595 204411 147598
rect 211797 147595 211863 147598
rect 71773 146978 71839 146981
rect 108481 146978 108547 146981
rect 259494 146978 259500 146980
rect 71773 146976 108547 146978
rect 71773 146920 71778 146976
rect 71834 146920 108486 146976
rect 108542 146920 108547 146976
rect 71773 146918 108547 146920
rect 71773 146915 71839 146918
rect 108481 146915 108547 146918
rect 229050 146918 259500 146978
rect 170581 146570 170647 146573
rect 226793 146570 226859 146573
rect 229050 146570 229110 146918
rect 259494 146916 259500 146918
rect 259564 146916 259570 146980
rect 170581 146568 229110 146570
rect 170581 146512 170586 146568
rect 170642 146512 226798 146568
rect 226854 146512 229110 146568
rect 170581 146510 229110 146512
rect 170581 146507 170647 146510
rect 226793 146507 226859 146510
rect 97942 146372 97948 146436
rect 98012 146434 98018 146436
rect 98821 146434 98887 146437
rect 229185 146434 229251 146437
rect 98012 146432 229251 146434
rect 98012 146376 98826 146432
rect 98882 146376 229190 146432
rect 229246 146376 229251 146432
rect 98012 146374 229251 146376
rect 98012 146372 98018 146374
rect 98821 146371 98887 146374
rect 229185 146371 229251 146374
rect 222009 146298 222075 146301
rect 226374 146298 226380 146300
rect 222009 146296 226380 146298
rect 222009 146240 222014 146296
rect 222070 146240 226380 146296
rect 222009 146238 226380 146240
rect 222009 146235 222075 146238
rect 226374 146236 226380 146238
rect 226444 146236 226450 146300
rect 3141 145754 3207 145757
rect 96705 145754 96771 145757
rect 104801 145754 104867 145757
rect 3141 145752 104867 145754
rect 3141 145696 3146 145752
rect 3202 145696 96710 145752
rect 96766 145696 104806 145752
rect 104862 145696 104867 145752
rect 3141 145694 104867 145696
rect 3141 145691 3207 145694
rect 96705 145691 96771 145694
rect 104801 145691 104867 145694
rect 74809 145618 74875 145621
rect 175181 145618 175247 145621
rect 201585 145618 201651 145621
rect 252461 145618 252527 145621
rect 74809 145616 201651 145618
rect 74809 145560 74814 145616
rect 74870 145560 175186 145616
rect 175242 145560 201590 145616
rect 201646 145560 201651 145616
rect 74809 145558 201651 145560
rect 74809 145555 74875 145558
rect 175181 145555 175247 145558
rect 201585 145555 201651 145558
rect 229050 145616 252527 145618
rect 229050 145560 252466 145616
rect 252522 145560 252527 145616
rect 229050 145558 252527 145560
rect 188521 145074 188587 145077
rect 226558 145074 226564 145076
rect 188521 145072 226564 145074
rect 188521 145016 188526 145072
rect 188582 145016 226564 145072
rect 188521 145014 226564 145016
rect 188521 145011 188587 145014
rect 226558 145012 226564 145014
rect 226628 145074 226634 145076
rect 229050 145074 229110 145558
rect 252461 145555 252527 145558
rect 226628 145014 229110 145074
rect 226628 145012 226634 145014
rect 102961 144938 103027 144941
rect 230473 144938 230539 144941
rect 231117 144938 231183 144941
rect 102961 144936 231183 144938
rect 102961 144880 102966 144936
rect 103022 144880 230478 144936
rect 230534 144880 231122 144936
rect 231178 144880 231183 144936
rect 102961 144878 231183 144880
rect 102961 144875 103027 144878
rect 230473 144875 230539 144878
rect 231117 144875 231183 144878
rect 213269 144802 213335 144805
rect 285857 144802 285923 144805
rect 286777 144802 286843 144805
rect 213269 144800 286843 144802
rect 213269 144744 213274 144800
rect 213330 144744 285862 144800
rect 285918 144744 286782 144800
rect 286838 144744 286843 144800
rect 213269 144742 286843 144744
rect 213269 144739 213335 144742
rect 285857 144739 285923 144742
rect 286777 144739 286843 144742
rect 222285 144666 222351 144669
rect 223021 144666 223087 144669
rect 222285 144664 223087 144666
rect 222285 144608 222290 144664
rect 222346 144608 223026 144664
rect 223082 144608 223087 144664
rect 222285 144606 223087 144608
rect 222285 144603 222351 144606
rect 223021 144603 223087 144606
rect 188613 144258 188679 144261
rect 193581 144258 193647 144261
rect 188613 144256 193647 144258
rect 188613 144200 188618 144256
rect 188674 144200 193586 144256
rect 193642 144200 193647 144256
rect 188613 144198 193647 144200
rect 188613 144195 188679 144198
rect 193581 144195 193647 144198
rect 187049 144122 187115 144125
rect 201309 144122 201375 144125
rect 187049 144120 201375 144122
rect 187049 144064 187054 144120
rect 187110 144064 201314 144120
rect 201370 144064 201375 144120
rect 187049 144062 201375 144064
rect 187049 144059 187115 144062
rect 201309 144059 201375 144062
rect 59169 143714 59235 143717
rect 108389 143714 108455 143717
rect 59169 143712 108455 143714
rect 59169 143656 59174 143712
rect 59230 143656 108394 143712
rect 108450 143656 108455 143712
rect 59169 143654 108455 143656
rect 59169 143651 59235 143654
rect 108389 143651 108455 143654
rect 183093 143714 183159 143717
rect 223021 143714 223087 143717
rect 183093 143712 223087 143714
rect 183093 143656 183098 143712
rect 183154 143656 223026 143712
rect 223082 143656 223087 143712
rect 183093 143654 223087 143656
rect 183093 143651 183159 143654
rect 223021 143651 223087 143654
rect 82997 143578 83063 143581
rect 188429 143578 188495 143581
rect 82997 143576 188495 143578
rect 82997 143520 83002 143576
rect 83058 143520 188434 143576
rect 188490 143520 188495 143576
rect 82997 143518 188495 143520
rect 82997 143515 83063 143518
rect 188429 143515 188495 143518
rect 196617 143578 196683 143581
rect 229277 143578 229343 143581
rect 231761 143578 231827 143581
rect 196617 143576 231827 143578
rect 196617 143520 196622 143576
rect 196678 143520 229282 143576
rect 229338 143520 231766 143576
rect 231822 143520 231827 143576
rect 196617 143518 231827 143520
rect 196617 143515 196683 143518
rect 229277 143515 229343 143518
rect 231761 143515 231827 143518
rect 70577 143442 70643 143445
rect 155861 143442 155927 143445
rect 194685 143442 194751 143445
rect 70577 143440 194751 143442
rect 70577 143384 70582 143440
rect 70638 143384 155866 143440
rect 155922 143384 194690 143440
rect 194746 143384 194751 143440
rect 70577 143382 194751 143384
rect 70577 143379 70643 143382
rect 155861 143379 155927 143382
rect 194685 143379 194751 143382
rect 196157 143442 196223 143445
rect 196566 143442 196572 143444
rect 196157 143440 196572 143442
rect 196157 143384 196162 143440
rect 196218 143384 196572 143440
rect 196157 143382 196572 143384
rect 196157 143379 196223 143382
rect 196566 143380 196572 143382
rect 196636 143380 196642 143444
rect 83457 142490 83523 142493
rect 212349 142490 212415 142493
rect 83457 142488 212415 142490
rect 83457 142432 83462 142488
rect 83518 142432 212354 142488
rect 212410 142432 212415 142488
rect 83457 142430 212415 142432
rect 83457 142427 83523 142430
rect 212349 142427 212415 142430
rect 218237 142490 218303 142493
rect 291837 142490 291903 142493
rect 218237 142488 291903 142490
rect 218237 142432 218242 142488
rect 218298 142432 291842 142488
rect 291898 142432 291903 142488
rect 218237 142430 291903 142432
rect 218237 142427 218303 142430
rect 291837 142427 291903 142430
rect 73470 142292 73476 142356
rect 73540 142354 73546 142356
rect 196566 142354 196572 142356
rect 73540 142294 196572 142354
rect 73540 142292 73546 142294
rect 196566 142292 196572 142294
rect 196636 142292 196642 142356
rect 221917 142218 221983 142221
rect 224350 142218 224356 142220
rect 221917 142216 224356 142218
rect 221917 142160 221922 142216
rect 221978 142160 224356 142216
rect 221917 142158 224356 142160
rect 221917 142155 221983 142158
rect 224350 142156 224356 142158
rect 224420 142156 224426 142220
rect 193070 141068 193076 141132
rect 193140 141130 193146 141132
rect 195237 141130 195303 141133
rect 193140 141128 195303 141130
rect 193140 141072 195242 141128
rect 195298 141072 195303 141128
rect 193140 141070 195303 141072
rect 193140 141068 193146 141070
rect 195237 141067 195303 141070
rect 69790 140932 69796 140996
rect 69860 140994 69866 140996
rect 75913 140994 75979 140997
rect 202873 140994 202939 140997
rect 69860 140934 74550 140994
rect 69860 140932 69866 140934
rect 66161 140858 66227 140861
rect 69289 140858 69355 140861
rect 66161 140856 69355 140858
rect 66161 140800 66166 140856
rect 66222 140800 69294 140856
rect 69350 140800 69355 140856
rect 66161 140798 69355 140800
rect 66161 140795 66227 140798
rect 69289 140795 69355 140798
rect 71129 140858 71195 140861
rect 73470 140858 73476 140860
rect 71129 140856 73476 140858
rect 71129 140800 71134 140856
rect 71190 140800 73476 140856
rect 71129 140798 73476 140800
rect 71129 140795 71195 140798
rect 73470 140796 73476 140798
rect 73540 140796 73546 140860
rect 74490 140858 74550 140934
rect 75913 140992 202939 140994
rect 75913 140936 75918 140992
rect 75974 140936 202878 140992
rect 202934 140936 202939 140992
rect 75913 140934 202939 140936
rect 75913 140931 75979 140934
rect 202873 140931 202939 140934
rect 205449 140994 205515 140997
rect 256601 140994 256667 140997
rect 260097 140994 260163 140997
rect 205449 140992 260163 140994
rect 205449 140936 205454 140992
rect 205510 140936 256606 140992
rect 256662 140936 260102 140992
rect 260158 140936 260163 140992
rect 205449 140934 260163 140936
rect 205449 140931 205515 140934
rect 256601 140931 256667 140934
rect 260097 140931 260163 140934
rect 91093 140858 91159 140861
rect 74490 140856 91159 140858
rect 74490 140800 91098 140856
rect 91154 140800 91159 140856
rect 74490 140798 91159 140800
rect 91093 140795 91159 140798
rect 93669 140858 93735 140861
rect 223573 140858 223639 140861
rect 93669 140856 223639 140858
rect 93669 140800 93674 140856
rect 93730 140800 223578 140856
rect 223634 140800 223639 140856
rect 93669 140798 223639 140800
rect 93669 140795 93735 140798
rect 223573 140795 223639 140798
rect 206553 140586 206619 140589
rect 200070 140584 206619 140586
rect 200070 140528 206558 140584
rect 206614 140528 206619 140584
rect 200070 140526 206619 140528
rect 196566 140388 196572 140452
rect 196636 140450 196642 140452
rect 196801 140450 196867 140453
rect 196636 140448 196867 140450
rect 196636 140392 196806 140448
rect 196862 140392 196867 140448
rect 196636 140390 196867 140392
rect 196636 140388 196642 140390
rect 196801 140387 196867 140390
rect 193438 140116 193444 140180
rect 193508 140178 193514 140180
rect 200070 140178 200130 140526
rect 206553 140523 206619 140526
rect 206553 140450 206619 140453
rect 206870 140450 206876 140452
rect 206553 140448 206876 140450
rect 206553 140392 206558 140448
rect 206614 140392 206876 140448
rect 206553 140390 206876 140392
rect 206553 140387 206619 140390
rect 206870 140388 206876 140390
rect 206940 140388 206946 140452
rect 224493 140450 224559 140453
rect 225270 140450 225276 140452
rect 224493 140448 225276 140450
rect 224493 140392 224498 140448
rect 224554 140392 225276 140448
rect 224493 140390 225276 140392
rect 224493 140387 224559 140390
rect 225270 140388 225276 140390
rect 225340 140388 225346 140452
rect 193508 140118 200130 140178
rect 193508 140116 193514 140118
rect 222326 140116 222332 140180
rect 222396 140178 222402 140180
rect 225321 140178 225387 140181
rect 222396 140176 225387 140178
rect 222396 140120 225326 140176
rect 225382 140120 225387 140176
rect 222396 140118 225387 140120
rect 222396 140116 222402 140118
rect 225321 140115 225387 140118
rect 94221 140042 94287 140045
rect 145649 140042 145715 140045
rect 94221 140040 145715 140042
rect 94221 139984 94226 140040
rect 94282 139984 145654 140040
rect 145710 139984 145715 140040
rect 94221 139982 145715 139984
rect 94221 139979 94287 139982
rect 145649 139979 145715 139982
rect 160921 140042 160987 140045
rect 193305 140042 193371 140045
rect 160921 140040 193371 140042
rect 160921 139984 160926 140040
rect 160982 139984 193310 140040
rect 193366 139984 193371 140040
rect 160921 139982 193371 139984
rect 160921 139979 160987 139982
rect 193305 139979 193371 139982
rect 191649 139906 191715 139909
rect 226558 139906 226564 139908
rect 191649 139904 193660 139906
rect 191649 139848 191654 139904
rect 191710 139848 193660 139904
rect 191649 139846 193660 139848
rect 224940 139846 226564 139906
rect 191649 139843 191715 139846
rect 226558 139844 226564 139846
rect 226628 139844 226634 139908
rect 63217 139634 63283 139637
rect 89989 139634 90055 139637
rect 63217 139632 90055 139634
rect 63217 139576 63222 139632
rect 63278 139576 89994 139632
rect 90050 139576 90055 139632
rect 63217 139574 90055 139576
rect 63217 139571 63283 139574
rect 89989 139571 90055 139574
rect 53281 139498 53347 139501
rect 53649 139498 53715 139501
rect 104341 139498 104407 139501
rect 53281 139496 104407 139498
rect 53281 139440 53286 139496
rect 53342 139440 53654 139496
rect 53710 139440 104346 139496
rect 104402 139440 104407 139496
rect 53281 139438 104407 139440
rect 53281 139435 53347 139438
rect 53649 139435 53715 139438
rect 104341 139435 104407 139438
rect 583017 139362 583083 139365
rect 583520 139362 584960 139452
rect 583017 139360 584960 139362
rect 583017 139304 583022 139360
rect 583078 139304 584960 139360
rect 583017 139302 584960 139304
rect 583017 139299 583083 139302
rect 583520 139212 584960 139302
rect 193070 139028 193076 139092
rect 193140 139090 193146 139092
rect 227621 139090 227687 139093
rect 193140 139030 193660 139090
rect 224940 139088 227687 139090
rect 224940 139032 227626 139088
rect 227682 139032 227687 139088
rect 224940 139030 227687 139032
rect 193140 139028 193146 139030
rect 227621 139027 227687 139030
rect 57605 138818 57671 138821
rect 82997 138818 83063 138821
rect 57605 138816 83063 138818
rect 57605 138760 57610 138816
rect 57666 138760 83002 138816
rect 83058 138760 83063 138816
rect 57605 138758 83063 138760
rect 57605 138755 57671 138758
rect 82997 138755 83063 138758
rect 84653 138818 84719 138821
rect 117957 138818 118023 138821
rect 84653 138816 118023 138818
rect 84653 138760 84658 138816
rect 84714 138760 117962 138816
rect 118018 138760 118023 138816
rect 84653 138758 118023 138760
rect 84653 138755 84719 138758
rect 117957 138755 118023 138758
rect 52177 138682 52243 138685
rect 72325 138682 72391 138685
rect 52177 138680 72391 138682
rect 52177 138624 52182 138680
rect 52238 138624 72330 138680
rect 72386 138624 72391 138680
rect 52177 138622 72391 138624
rect 52177 138619 52243 138622
rect 72325 138619 72391 138622
rect 78121 138682 78187 138685
rect 193397 138682 193463 138685
rect 227805 138682 227871 138685
rect 582649 138682 582715 138685
rect 78121 138680 193463 138682
rect 78121 138624 78126 138680
rect 78182 138624 193402 138680
rect 193458 138624 193463 138680
rect 78121 138622 193463 138624
rect 78121 138619 78187 138622
rect 193397 138619 193463 138622
rect 224910 138680 582715 138682
rect 224910 138624 227810 138680
rect 227866 138624 582654 138680
rect 582710 138624 582715 138680
rect 224910 138622 582715 138624
rect 192702 138212 192708 138276
rect 192772 138274 192778 138276
rect 193029 138274 193095 138277
rect 192772 138272 193660 138274
rect 192772 138216 193034 138272
rect 193090 138216 193660 138272
rect 224910 138244 224970 138622
rect 227805 138619 227871 138622
rect 582649 138619 582715 138622
rect 192772 138214 193660 138216
rect 192772 138212 192778 138214
rect 193029 138211 193095 138214
rect 67817 138002 67883 138005
rect 76097 138002 76163 138005
rect 84745 138004 84811 138005
rect 84694 138002 84700 138004
rect 67817 138000 76163 138002
rect 67817 137944 67822 138000
rect 67878 137944 76102 138000
rect 76158 137944 76163 138000
rect 67817 137942 76163 137944
rect 84654 137942 84700 138002
rect 84764 138000 84811 138004
rect 84806 137944 84811 138000
rect 67817 137939 67883 137942
rect 76097 137939 76163 137942
rect 84694 137940 84700 137942
rect 84764 137940 84811 137944
rect 84745 137939 84811 137940
rect 115933 138002 115999 138005
rect 116485 138002 116551 138005
rect 193438 138002 193444 138004
rect 115933 138000 193444 138002
rect 115933 137944 115938 138000
rect 115994 137944 116490 138000
rect 116546 137944 193444 138000
rect 115933 137942 193444 137944
rect 115933 137939 115999 137942
rect 116485 137939 116551 137942
rect 193438 137940 193444 137942
rect 193508 137940 193514 138004
rect 91093 137866 91159 137869
rect 166349 137866 166415 137869
rect 91093 137864 166415 137866
rect 91093 137808 91098 137864
rect 91154 137808 166354 137864
rect 166410 137808 166415 137864
rect 91093 137806 166415 137808
rect 91093 137803 91159 137806
rect 166349 137803 166415 137806
rect 69841 137458 69907 137461
rect 80697 137458 80763 137461
rect 69841 137456 80763 137458
rect 69841 137400 69846 137456
rect 69902 137400 80702 137456
rect 80758 137400 80763 137456
rect 69841 137398 80763 137400
rect 69841 137395 69907 137398
rect 80697 137395 80763 137398
rect 191649 137458 191715 137461
rect 191649 137456 193660 137458
rect 191649 137400 191654 137456
rect 191710 137400 193660 137456
rect 191649 137398 193660 137400
rect 191649 137395 191715 137398
rect 79317 137322 79383 137325
rect 116485 137322 116551 137325
rect 79317 137320 116551 137322
rect 79317 137264 79322 137320
rect 79378 137264 116490 137320
rect 116546 137264 116551 137320
rect 79317 137262 116551 137264
rect 79317 137259 79383 137262
rect 116485 137259 116551 137262
rect 225270 137260 225276 137324
rect 225340 137322 225346 137324
rect 313273 137322 313339 137325
rect 225340 137320 313339 137322
rect 225340 137264 313278 137320
rect 313334 137264 313339 137320
rect 225340 137262 313339 137264
rect 225340 137260 225346 137262
rect 313273 137259 313339 137262
rect 226517 137186 226583 137189
rect 224940 137184 226583 137186
rect 224940 137128 226522 137184
rect 226578 137128 226583 137184
rect 224940 137126 226583 137128
rect 226517 137123 226583 137126
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 51717 136778 51783 136781
rect 75361 136778 75427 136781
rect 51717 136776 75427 136778
rect 51717 136720 51722 136776
rect 51778 136720 75366 136776
rect 75422 136720 75427 136776
rect 51717 136718 75427 136720
rect 51717 136715 51783 136718
rect 75361 136715 75427 136718
rect 89713 136778 89779 136781
rect 90950 136778 90956 136780
rect 89713 136776 90956 136778
rect 89713 136720 89718 136776
rect 89774 136720 90956 136776
rect 89713 136718 90956 136720
rect 89713 136715 89779 136718
rect 90950 136716 90956 136718
rect 91020 136716 91026 136780
rect 92565 136778 92631 136781
rect 93526 136778 93532 136780
rect 92565 136776 93532 136778
rect 92565 136720 92570 136776
rect 92626 136720 93532 136776
rect 92565 136718 93532 136720
rect 92565 136715 92631 136718
rect 93526 136716 93532 136718
rect 93596 136716 93602 136780
rect 89989 136642 90055 136645
rect 158069 136642 158135 136645
rect 89989 136640 158135 136642
rect 89989 136584 89994 136640
rect 90050 136584 158074 136640
rect 158130 136584 158135 136640
rect 89989 136582 158135 136584
rect 89989 136579 90055 136582
rect 158069 136579 158135 136582
rect 191741 136370 191807 136373
rect 226793 136370 226859 136373
rect 191741 136368 193660 136370
rect 191741 136312 191746 136368
rect 191802 136312 193660 136368
rect 191741 136310 193660 136312
rect 224940 136368 226859 136370
rect 224940 136312 226798 136368
rect 226854 136312 226859 136368
rect 224940 136310 226859 136312
rect 191741 136307 191807 136310
rect 226793 136307 226859 136310
rect 65926 135900 65932 135964
rect 65996 135962 66002 135964
rect 161381 135962 161447 135965
rect 180057 135962 180123 135965
rect 65996 135960 180123 135962
rect 65996 135904 161386 135960
rect 161442 135904 180062 135960
rect 180118 135904 180123 135960
rect 65996 135902 180123 135904
rect 65996 135900 66002 135902
rect 161381 135899 161447 135902
rect 180057 135899 180123 135902
rect 191741 135554 191807 135557
rect 226517 135554 226583 135557
rect 191741 135552 193660 135554
rect 191741 135496 191746 135552
rect 191802 135496 193660 135552
rect 191741 135494 193660 135496
rect 224940 135552 226583 135554
rect 224940 135496 226522 135552
rect 226578 135496 226583 135552
rect 224940 135494 226583 135496
rect 191741 135491 191807 135494
rect 226517 135491 226583 135494
rect 70301 135010 70367 135013
rect 69430 135008 70367 135010
rect 69430 134952 70306 135008
rect 70362 134952 70367 135008
rect 69430 134950 70367 134952
rect 69430 134436 69490 134950
rect 70301 134947 70367 134950
rect 226701 134738 226767 134741
rect 226977 134738 227043 134741
rect 224940 134736 227043 134738
rect 190269 134194 190335 134197
rect 193630 134194 193690 134708
rect 224940 134680 226706 134736
rect 226762 134680 226982 134736
rect 227038 134680 227043 134736
rect 224940 134678 227043 134680
rect 226701 134675 226767 134678
rect 226977 134675 227043 134678
rect 190269 134192 193690 134194
rect 190269 134136 190274 134192
rect 190330 134136 193690 134192
rect 190269 134134 193690 134136
rect 190269 134131 190335 134134
rect 95182 133996 95188 134060
rect 95252 134058 95258 134060
rect 96061 134058 96127 134061
rect 95252 134056 96127 134058
rect 95252 134000 96066 134056
rect 96122 134000 96127 134056
rect 95252 133998 96127 134000
rect 95252 133996 95258 133998
rect 96061 133995 96127 133998
rect 96797 133922 96863 133925
rect 94668 133920 96863 133922
rect 94668 133864 96802 133920
rect 96858 133864 96863 133920
rect 94668 133862 96863 133864
rect 96797 133859 96863 133862
rect 186957 133922 187023 133925
rect 186957 133920 193660 133922
rect 186957 133864 186962 133920
rect 187018 133864 193660 133920
rect 186957 133862 193660 133864
rect 186957 133859 187023 133862
rect 226701 133650 226767 133653
rect 224940 133648 226767 133650
rect 69430 133516 69490 133620
rect 224940 133592 226706 133648
rect 226762 133592 226767 133648
rect 224940 133590 226767 133592
rect 226701 133587 226767 133590
rect 69422 133452 69428 133516
rect 69492 133452 69498 133516
rect 96613 133106 96679 133109
rect 94668 133104 96679 133106
rect 94668 133048 96618 133104
rect 96674 133048 96679 133104
rect 94668 133046 96679 133048
rect 96613 133043 96679 133046
rect 67725 132834 67791 132837
rect 191741 132834 191807 132837
rect 226885 132834 226951 132837
rect 67725 132832 68908 132834
rect 67725 132776 67730 132832
rect 67786 132776 68908 132832
rect 67725 132774 68908 132776
rect 191741 132832 193660 132834
rect 191741 132776 191746 132832
rect 191802 132776 193660 132832
rect 191741 132774 193660 132776
rect 224940 132832 226951 132834
rect 224940 132776 226890 132832
rect 226946 132776 226951 132832
rect 224940 132774 226951 132776
rect 67725 132771 67791 132774
rect 191741 132771 191807 132774
rect 226885 132771 226951 132774
rect 96613 132290 96679 132293
rect 94668 132288 96679 132290
rect 94668 132232 96618 132288
rect 96674 132232 96679 132288
rect 94668 132230 96679 132232
rect 96613 132227 96679 132230
rect 66897 132018 66963 132021
rect 192937 132018 193003 132021
rect 226701 132018 226767 132021
rect 66897 132016 68908 132018
rect 66897 131960 66902 132016
rect 66958 131960 68908 132016
rect 66897 131958 68908 131960
rect 192937 132016 193660 132018
rect 192937 131960 192942 132016
rect 192998 131960 193660 132016
rect 192937 131958 193660 131960
rect 224940 132016 226767 132018
rect 224940 131960 226706 132016
rect 226762 131960 226767 132016
rect 224940 131958 226767 131960
rect 66897 131955 66963 131958
rect 192937 131955 193003 131958
rect 226701 131955 226767 131958
rect 224350 131684 224356 131748
rect 224420 131746 224426 131748
rect 276013 131746 276079 131749
rect 224420 131744 276079 131746
rect 224420 131688 276018 131744
rect 276074 131688 276079 131744
rect 224420 131686 276079 131688
rect 224420 131684 224426 131686
rect 276013 131683 276079 131686
rect 97349 131474 97415 131477
rect 94668 131472 97415 131474
rect 94668 131416 97354 131472
rect 97410 131416 97415 131472
rect 94668 131414 97415 131416
rect 97349 131411 97415 131414
rect 66345 131202 66411 131205
rect 184197 131202 184263 131205
rect 66345 131200 68908 131202
rect 66345 131144 66350 131200
rect 66406 131144 68908 131200
rect 66345 131142 68908 131144
rect 184197 131200 193660 131202
rect 184197 131144 184202 131200
rect 184258 131144 193660 131200
rect 184197 131142 193660 131144
rect 66345 131139 66411 131142
rect 184197 131139 184263 131142
rect 96613 130930 96679 130933
rect 225413 130930 225479 130933
rect 94668 130928 96679 130930
rect 94668 130872 96618 130928
rect 96674 130872 96679 130928
rect 94668 130870 96679 130872
rect 224940 130928 225479 130930
rect 224940 130872 225418 130928
rect 225474 130872 225479 130928
rect 224940 130870 225479 130872
rect 96613 130867 96679 130870
rect 225413 130867 225479 130870
rect 65885 130658 65951 130661
rect 65885 130656 68908 130658
rect 65885 130600 65890 130656
rect 65946 130600 68908 130656
rect 65885 130598 68908 130600
rect 65885 130595 65951 130598
rect 96613 130114 96679 130117
rect 94668 130112 96679 130114
rect 94668 130056 96618 130112
rect 96674 130056 96679 130112
rect 94668 130054 96679 130056
rect 96613 130051 96679 130054
rect 191005 130114 191071 130117
rect 226609 130114 226675 130117
rect 191005 130112 193660 130114
rect 191005 130056 191010 130112
rect 191066 130056 193660 130112
rect 191005 130054 193660 130056
rect 224940 130112 226675 130114
rect 224940 130056 226614 130112
rect 226670 130056 226675 130112
rect 224940 130054 226675 130056
rect 191005 130051 191071 130054
rect 226609 130051 226675 130054
rect 67541 129842 67607 129845
rect 185485 129842 185551 129845
rect 190269 129842 190335 129845
rect 67541 129840 68908 129842
rect 67541 129784 67546 129840
rect 67602 129784 68908 129840
rect 67541 129782 68908 129784
rect 185485 129840 190335 129842
rect 185485 129784 185490 129840
rect 185546 129784 190274 129840
rect 190330 129784 190335 129840
rect 185485 129782 190335 129784
rect 67541 129779 67607 129782
rect 185485 129779 185551 129782
rect 190269 129779 190335 129782
rect 98494 129298 98500 129300
rect 94668 129238 98500 129298
rect 98494 129236 98500 129238
rect 98564 129236 98570 129300
rect 191189 129298 191255 129301
rect 227161 129298 227227 129301
rect 191189 129296 193660 129298
rect 191189 129240 191194 129296
rect 191250 129240 193660 129296
rect 191189 129238 193660 129240
rect 224940 129296 227227 129298
rect 224940 129240 227166 129296
rect 227222 129240 227227 129296
rect 224940 129238 227227 129240
rect 191189 129235 191255 129238
rect 227161 129235 227227 129238
rect 67725 129026 67791 129029
rect 225045 129026 225111 129029
rect 67725 129024 68908 129026
rect 67725 128968 67730 129024
rect 67786 128968 68908 129024
rect 67725 128966 68908 128968
rect 224910 129024 225111 129026
rect 224910 128968 225050 129024
rect 225106 128968 225111 129024
rect 224910 128966 225111 128968
rect 67725 128963 67791 128966
rect 67541 128890 67607 128893
rect 68134 128890 68140 128892
rect 67541 128888 68140 128890
rect 67541 128832 67546 128888
rect 67602 128832 68140 128888
rect 67541 128830 68140 128832
rect 67541 128827 67607 128830
rect 68134 128828 68140 128830
rect 68204 128828 68210 128892
rect 160921 128482 160987 128485
rect 94668 128480 160987 128482
rect 94668 128424 160926 128480
rect 160982 128424 160987 128480
rect 94668 128422 160987 128424
rect 160921 128419 160987 128422
rect 191189 128482 191255 128485
rect 224910 128482 224970 128966
rect 225045 128963 225111 128966
rect 226149 128482 226215 128485
rect 191189 128480 193660 128482
rect 191189 128424 191194 128480
rect 191250 128424 193660 128480
rect 224910 128480 226215 128482
rect 224910 128452 226154 128480
rect 191189 128422 193660 128424
rect 224940 128424 226154 128452
rect 226210 128424 226215 128480
rect 224940 128422 226215 128424
rect 191189 128419 191255 128422
rect 226149 128419 226215 128422
rect 67909 128210 67975 128213
rect 67909 128208 68908 128210
rect 67909 128152 67914 128208
rect 67970 128152 68908 128208
rect 67909 128150 68908 128152
rect 67909 128147 67975 128150
rect 66897 127666 66963 127669
rect 96705 127666 96771 127669
rect 66897 127664 68908 127666
rect 66897 127608 66902 127664
rect 66958 127608 68908 127664
rect 66897 127606 68908 127608
rect 94668 127664 96771 127666
rect 94668 127608 96710 127664
rect 96766 127608 96771 127664
rect 94668 127606 96771 127608
rect 66897 127603 66963 127606
rect 96705 127603 96771 127606
rect 191741 127666 191807 127669
rect 192334 127666 192340 127668
rect 191741 127664 192340 127666
rect 191741 127608 191746 127664
rect 191802 127608 192340 127664
rect 191741 127606 192340 127608
rect 191741 127603 191807 127606
rect 192334 127604 192340 127606
rect 192404 127666 192410 127668
rect 192404 127606 193660 127666
rect 192404 127604 192410 127606
rect 226609 127394 226675 127397
rect 224940 127392 226675 127394
rect 224940 127336 226614 127392
rect 226670 127336 226675 127392
rect 224940 127334 226675 127336
rect 226609 127331 226675 127334
rect 97533 127122 97599 127125
rect 94668 127120 97599 127122
rect 94668 127064 97538 127120
rect 97594 127064 97599 127120
rect 94668 127062 97599 127064
rect 97533 127059 97599 127062
rect 66805 126850 66871 126853
rect 66805 126848 68908 126850
rect 66805 126792 66810 126848
rect 66866 126792 68908 126848
rect 66805 126790 68908 126792
rect 66805 126787 66871 126790
rect 191557 126578 191623 126581
rect 226885 126578 226951 126581
rect 191557 126576 193660 126578
rect 191557 126520 191562 126576
rect 191618 126520 193660 126576
rect 191557 126518 193660 126520
rect 224940 126576 226951 126578
rect 224940 126520 226890 126576
rect 226946 126520 226951 126576
rect 224940 126518 226951 126520
rect 191557 126515 191623 126518
rect 226885 126515 226951 126518
rect 97809 126306 97875 126309
rect 94668 126304 97875 126306
rect 94668 126248 97814 126304
rect 97870 126248 97875 126304
rect 94668 126246 97875 126248
rect 97809 126243 97875 126246
rect 66713 126034 66779 126037
rect 582373 126034 582439 126037
rect 583520 126034 584960 126124
rect 66713 126032 68908 126034
rect 66713 125976 66718 126032
rect 66774 125976 68908 126032
rect 66713 125974 68908 125976
rect 582373 126032 584960 126034
rect 582373 125976 582378 126032
rect 582434 125976 584960 126032
rect 582373 125974 584960 125976
rect 66713 125971 66779 125974
rect 582373 125971 582439 125974
rect 583520 125884 584960 125974
rect 191046 125700 191052 125764
rect 191116 125762 191122 125764
rect 193254 125762 193260 125764
rect 191116 125702 193260 125762
rect 191116 125700 191122 125702
rect 193254 125700 193260 125702
rect 193324 125762 193330 125764
rect 226425 125762 226491 125765
rect 193324 125702 193660 125762
rect 224940 125760 226491 125762
rect 224940 125704 226430 125760
rect 226486 125704 226491 125760
rect 224940 125702 226491 125704
rect 193324 125700 193330 125702
rect 226425 125699 226491 125702
rect 97942 125490 97948 125492
rect 94668 125430 97948 125490
rect 97942 125428 97948 125430
rect 98012 125490 98018 125492
rect 98453 125490 98519 125493
rect 98012 125488 98519 125490
rect 98012 125432 98458 125488
rect 98514 125432 98519 125488
rect 98012 125430 98519 125432
rect 98012 125428 98018 125430
rect 98453 125427 98519 125430
rect 67541 125218 67607 125221
rect 67541 125216 68908 125218
rect 67541 125160 67546 125216
rect 67602 125160 68908 125216
rect 67541 125158 68908 125160
rect 67541 125155 67607 125158
rect 69422 124884 69428 124948
rect 69492 124884 69498 124948
rect 193121 124946 193187 124949
rect 193121 124944 193660 124946
rect 193121 124888 193126 124944
rect 193182 124888 193660 124944
rect 193121 124886 193660 124888
rect 69430 124372 69490 124884
rect 193121 124883 193187 124886
rect 97073 124674 97139 124677
rect 226609 124674 226675 124677
rect 94668 124672 97139 124674
rect 94668 124616 97078 124672
rect 97134 124616 97139 124672
rect 94668 124614 97139 124616
rect 224940 124672 226675 124674
rect 224940 124616 226614 124672
rect 226670 124616 226675 124672
rect 224940 124614 226675 124616
rect 97073 124611 97139 124614
rect 226609 124611 226675 124614
rect 97809 124130 97875 124133
rect 94668 124128 97875 124130
rect 94668 124072 97814 124128
rect 97870 124072 97875 124128
rect 94668 124070 97875 124072
rect 97809 124067 97875 124070
rect 66253 123858 66319 123861
rect 191465 123858 191531 123861
rect 226517 123858 226583 123861
rect 66253 123856 68908 123858
rect -960 123572 480 123812
rect 66253 123800 66258 123856
rect 66314 123800 68908 123856
rect 66253 123798 68908 123800
rect 191465 123856 193660 123858
rect 191465 123800 191470 123856
rect 191526 123800 193660 123856
rect 191465 123798 193660 123800
rect 224940 123856 226583 123858
rect 224940 123800 226522 123856
rect 226578 123800 226583 123856
rect 224940 123798 226583 123800
rect 66253 123795 66319 123798
rect 191465 123795 191531 123798
rect 226517 123795 226583 123798
rect 97165 123314 97231 123317
rect 94668 123312 97231 123314
rect 94668 123256 97170 123312
rect 97226 123256 97231 123312
rect 94668 123254 97231 123256
rect 97165 123251 97231 123254
rect 66621 123042 66687 123045
rect 191005 123042 191071 123045
rect 226701 123042 226767 123045
rect 66621 123040 68908 123042
rect 66621 122984 66626 123040
rect 66682 122984 68908 123040
rect 66621 122982 68908 122984
rect 191005 123040 193660 123042
rect 191005 122984 191010 123040
rect 191066 122984 193660 123040
rect 191005 122982 193660 122984
rect 224940 123040 226767 123042
rect 224940 122984 226706 123040
rect 226762 122984 226767 123040
rect 224940 122982 226767 122984
rect 66621 122979 66687 122982
rect 191005 122979 191071 122982
rect 226701 122979 226767 122982
rect 97257 122498 97323 122501
rect 94668 122496 97323 122498
rect 94668 122440 97262 122496
rect 97318 122440 97323 122496
rect 94668 122438 97323 122440
rect 97257 122435 97323 122438
rect 65977 122226 66043 122229
rect 191741 122226 191807 122229
rect 226517 122226 226583 122229
rect 65977 122224 68908 122226
rect 65977 122168 65982 122224
rect 66038 122168 68908 122224
rect 65977 122166 68908 122168
rect 191741 122224 193660 122226
rect 191741 122168 191746 122224
rect 191802 122168 193660 122224
rect 191741 122166 193660 122168
rect 224940 122224 226583 122226
rect 224940 122168 226522 122224
rect 226578 122168 226583 122224
rect 224940 122166 226583 122168
rect 65977 122163 66043 122166
rect 191741 122163 191807 122166
rect 226517 122163 226583 122166
rect 97533 121682 97599 121685
rect 94668 121680 97599 121682
rect 94668 121624 97538 121680
rect 97594 121624 97599 121680
rect 94668 121622 97599 121624
rect 97533 121619 97599 121622
rect 66805 121410 66871 121413
rect 191741 121410 191807 121413
rect 66805 121408 68908 121410
rect 66805 121352 66810 121408
rect 66866 121352 68908 121408
rect 66805 121350 68908 121352
rect 191741 121408 193660 121410
rect 191741 121352 191746 121408
rect 191802 121352 193660 121408
rect 191741 121350 193660 121352
rect 66805 121347 66871 121350
rect 191741 121347 191807 121350
rect 224902 121348 224908 121412
rect 224972 121348 224978 121412
rect 224910 121108 224970 121348
rect 96981 120866 97047 120869
rect 94668 120864 97047 120866
rect 94668 120808 96986 120864
rect 97042 120808 97047 120864
rect 94668 120806 97047 120808
rect 96981 120803 97047 120806
rect 66897 120594 66963 120597
rect 66897 120592 68908 120594
rect 66897 120536 66902 120592
rect 66958 120536 68908 120592
rect 66897 120534 68908 120536
rect 66897 120531 66963 120534
rect 95325 120322 95391 120325
rect 96061 120322 96127 120325
rect 94668 120320 96127 120322
rect 94668 120264 95330 120320
rect 95386 120264 96066 120320
rect 96122 120264 96127 120320
rect 94668 120262 96127 120264
rect 95325 120259 95391 120262
rect 96061 120259 96127 120262
rect 191741 120322 191807 120325
rect 226701 120322 226767 120325
rect 191741 120320 193660 120322
rect 191741 120264 191746 120320
rect 191802 120264 193660 120320
rect 191741 120262 193660 120264
rect 224940 120320 226767 120322
rect 224940 120264 226706 120320
rect 226762 120264 226767 120320
rect 224940 120262 226767 120264
rect 191741 120259 191807 120262
rect 226701 120259 226767 120262
rect 66805 120050 66871 120053
rect 66805 120048 68908 120050
rect 66805 119992 66810 120048
rect 66866 119992 68908 120048
rect 66805 119990 68908 119992
rect 66805 119987 66871 119990
rect 97901 119506 97967 119509
rect 94668 119504 97967 119506
rect 94668 119448 97906 119504
rect 97962 119448 97967 119504
rect 94668 119446 97967 119448
rect 97901 119443 97967 119446
rect 191741 119506 191807 119509
rect 226374 119506 226380 119508
rect 191741 119504 193660 119506
rect 191741 119448 191746 119504
rect 191802 119448 193660 119504
rect 191741 119446 193660 119448
rect 224940 119446 226380 119506
rect 191741 119443 191807 119446
rect 226374 119444 226380 119446
rect 226444 119444 226450 119508
rect 66897 119234 66963 119237
rect 66897 119232 68908 119234
rect 66897 119176 66902 119232
rect 66958 119176 68908 119232
rect 66897 119174 68908 119176
rect 66897 119171 66963 119174
rect 97901 118690 97967 118693
rect 94668 118688 97967 118690
rect 94668 118632 97906 118688
rect 97962 118632 97967 118688
rect 94668 118630 97967 118632
rect 97901 118627 97967 118630
rect 190545 118690 190611 118693
rect 191005 118690 191071 118693
rect 190545 118688 193660 118690
rect 190545 118632 190550 118688
rect 190606 118632 191010 118688
rect 191066 118632 193660 118688
rect 190545 118630 193660 118632
rect 190545 118627 190611 118630
rect 191005 118627 191071 118630
rect 65926 118356 65932 118420
rect 65996 118418 66002 118420
rect 226701 118418 226767 118421
rect 65996 118358 68908 118418
rect 224940 118416 226767 118418
rect 224940 118360 226706 118416
rect 226762 118360 226767 118416
rect 224940 118358 226767 118360
rect 65996 118356 66002 118358
rect 226701 118355 226767 118358
rect 66713 117602 66779 117605
rect 66713 117600 68908 117602
rect 66713 117544 66718 117600
rect 66774 117544 68908 117600
rect 66713 117542 68908 117544
rect 66713 117539 66779 117542
rect 94638 117330 94698 117844
rect 191649 117602 191715 117605
rect 226609 117602 226675 117605
rect 191649 117600 193660 117602
rect 191649 117544 191654 117600
rect 191710 117544 193660 117600
rect 191649 117542 193660 117544
rect 224940 117600 226675 117602
rect 224940 117544 226614 117600
rect 226670 117544 226675 117600
rect 224940 117542 226675 117544
rect 191649 117539 191715 117542
rect 226609 117539 226675 117542
rect 116669 117330 116735 117333
rect 94638 117328 116735 117330
rect 94638 117272 116674 117328
rect 116730 117272 116735 117328
rect 94638 117270 116735 117272
rect 116669 117267 116735 117270
rect 66805 117058 66871 117061
rect 97349 117058 97415 117061
rect 66805 117056 68908 117058
rect 66805 117000 66810 117056
rect 66866 117000 68908 117056
rect 66805 116998 68908 117000
rect 94668 117056 97415 117058
rect 94668 117000 97354 117056
rect 97410 117000 97415 117056
rect 94668 116998 97415 117000
rect 66805 116995 66871 116998
rect 97349 116995 97415 116998
rect 191741 116786 191807 116789
rect 225229 116786 225295 116789
rect 191741 116784 193660 116786
rect 191741 116728 191746 116784
rect 191802 116728 193660 116784
rect 191741 116726 193660 116728
rect 224940 116784 225295 116786
rect 224940 116728 225234 116784
rect 225290 116728 225295 116784
rect 224940 116726 225295 116728
rect 191741 116723 191807 116726
rect 225229 116723 225295 116726
rect 97901 116514 97967 116517
rect 94668 116512 97967 116514
rect 94668 116456 97906 116512
rect 97962 116456 97967 116512
rect 94668 116454 97967 116456
rect 97901 116451 97967 116454
rect 66253 116242 66319 116245
rect 66253 116240 68908 116242
rect 66253 116184 66258 116240
rect 66314 116184 68908 116240
rect 66253 116182 68908 116184
rect 66253 116179 66319 116182
rect 191005 115970 191071 115973
rect 226701 115970 226767 115973
rect 191005 115968 193660 115970
rect 191005 115912 191010 115968
rect 191066 115912 193660 115968
rect 191005 115910 193660 115912
rect 224940 115968 226767 115970
rect 224940 115912 226706 115968
rect 226762 115912 226767 115968
rect 224940 115910 226767 115912
rect 191005 115907 191071 115910
rect 226701 115907 226767 115910
rect 97901 115698 97967 115701
rect 94668 115696 97967 115698
rect 94668 115640 97906 115696
rect 97962 115640 97967 115696
rect 94668 115638 97967 115640
rect 97901 115635 97967 115638
rect 66897 115426 66963 115429
rect 66897 115424 68908 115426
rect 66897 115368 66902 115424
rect 66958 115368 68908 115424
rect 66897 115366 68908 115368
rect 66897 115363 66963 115366
rect 190821 115154 190887 115157
rect 190821 115152 193660 115154
rect 190821 115096 190826 115152
rect 190882 115096 193660 115152
rect 190821 115094 193660 115096
rect 190821 115091 190887 115094
rect 97809 114882 97875 114885
rect 226701 114882 226767 114885
rect 94668 114880 97875 114882
rect 94668 114824 97814 114880
rect 97870 114824 97875 114880
rect 94668 114822 97875 114824
rect 224940 114880 226767 114882
rect 224940 114824 226706 114880
rect 226762 114824 226767 114880
rect 224940 114822 226767 114824
rect 97809 114819 97875 114822
rect 226701 114819 226767 114822
rect 66805 114610 66871 114613
rect 66805 114608 68908 114610
rect 66805 114552 66810 114608
rect 66866 114552 68908 114608
rect 66805 114550 68908 114552
rect 66805 114547 66871 114550
rect 97809 114066 97875 114069
rect 94668 114064 97875 114066
rect 94668 114008 97814 114064
rect 97870 114008 97875 114064
rect 94668 114006 97875 114008
rect 97809 114003 97875 114006
rect 191833 114066 191899 114069
rect 226609 114066 226675 114069
rect 191833 114064 193660 114066
rect 191833 114008 191838 114064
rect 191894 114008 193660 114064
rect 191833 114006 193660 114008
rect 224940 114064 226675 114066
rect 224940 114008 226614 114064
rect 226670 114008 226675 114064
rect 224940 114006 226675 114008
rect 191833 114003 191899 114006
rect 226609 114003 226675 114006
rect 66805 113794 66871 113797
rect 225045 113794 225111 113797
rect 66805 113792 68908 113794
rect 66805 113736 66810 113792
rect 66866 113736 68908 113792
rect 66805 113734 68908 113736
rect 224910 113792 225111 113794
rect 224910 113736 225050 113792
rect 225106 113736 225111 113792
rect 224910 113734 225111 113736
rect 66805 113731 66871 113734
rect 97901 113522 97967 113525
rect 94668 113520 97967 113522
rect 94668 113464 97906 113520
rect 97962 113464 97967 113520
rect 94668 113462 97967 113464
rect 97901 113459 97967 113462
rect 66897 113250 66963 113253
rect 191741 113250 191807 113253
rect 66897 113248 68908 113250
rect 66897 113192 66902 113248
rect 66958 113192 68908 113248
rect 66897 113190 68908 113192
rect 191741 113248 193660 113250
rect 191741 113192 191746 113248
rect 191802 113192 193660 113248
rect 224910 113220 224970 113734
rect 225045 113731 225111 113734
rect 191741 113190 193660 113192
rect 66897 113187 66963 113190
rect 191741 113187 191807 113190
rect 582833 112842 582899 112845
rect 583520 112842 584960 112932
rect 582833 112840 584960 112842
rect 582833 112784 582838 112840
rect 582894 112784 584960 112840
rect 582833 112782 584960 112784
rect 582833 112779 582899 112782
rect 583520 112692 584960 112782
rect 67817 112434 67883 112437
rect 67817 112432 68908 112434
rect 67817 112376 67822 112432
rect 67878 112376 68908 112432
rect 67817 112374 68908 112376
rect 67817 112371 67883 112374
rect 94638 112162 94698 112676
rect 191741 112434 191807 112437
rect 191741 112432 193660 112434
rect 191741 112376 191746 112432
rect 191802 112376 193660 112432
rect 191741 112374 193660 112376
rect 191741 112371 191807 112374
rect 178769 112162 178835 112165
rect 226701 112162 226767 112165
rect 94638 112160 178835 112162
rect 94638 112104 178774 112160
rect 178830 112104 178835 112160
rect 94638 112102 178835 112104
rect 224940 112160 226767 112162
rect 224940 112104 226706 112160
rect 226762 112104 226767 112160
rect 224940 112102 226767 112104
rect 178769 112099 178835 112102
rect 226701 112099 226767 112102
rect 97073 111890 97139 111893
rect 94668 111888 97139 111890
rect 94668 111832 97078 111888
rect 97134 111832 97139 111888
rect 94668 111830 97139 111832
rect 97073 111827 97139 111830
rect 66805 111618 66871 111621
rect 66805 111616 68908 111618
rect 66805 111560 66810 111616
rect 66866 111560 68908 111616
rect 66805 111558 68908 111560
rect 66805 111555 66871 111558
rect 96705 111074 96771 111077
rect 94668 111072 96771 111074
rect 94668 111016 96710 111072
rect 96766 111016 96771 111072
rect 94668 111014 96771 111016
rect 96705 111011 96771 111014
rect 66805 110802 66871 110805
rect 189073 110802 189139 110805
rect 193630 110802 193690 111316
rect 66805 110800 68908 110802
rect -960 110666 480 110756
rect 66805 110744 66810 110800
rect 66866 110744 68908 110800
rect 66805 110742 68908 110744
rect 189073 110800 193690 110802
rect 189073 110744 189078 110800
rect 189134 110744 193690 110800
rect 189073 110742 193690 110744
rect 224910 110802 224970 111316
rect 227713 110802 227779 110805
rect 224910 110800 227779 110802
rect 224910 110744 227718 110800
rect 227774 110744 227779 110800
rect 224910 110742 227779 110744
rect 66805 110739 66871 110742
rect 189073 110739 189139 110742
rect 227713 110739 227779 110742
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 191741 110530 191807 110533
rect 227069 110530 227135 110533
rect 191741 110528 193660 110530
rect 191741 110472 191746 110528
rect 191802 110472 193660 110528
rect 191741 110470 193660 110472
rect 224940 110528 227135 110530
rect 224940 110472 227074 110528
rect 227130 110472 227135 110528
rect 224940 110470 227135 110472
rect 191741 110467 191807 110470
rect 227069 110467 227135 110470
rect 66805 110258 66871 110261
rect 97901 110258 97967 110261
rect 66805 110256 68908 110258
rect 66805 110200 66810 110256
rect 66866 110200 68908 110256
rect 66805 110198 68908 110200
rect 94668 110256 97967 110258
rect 94668 110200 97906 110256
rect 97962 110200 97967 110256
rect 94668 110198 97967 110200
rect 66805 110195 66871 110198
rect 97901 110195 97967 110198
rect 97809 109714 97875 109717
rect 94668 109712 97875 109714
rect 94668 109656 97814 109712
rect 97870 109656 97875 109712
rect 94668 109654 97875 109656
rect 97809 109651 97875 109654
rect 191097 109714 191163 109717
rect 225137 109714 225203 109717
rect 191097 109712 193660 109714
rect 191097 109656 191102 109712
rect 191158 109656 193660 109712
rect 191097 109654 193660 109656
rect 224940 109712 225203 109714
rect 224940 109656 225142 109712
rect 225198 109656 225203 109712
rect 224940 109654 225203 109656
rect 191097 109651 191163 109654
rect 225137 109651 225203 109654
rect 67541 109442 67607 109445
rect 67541 109440 68908 109442
rect 67541 109384 67546 109440
rect 67602 109384 68908 109440
rect 67541 109382 68908 109384
rect 67541 109379 67607 109382
rect 107469 109034 107535 109037
rect 114553 109034 114619 109037
rect 115289 109034 115355 109037
rect 107469 109032 115355 109034
rect 107469 108976 107474 109032
rect 107530 108976 114558 109032
rect 114614 108976 115294 109032
rect 115350 108976 115355 109032
rect 107469 108974 115355 108976
rect 107469 108971 107535 108974
rect 114553 108971 114619 108974
rect 115289 108971 115355 108974
rect 98085 108898 98151 108901
rect 94668 108896 98151 108898
rect 94668 108840 98090 108896
rect 98146 108840 98151 108896
rect 94668 108838 98151 108840
rect 98085 108835 98151 108838
rect 65977 108626 66043 108629
rect 65977 108624 68908 108626
rect 65977 108568 65982 108624
rect 66038 108568 68908 108624
rect 65977 108566 68908 108568
rect 65977 108563 66043 108566
rect 192017 108354 192083 108357
rect 193630 108354 193690 108868
rect 226425 108626 226491 108629
rect 224940 108624 226491 108626
rect 224940 108596 226430 108624
rect 192017 108352 193690 108354
rect 192017 108296 192022 108352
rect 192078 108296 193690 108352
rect 192017 108294 193690 108296
rect 224910 108568 226430 108596
rect 226486 108568 226491 108624
rect 224910 108566 226491 108568
rect 192017 108291 192083 108294
rect 184749 108218 184815 108221
rect 186313 108218 186379 108221
rect 184749 108216 186379 108218
rect 184749 108160 184754 108216
rect 184810 108160 186318 108216
rect 186374 108160 186379 108216
rect 184749 108158 186379 108160
rect 184749 108155 184815 108158
rect 186313 108155 186379 108158
rect 97901 108082 97967 108085
rect 224910 108084 224970 108566
rect 226425 108563 226491 108566
rect 94668 108080 97967 108082
rect 94668 108024 97906 108080
rect 97962 108024 97967 108080
rect 94668 108022 97967 108024
rect 97901 108019 97967 108022
rect 224902 108020 224908 108084
rect 224972 108020 224978 108084
rect 66805 107810 66871 107813
rect 186313 107810 186379 107813
rect 226701 107810 226767 107813
rect 66805 107808 68908 107810
rect 66805 107752 66810 107808
rect 66866 107752 68908 107808
rect 66805 107750 68908 107752
rect 186313 107808 193660 107810
rect 186313 107752 186318 107808
rect 186374 107752 193660 107808
rect 186313 107750 193660 107752
rect 224940 107808 226767 107810
rect 224940 107752 226706 107808
rect 226762 107752 226767 107808
rect 224940 107750 226767 107752
rect 66805 107747 66871 107750
rect 186313 107747 186379 107750
rect 226701 107747 226767 107750
rect 179229 107674 179295 107677
rect 192017 107674 192083 107677
rect 179229 107672 192083 107674
rect 179229 107616 179234 107672
rect 179290 107616 192022 107672
rect 192078 107616 192083 107672
rect 179229 107614 192083 107616
rect 179229 107611 179295 107614
rect 192017 107611 192083 107614
rect 96705 107266 96771 107269
rect 94668 107264 96771 107266
rect 94668 107208 96710 107264
rect 96766 107208 96771 107264
rect 94668 107206 96771 107208
rect 96705 107203 96771 107206
rect 66805 106994 66871 106997
rect 191741 106994 191807 106997
rect 226793 106994 226859 106997
rect 66805 106992 68908 106994
rect 66805 106936 66810 106992
rect 66866 106936 68908 106992
rect 66805 106934 68908 106936
rect 191741 106992 193660 106994
rect 191741 106936 191746 106992
rect 191802 106936 193660 106992
rect 191741 106934 193660 106936
rect 224940 106992 226859 106994
rect 224940 106936 226798 106992
rect 226854 106936 226859 106992
rect 224940 106934 226859 106936
rect 66805 106931 66871 106934
rect 191741 106931 191807 106934
rect 226793 106931 226859 106934
rect 66110 106388 66116 106452
rect 66180 106450 66186 106452
rect 66180 106390 68908 106450
rect 66180 106388 66186 106390
rect 94638 106314 94698 106692
rect 177389 106314 177455 106317
rect 94638 106312 177455 106314
rect 94638 106256 177394 106312
rect 177450 106256 177455 106312
rect 94638 106254 177455 106256
rect 177389 106251 177455 106254
rect 191189 106178 191255 106181
rect 191189 106176 193660 106178
rect 191189 106120 191194 106176
rect 191250 106120 193660 106176
rect 191189 106118 193660 106120
rect 191189 106115 191255 106118
rect 100702 105906 100708 105908
rect 94668 105846 100708 105906
rect 100702 105844 100708 105846
rect 100772 105844 100778 105908
rect 226701 105906 226767 105909
rect 224940 105904 226767 105906
rect 224940 105848 226706 105904
rect 226762 105848 226767 105904
rect 224940 105846 226767 105848
rect 226701 105843 226767 105846
rect 66529 105634 66595 105637
rect 66529 105632 68908 105634
rect 66529 105576 66534 105632
rect 66590 105576 68908 105632
rect 66529 105574 68908 105576
rect 66529 105571 66595 105574
rect 95969 105090 96035 105093
rect 94668 105088 96035 105090
rect 94668 105032 95974 105088
rect 96030 105032 96035 105088
rect 94668 105030 96035 105032
rect 95969 105027 96035 105030
rect 191741 105090 191807 105093
rect 226425 105090 226491 105093
rect 191741 105088 193660 105090
rect 191741 105032 191746 105088
rect 191802 105032 193660 105088
rect 191741 105030 193660 105032
rect 224940 105088 226491 105090
rect 224940 105032 226430 105088
rect 226486 105032 226491 105088
rect 224940 105030 226491 105032
rect 191741 105027 191807 105030
rect 226425 105027 226491 105030
rect 66805 104818 66871 104821
rect 66805 104816 68908 104818
rect 66805 104760 66810 104816
rect 66866 104760 68908 104816
rect 66805 104758 68908 104760
rect 66805 104755 66871 104758
rect 193806 104484 193812 104548
rect 193876 104484 193882 104548
rect 96797 104274 96863 104277
rect 94668 104272 96863 104274
rect 94668 104216 96802 104272
rect 96858 104216 96863 104272
rect 94668 104214 96863 104216
rect 96797 104211 96863 104214
rect 192477 104274 192543 104277
rect 193814 104274 193874 104484
rect 226701 104274 226767 104277
rect 192477 104272 193874 104274
rect 192477 104216 192482 104272
rect 192538 104244 193874 104272
rect 224940 104272 226767 104274
rect 192538 104216 193844 104244
rect 192477 104214 193844 104216
rect 224940 104216 226706 104272
rect 226762 104216 226767 104272
rect 224940 104214 226767 104216
rect 192477 104211 192543 104214
rect 226701 104211 226767 104214
rect 193213 104138 193279 104141
rect 194174 104138 194180 104140
rect 193213 104136 194180 104138
rect 193213 104080 193218 104136
rect 193274 104080 194180 104136
rect 193213 104078 194180 104080
rect 193213 104075 193279 104078
rect 194174 104076 194180 104078
rect 194244 104076 194250 104140
rect 67357 104002 67423 104005
rect 67357 104000 68908 104002
rect 67357 103944 67362 104000
rect 67418 103944 68908 104000
rect 67357 103942 68908 103944
rect 67357 103939 67423 103942
rect 95141 103594 95207 103597
rect 95141 103592 95250 103594
rect 95141 103536 95146 103592
rect 95202 103536 95250 103592
rect 95141 103531 95250 103536
rect 95190 103458 95250 103531
rect 96521 103458 96587 103461
rect 94668 103456 96587 103458
rect 94668 103400 96526 103456
rect 96582 103400 96587 103456
rect 94668 103398 96587 103400
rect 96521 103395 96587 103398
rect 191741 103458 191807 103461
rect 226609 103458 226675 103461
rect 191741 103456 193660 103458
rect 191741 103400 191746 103456
rect 191802 103400 193660 103456
rect 191741 103398 193660 103400
rect 224940 103456 226675 103458
rect 224940 103400 226614 103456
rect 226670 103400 226675 103456
rect 224940 103398 226675 103400
rect 191741 103395 191807 103398
rect 226609 103395 226675 103398
rect 66805 103186 66871 103189
rect 66805 103184 68908 103186
rect 66805 103128 66810 103184
rect 66866 103128 68908 103184
rect 66805 103126 68908 103128
rect 66805 103123 66871 103126
rect 97901 102914 97967 102917
rect 94668 102912 97967 102914
rect 94668 102856 97906 102912
rect 97962 102856 97967 102912
rect 94668 102854 97967 102856
rect 97901 102851 97967 102854
rect 66069 102642 66135 102645
rect 193029 102642 193095 102645
rect 66069 102640 68908 102642
rect 66069 102584 66074 102640
rect 66130 102584 68908 102640
rect 66069 102582 68908 102584
rect 193029 102640 193660 102642
rect 193029 102584 193034 102640
rect 193090 102584 193660 102640
rect 193029 102582 193660 102584
rect 66069 102579 66135 102582
rect 193029 102579 193095 102582
rect 226701 102370 226767 102373
rect 224940 102368 226767 102370
rect 224940 102312 226706 102368
rect 226762 102312 226767 102368
rect 224940 102310 226767 102312
rect 226701 102307 226767 102310
rect 97901 102098 97967 102101
rect 94668 102096 97967 102098
rect 94668 102040 97906 102096
rect 97962 102040 97967 102096
rect 94668 102038 97967 102040
rect 97901 102035 97967 102038
rect 66621 101826 66687 101829
rect 66621 101824 68908 101826
rect 66621 101768 66626 101824
rect 66682 101768 68908 101824
rect 66621 101766 68908 101768
rect 66621 101763 66687 101766
rect 191741 101554 191807 101557
rect 226517 101554 226583 101557
rect 191741 101552 193660 101554
rect 191741 101496 191746 101552
rect 191802 101496 193660 101552
rect 191741 101494 193660 101496
rect 224940 101552 226583 101554
rect 224940 101496 226522 101552
rect 226578 101496 226583 101552
rect 224940 101494 226583 101496
rect 191741 101491 191807 101494
rect 226517 101491 226583 101494
rect 99465 101282 99531 101285
rect 94668 101280 99531 101282
rect 94668 101224 99470 101280
rect 99526 101224 99531 101280
rect 94668 101222 99531 101224
rect 99465 101219 99531 101222
rect 67817 101010 67883 101013
rect 67817 101008 68908 101010
rect 67817 100952 67822 101008
rect 67878 100952 68908 101008
rect 67817 100950 68908 100952
rect 67817 100947 67883 100950
rect 191557 100738 191623 100741
rect 226701 100738 226767 100741
rect 191557 100736 193660 100738
rect 191557 100680 191562 100736
rect 191618 100680 193660 100736
rect 191557 100678 193660 100680
rect 224940 100736 226767 100738
rect 224940 100680 226706 100736
rect 226762 100680 226767 100736
rect 224940 100678 226767 100680
rect 191557 100675 191623 100678
rect 226701 100675 226767 100678
rect 97533 100466 97599 100469
rect 94668 100464 97599 100466
rect 94668 100408 97538 100464
rect 97594 100408 97599 100464
rect 94668 100406 97599 100408
rect 97533 100403 97599 100406
rect 67357 100194 67423 100197
rect 67357 100192 68908 100194
rect 67357 100136 67362 100192
rect 67418 100136 68908 100192
rect 67357 100134 68908 100136
rect 67357 100131 67423 100134
rect 100293 100058 100359 100061
rect 120073 100058 120139 100061
rect 191046 100058 191052 100060
rect 100293 100056 191052 100058
rect 100293 100000 100298 100056
rect 100354 100000 120078 100056
rect 120134 100000 191052 100056
rect 100293 99998 191052 100000
rect 100293 99995 100359 99998
rect 120073 99995 120139 99998
rect 191046 99996 191052 99998
rect 191116 99996 191122 100060
rect 191741 99922 191807 99925
rect 191741 99920 193660 99922
rect 191741 99864 191746 99920
rect 191802 99864 193660 99920
rect 191741 99862 193660 99864
rect 191741 99859 191807 99862
rect 66805 99650 66871 99653
rect 97901 99650 97967 99653
rect 226609 99650 226675 99653
rect 66805 99648 68908 99650
rect 66805 99592 66810 99648
rect 66866 99592 68908 99648
rect 66805 99590 68908 99592
rect 94668 99648 97967 99650
rect 94668 99592 97906 99648
rect 97962 99592 97967 99648
rect 94668 99590 97967 99592
rect 224940 99648 226675 99650
rect 224940 99592 226614 99648
rect 226670 99592 226675 99648
rect 224940 99590 226675 99592
rect 66805 99587 66871 99590
rect 97901 99587 97967 99590
rect 226609 99587 226675 99590
rect 582833 99514 582899 99517
rect 583520 99514 584960 99604
rect 582833 99512 584960 99514
rect 582833 99456 582838 99512
rect 582894 99456 584960 99512
rect 582833 99454 584960 99456
rect 582833 99451 582899 99454
rect 583520 99364 584960 99454
rect 97809 99106 97875 99109
rect 94668 99104 97875 99106
rect 94668 99048 97814 99104
rect 97870 99048 97875 99104
rect 94668 99046 97875 99048
rect 97809 99043 97875 99046
rect 66805 98834 66871 98837
rect 226374 98834 226380 98836
rect 66805 98832 68908 98834
rect 66805 98776 66810 98832
rect 66866 98776 68908 98832
rect 66805 98774 68908 98776
rect 66805 98771 66871 98774
rect 94814 98500 94820 98564
rect 94884 98562 94890 98564
rect 193630 98562 193690 98804
rect 224940 98774 226380 98834
rect 226374 98772 226380 98774
rect 226444 98772 226450 98836
rect 94884 98502 193690 98562
rect 94884 98500 94890 98502
rect 97901 98290 97967 98293
rect 94668 98288 97967 98290
rect 94668 98232 97906 98288
rect 97962 98232 97967 98288
rect 94668 98230 97967 98232
rect 97901 98227 97967 98230
rect 66662 97956 66668 98020
rect 66732 98018 66738 98020
rect 190545 98018 190611 98021
rect 227345 98018 227411 98021
rect 227713 98018 227779 98021
rect 66732 97958 68908 98018
rect 190545 98016 193660 98018
rect 190545 97960 190550 98016
rect 190606 97960 193660 98016
rect 190545 97958 193660 97960
rect 224940 98016 227779 98018
rect 224940 97960 227350 98016
rect 227406 97960 227718 98016
rect 227774 97960 227779 98016
rect 224940 97958 227779 97960
rect 66732 97956 66738 97958
rect 190545 97955 190611 97958
rect 227345 97955 227411 97958
rect 227713 97955 227779 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 67449 97202 67515 97205
rect 67449 97200 68908 97202
rect 67449 97144 67454 97200
rect 67510 97144 68908 97200
rect 67449 97142 68908 97144
rect 67449 97139 67515 97142
rect 94638 96930 94698 97444
rect 224534 97412 224540 97476
rect 224604 97474 224610 97476
rect 280153 97474 280219 97477
rect 224604 97472 280219 97474
rect 224604 97416 280158 97472
rect 280214 97416 280219 97472
rect 224604 97414 280219 97416
rect 224604 97412 224610 97414
rect 280153 97411 280219 97414
rect 190453 97202 190519 97205
rect 225229 97202 225295 97205
rect 226241 97202 226307 97205
rect 190453 97200 193660 97202
rect 190453 97144 190458 97200
rect 190514 97144 193660 97200
rect 190453 97142 193660 97144
rect 224940 97200 226307 97202
rect 224940 97144 225234 97200
rect 225290 97144 226246 97200
rect 226302 97144 226307 97200
rect 224940 97142 226307 97144
rect 190453 97139 190519 97142
rect 225229 97139 225295 97142
rect 226241 97139 226307 97142
rect 188061 96930 188127 96933
rect 94638 96928 188127 96930
rect 94638 96872 188066 96928
rect 188122 96872 188127 96928
rect 94638 96870 188127 96872
rect 188061 96867 188127 96870
rect 96705 96658 96771 96661
rect 94668 96656 96771 96658
rect 94668 96600 96710 96656
rect 96766 96600 96771 96656
rect 94668 96598 96771 96600
rect 96705 96595 96771 96598
rect 66437 96386 66503 96389
rect 193213 96386 193279 96389
rect 66437 96384 68908 96386
rect 66437 96328 66442 96384
rect 66498 96328 68908 96384
rect 66437 96326 68908 96328
rect 193213 96384 193660 96386
rect 193213 96328 193218 96384
rect 193274 96328 193660 96384
rect 193213 96326 193660 96328
rect 66437 96323 66503 96326
rect 193213 96323 193279 96326
rect 97901 96114 97967 96117
rect 226701 96114 226767 96117
rect 94668 96112 97967 96114
rect 94668 96056 97906 96112
rect 97962 96056 97967 96112
rect 94668 96054 97967 96056
rect 224940 96112 226767 96114
rect 224940 96056 226706 96112
rect 226762 96056 226767 96112
rect 224940 96054 226767 96056
rect 97901 96051 97967 96054
rect 226701 96051 226767 96054
rect 227805 95842 227871 95845
rect 246297 95842 246363 95845
rect 224910 95840 246363 95842
rect 69430 95300 69490 95812
rect 224910 95784 227810 95840
rect 227866 95784 246302 95840
rect 246358 95784 246363 95840
rect 224910 95782 246363 95784
rect 94814 95508 94820 95572
rect 94884 95570 94890 95572
rect 94884 95510 180810 95570
rect 94884 95508 94890 95510
rect 69422 95236 69428 95300
rect 69492 95236 69498 95300
rect 97073 95298 97139 95301
rect 94668 95296 97139 95298
rect 94668 95240 97078 95296
rect 97134 95240 97139 95296
rect 94668 95238 97139 95240
rect 180750 95298 180810 95510
rect 191373 95434 191439 95437
rect 193213 95434 193279 95437
rect 186270 95432 193279 95434
rect 186270 95376 191378 95432
rect 191434 95376 193218 95432
rect 193274 95376 193279 95432
rect 186270 95374 193279 95376
rect 186270 95298 186330 95374
rect 191373 95371 191439 95374
rect 193213 95371 193279 95374
rect 180750 95238 186330 95298
rect 97073 95235 97139 95238
rect 186814 95236 186820 95300
rect 186884 95298 186890 95300
rect 186884 95238 193660 95298
rect 224910 95268 224970 95782
rect 227805 95779 227871 95782
rect 246297 95779 246363 95782
rect 186884 95236 186890 95238
rect 226333 95162 226399 95165
rect 227529 95162 227595 95165
rect 226333 95160 227595 95162
rect 226333 95104 226338 95160
rect 226394 95104 227534 95160
rect 227590 95104 227595 95160
rect 226333 95102 227595 95104
rect 226333 95099 226399 95102
rect 227529 95099 227595 95102
rect 66805 95026 66871 95029
rect 66805 95024 68908 95026
rect 66805 94968 66810 95024
rect 66866 94968 68908 95024
rect 66805 94966 68908 94968
rect 66805 94963 66871 94966
rect 224718 94692 224724 94756
rect 224788 94754 224794 94756
rect 270493 94754 270559 94757
rect 224788 94752 270559 94754
rect 224788 94696 270498 94752
rect 270554 94696 270559 94752
rect 224788 94694 270559 94696
rect 224788 94692 224794 94694
rect 270493 94691 270559 94694
rect 64781 94482 64847 94485
rect 69238 94482 69244 94484
rect 64781 94480 69244 94482
rect 64781 94424 64786 94480
rect 64842 94424 69244 94480
rect 64781 94422 69244 94424
rect 64781 94419 64847 94422
rect 69238 94420 69244 94422
rect 69308 94420 69314 94484
rect 97809 94482 97875 94485
rect 94668 94480 97875 94482
rect 94668 94424 97814 94480
rect 97870 94424 97875 94480
rect 94668 94422 97875 94424
rect 97809 94419 97875 94422
rect 166441 94482 166507 94485
rect 166901 94482 166967 94485
rect 190177 94482 190243 94485
rect 226333 94482 226399 94485
rect 166441 94480 193660 94482
rect 166441 94424 166446 94480
rect 166502 94424 166906 94480
rect 166962 94424 190182 94480
rect 190238 94424 193660 94480
rect 166441 94422 193660 94424
rect 224940 94480 226399 94482
rect 224940 94424 226338 94480
rect 226394 94424 226399 94480
rect 224940 94422 226399 94424
rect 166441 94419 166507 94422
rect 166901 94419 166967 94422
rect 190177 94419 190243 94422
rect 226333 94419 226399 94422
rect 67909 93938 67975 93941
rect 68878 93938 68938 94180
rect 67909 93936 68938 93938
rect 67909 93880 67914 93936
rect 67970 93880 68938 93936
rect 67909 93878 68938 93880
rect 67909 93875 67975 93878
rect 192334 93740 192340 93804
rect 192404 93802 192410 93804
rect 192845 93802 192911 93805
rect 192404 93800 192911 93802
rect 192404 93744 192850 93800
rect 192906 93744 192911 93800
rect 192404 93742 192911 93744
rect 192404 93740 192410 93742
rect 192845 93739 192911 93742
rect 97901 93666 97967 93669
rect 94668 93664 97967 93666
rect 94668 93608 97906 93664
rect 97962 93608 97967 93664
rect 94668 93606 97967 93608
rect 97901 93603 97967 93606
rect 190453 93666 190519 93669
rect 226885 93666 226951 93669
rect 190453 93664 193660 93666
rect 190453 93608 190458 93664
rect 190514 93608 193660 93664
rect 190453 93606 193660 93608
rect 224940 93664 226951 93666
rect 224940 93608 226890 93664
rect 226946 93608 226951 93664
rect 224940 93606 226951 93608
rect 190453 93603 190519 93606
rect 226885 93603 226951 93606
rect 66989 93394 67055 93397
rect 66989 93392 68908 93394
rect 66989 93336 66994 93392
rect 67050 93336 68908 93392
rect 66989 93334 68908 93336
rect 66989 93331 67055 93334
rect 202086 93332 202092 93396
rect 202156 93394 202162 93396
rect 202229 93394 202295 93397
rect 224769 93396 224835 93397
rect 202156 93392 202295 93394
rect 202156 93336 202234 93392
rect 202290 93336 202295 93392
rect 202156 93334 202295 93336
rect 202156 93332 202162 93334
rect 202229 93331 202295 93334
rect 224718 93332 224724 93396
rect 224788 93394 224835 93396
rect 224788 93392 224880 93394
rect 224830 93336 224880 93392
rect 224788 93334 224880 93336
rect 224788 93332 224835 93334
rect 224769 93331 224835 93332
rect 224493 93258 224559 93261
rect 227662 93258 227668 93260
rect 224493 93256 227668 93258
rect 224493 93200 224498 93256
rect 224554 93200 227668 93256
rect 224493 93198 227668 93200
rect 224493 93195 224559 93198
rect 227662 93196 227668 93198
rect 227732 93196 227738 93260
rect 95877 92986 95943 92989
rect 210417 92988 210483 92989
rect 210366 92986 210372 92988
rect 95877 92984 103530 92986
rect 95877 92928 95882 92984
rect 95938 92928 103530 92984
rect 95877 92926 103530 92928
rect 210326 92926 210372 92986
rect 210436 92984 210483 92988
rect 210478 92928 210483 92984
rect 95877 92923 95943 92926
rect 97206 92850 97212 92852
rect 94668 92790 97212 92850
rect 97206 92788 97212 92790
rect 97276 92788 97282 92852
rect 103470 92850 103530 92926
rect 210366 92924 210372 92926
rect 210436 92924 210483 92928
rect 210417 92923 210483 92924
rect 200297 92850 200363 92853
rect 200614 92850 200620 92852
rect 103470 92848 200620 92850
rect 103470 92792 200302 92848
rect 200358 92792 200620 92848
rect 103470 92790 200620 92792
rect 200297 92787 200363 92790
rect 200614 92788 200620 92790
rect 200684 92850 200690 92852
rect 201033 92850 201099 92853
rect 208393 92852 208459 92853
rect 208342 92850 208348 92852
rect 200684 92848 201099 92850
rect 200684 92792 201038 92848
rect 201094 92792 201099 92848
rect 200684 92790 201099 92792
rect 208302 92790 208348 92850
rect 208412 92848 208459 92852
rect 208454 92792 208459 92848
rect 200684 92788 200690 92790
rect 201033 92787 201099 92790
rect 208342 92788 208348 92790
rect 208412 92788 208459 92792
rect 208393 92787 208459 92788
rect 224033 92850 224099 92853
rect 224534 92850 224540 92852
rect 224033 92848 224540 92850
rect 224033 92792 224038 92848
rect 224094 92792 224540 92848
rect 224033 92790 224540 92792
rect 224033 92787 224099 92790
rect 224534 92788 224540 92790
rect 224604 92788 224610 92852
rect 68870 92652 68876 92716
rect 68940 92714 68946 92716
rect 69703 92714 69769 92717
rect 68940 92712 69769 92714
rect 68940 92656 69708 92712
rect 69764 92656 69769 92712
rect 68940 92654 69769 92656
rect 68940 92652 68946 92654
rect 69703 92651 69769 92654
rect 71175 92714 71241 92717
rect 71446 92714 71452 92716
rect 71175 92712 71452 92714
rect 71175 92656 71180 92712
rect 71236 92656 71452 92712
rect 71175 92654 71452 92656
rect 71175 92651 71241 92654
rect 71446 92652 71452 92654
rect 71516 92652 71522 92716
rect 93255 92714 93321 92717
rect 93710 92714 93716 92716
rect 93255 92712 93716 92714
rect 93255 92656 93260 92712
rect 93316 92656 93716 92712
rect 93255 92654 93716 92656
rect 93255 92651 93321 92654
rect 93710 92652 93716 92654
rect 93780 92652 93786 92716
rect 193438 92652 193444 92716
rect 193508 92714 193514 92716
rect 194501 92714 194567 92717
rect 212165 92714 212231 92717
rect 193508 92712 194567 92714
rect 193508 92656 194506 92712
rect 194562 92656 194567 92712
rect 193508 92654 194567 92656
rect 193508 92652 193514 92654
rect 194501 92651 194567 92654
rect 195930 92712 212231 92714
rect 195930 92656 212170 92712
rect 212226 92656 212231 92712
rect 195930 92654 212231 92656
rect 191046 92516 191052 92580
rect 191116 92578 191122 92580
rect 195930 92578 195990 92654
rect 212165 92651 212231 92654
rect 191116 92518 195990 92578
rect 218789 92578 218855 92581
rect 252553 92578 252619 92581
rect 218789 92576 252619 92578
rect 218789 92520 218794 92576
rect 218850 92520 252558 92576
rect 252614 92520 252619 92576
rect 218789 92518 252619 92520
rect 191116 92516 191122 92518
rect 218789 92515 218855 92518
rect 252553 92515 252619 92518
rect 72550 92380 72556 92444
rect 72620 92442 72626 92444
rect 73337 92442 73403 92445
rect 72620 92440 73403 92442
rect 72620 92384 73342 92440
rect 73398 92384 73403 92440
rect 72620 92382 73403 92384
rect 72620 92380 72626 92382
rect 73337 92379 73403 92382
rect 91829 92442 91895 92445
rect 95182 92442 95188 92444
rect 91829 92440 95188 92442
rect 91829 92384 91834 92440
rect 91890 92384 95188 92440
rect 91829 92382 95188 92384
rect 91829 92379 91895 92382
rect 95182 92380 95188 92382
rect 95252 92380 95258 92444
rect 206093 92442 206159 92445
rect 207054 92442 207060 92444
rect 206093 92440 207060 92442
rect 206093 92384 206098 92440
rect 206154 92384 207060 92440
rect 206093 92382 207060 92384
rect 206093 92379 206159 92382
rect 207054 92380 207060 92382
rect 207124 92380 207130 92444
rect 211654 92380 211660 92444
rect 211724 92442 211730 92444
rect 214557 92442 214623 92445
rect 211724 92440 214623 92442
rect 211724 92384 214562 92440
rect 214618 92384 214623 92440
rect 211724 92382 214623 92384
rect 211724 92380 211730 92382
rect 214557 92379 214623 92382
rect 84653 92306 84719 92309
rect 100293 92306 100359 92309
rect 84653 92304 100359 92306
rect 84653 92248 84658 92304
rect 84714 92248 100298 92304
rect 100354 92248 100359 92304
rect 84653 92246 100359 92248
rect 84653 92243 84719 92246
rect 100293 92243 100359 92246
rect 193213 92306 193279 92309
rect 231945 92306 232011 92309
rect 193213 92304 232011 92306
rect 193213 92248 193218 92304
rect 193274 92248 231950 92304
rect 232006 92248 232011 92304
rect 193213 92246 232011 92248
rect 193213 92243 193279 92246
rect 231945 92243 232011 92246
rect 86677 92170 86743 92173
rect 100109 92170 100175 92173
rect 86677 92168 100175 92170
rect 86677 92112 86682 92168
rect 86738 92112 100114 92168
rect 100170 92112 100175 92168
rect 86677 92110 100175 92112
rect 86677 92107 86743 92110
rect 100109 92107 100175 92110
rect 176009 92170 176075 92173
rect 200757 92170 200823 92173
rect 176009 92168 200823 92170
rect 176009 92112 176014 92168
rect 176070 92112 200762 92168
rect 200818 92112 200823 92168
rect 176009 92110 200823 92112
rect 176009 92107 176075 92110
rect 200757 92107 200823 92110
rect 205541 92170 205607 92173
rect 250437 92170 250503 92173
rect 205541 92168 250503 92170
rect 205541 92112 205546 92168
rect 205602 92112 250442 92168
rect 250498 92112 250503 92168
rect 205541 92110 250503 92112
rect 205541 92107 205607 92110
rect 250437 92107 250503 92110
rect 67449 92034 67515 92037
rect 187509 92034 187575 92037
rect 67449 92032 187575 92034
rect 67449 91976 67454 92032
rect 67510 91976 187514 92032
rect 187570 91976 187575 92032
rect 67449 91974 187575 91976
rect 67449 91971 67515 91974
rect 187509 91971 187575 91974
rect 188061 92034 188127 92037
rect 205633 92034 205699 92037
rect 188061 92032 205699 92034
rect 188061 91976 188066 92032
rect 188122 91976 205638 92032
rect 205694 91976 205699 92032
rect 188061 91974 205699 91976
rect 188061 91971 188127 91974
rect 205633 91971 205699 91974
rect 71773 91082 71839 91085
rect 72734 91082 72740 91084
rect 71773 91080 72740 91082
rect 71773 91024 71778 91080
rect 71834 91024 72740 91080
rect 71773 91022 72740 91024
rect 71773 91019 71839 91022
rect 72734 91020 72740 91022
rect 72804 91020 72810 91084
rect 69238 90884 69244 90948
rect 69308 90946 69314 90948
rect 76281 90946 76347 90949
rect 69308 90944 76347 90946
rect 69308 90888 76286 90944
rect 76342 90888 76347 90944
rect 69308 90886 76347 90888
rect 69308 90884 69314 90886
rect 76281 90883 76347 90886
rect 212165 90946 212231 90949
rect 239397 90946 239463 90949
rect 212165 90944 239463 90946
rect 212165 90888 212170 90944
rect 212226 90888 239402 90944
rect 239458 90888 239463 90944
rect 212165 90886 239463 90888
rect 212165 90883 212231 90886
rect 239397 90883 239463 90886
rect 46749 90810 46815 90813
rect 74257 90810 74323 90813
rect 46749 90808 74323 90810
rect 46749 90752 46754 90808
rect 46810 90752 74262 90808
rect 74318 90752 74323 90808
rect 46749 90750 74323 90752
rect 46749 90747 46815 90750
rect 74257 90747 74323 90750
rect 108297 90674 108363 90677
rect 203701 90674 203767 90677
rect 108297 90672 203767 90674
rect 108297 90616 108302 90672
rect 108358 90616 203706 90672
rect 203762 90616 203767 90672
rect 108297 90614 203767 90616
rect 108297 90611 108363 90614
rect 203701 90611 203767 90614
rect 105445 90538 105511 90541
rect 105629 90538 105695 90541
rect 204437 90538 204503 90541
rect 105445 90536 204503 90538
rect 105445 90480 105450 90536
rect 105506 90480 105634 90536
rect 105690 90480 204442 90536
rect 204498 90480 204503 90536
rect 105445 90478 204503 90480
rect 105445 90475 105511 90478
rect 105629 90475 105695 90478
rect 204437 90475 204503 90478
rect 96705 90404 96771 90405
rect 96654 90402 96660 90404
rect 96614 90342 96660 90402
rect 96724 90400 96771 90404
rect 96766 90344 96771 90400
rect 96654 90340 96660 90342
rect 96724 90340 96771 90344
rect 96705 90339 96771 90340
rect 102777 90402 102843 90405
rect 203517 90402 203583 90405
rect 102777 90400 203583 90402
rect 102777 90344 102782 90400
rect 102838 90344 203522 90400
rect 203578 90344 203583 90400
rect 102777 90342 203583 90344
rect 102777 90339 102843 90342
rect 203517 90339 203583 90342
rect 208669 90266 208735 90269
rect 209681 90266 209747 90269
rect 215293 90268 215359 90269
rect 215293 90266 215340 90268
rect 208669 90264 209747 90266
rect 208669 90208 208674 90264
rect 208730 90208 209686 90264
rect 209742 90208 209747 90264
rect 208669 90206 209747 90208
rect 215212 90264 215340 90266
rect 215404 90266 215410 90268
rect 216397 90266 216463 90269
rect 215404 90264 216463 90266
rect 215212 90208 215298 90264
rect 215404 90208 216402 90264
rect 216458 90208 216463 90264
rect 215212 90206 215340 90208
rect 208669 90203 208735 90206
rect 209681 90203 209747 90206
rect 215293 90204 215340 90206
rect 215404 90206 216463 90208
rect 215404 90204 215410 90206
rect 215293 90203 215359 90204
rect 216397 90203 216463 90206
rect 210325 89858 210391 89861
rect 209730 89856 210391 89858
rect 209730 89800 210330 89856
rect 210386 89800 210391 89856
rect 209730 89798 210391 89800
rect 82997 89722 83063 89725
rect 209730 89722 209790 89798
rect 210325 89795 210391 89798
rect 82997 89720 209790 89722
rect 82997 89664 83002 89720
rect 83058 89664 209790 89720
rect 82997 89662 209790 89664
rect 211613 89722 211679 89725
rect 236729 89722 236795 89725
rect 211613 89720 236795 89722
rect 211613 89664 211618 89720
rect 211674 89664 236734 89720
rect 236790 89664 236795 89720
rect 211613 89662 236795 89664
rect 82997 89659 83063 89662
rect 211613 89659 211679 89662
rect 236729 89659 236795 89662
rect 78029 89586 78095 89589
rect 105445 89586 105511 89589
rect 78029 89584 105511 89586
rect 78029 89528 78034 89584
rect 78090 89528 105450 89584
rect 105506 89528 105511 89584
rect 78029 89526 105511 89528
rect 78029 89523 78095 89526
rect 105445 89523 105511 89526
rect 196525 89586 196591 89589
rect 253933 89586 253999 89589
rect 196525 89584 253999 89586
rect 196525 89528 196530 89584
rect 196586 89528 253938 89584
rect 253994 89528 253999 89584
rect 196525 89526 253999 89528
rect 196525 89523 196591 89526
rect 253933 89523 253999 89526
rect 66662 89388 66668 89452
rect 66732 89450 66738 89452
rect 94630 89450 94636 89452
rect 66732 89390 94636 89450
rect 66732 89388 66738 89390
rect 94630 89388 94636 89390
rect 94700 89388 94706 89452
rect 64597 88226 64663 88229
rect 101673 88226 101739 88229
rect 64597 88224 101739 88226
rect 64597 88168 64602 88224
rect 64658 88168 101678 88224
rect 101734 88168 101739 88224
rect 64597 88166 101739 88168
rect 64597 88163 64663 88166
rect 101673 88163 101739 88166
rect 198365 88226 198431 88229
rect 287053 88226 287119 88229
rect 582833 88226 582899 88229
rect 198365 88224 582899 88226
rect 198365 88168 198370 88224
rect 198426 88168 287058 88224
rect 287114 88168 582838 88224
rect 582894 88168 582899 88224
rect 198365 88166 582899 88168
rect 198365 88163 198431 88166
rect 287053 88163 287119 88166
rect 582833 88163 582899 88166
rect 87229 88090 87295 88093
rect 121453 88090 121519 88093
rect 87229 88088 121519 88090
rect 87229 88032 87234 88088
rect 87290 88032 121458 88088
rect 121514 88032 121519 88088
rect 87229 88030 121519 88032
rect 87229 88027 87295 88030
rect 121453 88027 121519 88030
rect 80973 87954 81039 87957
rect 109677 87954 109743 87957
rect 80973 87952 109743 87954
rect 80973 87896 80978 87952
rect 81034 87896 109682 87952
rect 109738 87896 109743 87952
rect 80973 87894 109743 87896
rect 80973 87891 81039 87894
rect 109677 87891 109743 87894
rect 112529 87954 112595 87957
rect 112989 87954 113055 87957
rect 209221 87954 209287 87957
rect 112529 87952 209287 87954
rect 112529 87896 112534 87952
rect 112590 87896 112994 87952
rect 113050 87896 209226 87952
rect 209282 87896 209287 87952
rect 112529 87894 209287 87896
rect 112529 87891 112595 87894
rect 112989 87891 113055 87894
rect 209221 87891 209287 87894
rect 204437 87546 204503 87549
rect 259361 87546 259427 87549
rect 204437 87544 259427 87546
rect 204437 87488 204442 87544
rect 204498 87488 259366 87544
rect 259422 87488 259427 87544
rect 204437 87486 259427 87488
rect 204437 87483 204503 87486
rect 259361 87483 259427 87486
rect 71773 86866 71839 86869
rect 197077 86866 197143 86869
rect 71773 86864 197143 86866
rect 71773 86808 71778 86864
rect 71834 86808 197082 86864
rect 197138 86808 197143 86864
rect 71773 86806 197143 86808
rect 71773 86803 71839 86806
rect 197077 86803 197143 86806
rect 92749 86730 92815 86733
rect 116577 86730 116643 86733
rect 221917 86730 221983 86733
rect 92749 86728 221983 86730
rect 92749 86672 92754 86728
rect 92810 86672 116582 86728
rect 116638 86672 221922 86728
rect 221978 86672 221983 86728
rect 92749 86670 221983 86672
rect 92749 86667 92815 86670
rect 116577 86667 116643 86670
rect 221917 86667 221983 86670
rect 84101 86594 84167 86597
rect 101581 86594 101647 86597
rect 84101 86592 101647 86594
rect 84101 86536 84106 86592
rect 84162 86536 101586 86592
rect 101642 86536 101647 86592
rect 84101 86534 101647 86536
rect 84101 86531 84167 86534
rect 101581 86531 101647 86534
rect 192937 86186 193003 86189
rect 273253 86186 273319 86189
rect 192937 86184 273319 86186
rect 192937 86128 192942 86184
rect 192998 86128 273258 86184
rect 273314 86128 273319 86184
rect 192937 86126 273319 86128
rect 192937 86123 193003 86126
rect 273253 86123 273319 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 98637 85506 98703 85509
rect 190361 85506 190427 85509
rect 220077 85506 220143 85509
rect 98637 85504 220143 85506
rect 98637 85448 98642 85504
rect 98698 85448 190366 85504
rect 190422 85448 220082 85504
rect 220138 85448 220143 85504
rect 98637 85446 220143 85448
rect 98637 85443 98703 85446
rect 190361 85443 190427 85446
rect 220077 85443 220143 85446
rect 78397 85370 78463 85373
rect 107653 85370 107719 85373
rect 108113 85370 108179 85373
rect 78397 85368 108179 85370
rect 78397 85312 78402 85368
rect 78458 85312 107658 85368
rect 107714 85312 108118 85368
rect 108174 85312 108179 85368
rect 78397 85310 108179 85312
rect 78397 85307 78463 85310
rect 107653 85307 107719 85310
rect 108113 85307 108179 85310
rect 91277 85234 91343 85237
rect 98637 85234 98703 85237
rect 91277 85232 98703 85234
rect 91277 85176 91282 85232
rect 91338 85176 98642 85232
rect 98698 85176 98703 85232
rect 91277 85174 98703 85176
rect 91277 85171 91343 85174
rect 98637 85171 98703 85174
rect 191373 84826 191439 84829
rect 327717 84826 327783 84829
rect 191373 84824 327783 84826
rect -960 84690 480 84780
rect 191373 84768 191378 84824
rect 191434 84768 327722 84824
rect 327778 84768 327783 84824
rect 191373 84766 327783 84768
rect 191373 84763 191439 84766
rect 327717 84763 327783 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 65885 84146 65951 84149
rect 186313 84146 186379 84149
rect 65885 84144 186379 84146
rect 65885 84088 65890 84144
rect 65946 84088 186318 84144
rect 186374 84088 186379 84144
rect 65885 84086 186379 84088
rect 65885 84083 65951 84086
rect 186313 84083 186379 84086
rect 188337 84146 188403 84149
rect 227805 84146 227871 84149
rect 188337 84144 227871 84146
rect 188337 84088 188342 84144
rect 188398 84088 227810 84144
rect 227866 84088 227871 84144
rect 188337 84086 227871 84088
rect 188337 84083 188403 84086
rect 227805 84083 227871 84086
rect 85665 84010 85731 84013
rect 104157 84010 104223 84013
rect 85665 84008 104223 84010
rect 85665 83952 85670 84008
rect 85726 83952 104162 84008
rect 104218 83952 104223 84008
rect 85665 83950 104223 83952
rect 85665 83947 85731 83950
rect 104157 83947 104223 83950
rect 93117 83466 93183 83469
rect 96613 83466 96679 83469
rect 93117 83464 96679 83466
rect 93117 83408 93122 83464
rect 93178 83408 96618 83464
rect 96674 83408 96679 83464
rect 93117 83406 96679 83408
rect 93117 83403 93183 83406
rect 96613 83403 96679 83406
rect 192702 83404 192708 83468
rect 192772 83466 192778 83468
rect 259545 83466 259611 83469
rect 192772 83464 259611 83466
rect 192772 83408 259550 83464
rect 259606 83408 259611 83464
rect 192772 83406 259611 83408
rect 192772 83404 192778 83406
rect 259545 83403 259611 83406
rect 186313 82922 186379 82925
rect 186957 82922 187023 82925
rect 186313 82920 187023 82922
rect 186313 82864 186318 82920
rect 186374 82864 186962 82920
rect 187018 82864 187023 82920
rect 186313 82862 187023 82864
rect 186313 82859 186379 82862
rect 186957 82859 187023 82862
rect 89989 82786 90055 82789
rect 124857 82786 124923 82789
rect 89989 82784 124923 82786
rect 89989 82728 89994 82784
rect 90050 82728 124862 82784
rect 124918 82728 124923 82784
rect 89989 82726 124923 82728
rect 89989 82723 90055 82726
rect 124857 82723 124923 82726
rect 69606 82588 69612 82652
rect 69676 82650 69682 82652
rect 94446 82650 94452 82652
rect 69676 82590 94452 82650
rect 69676 82588 69682 82590
rect 94446 82588 94452 82590
rect 94516 82588 94522 82652
rect 70301 82106 70367 82109
rect 189942 82106 189948 82108
rect 70301 82104 189948 82106
rect 70301 82048 70306 82104
rect 70362 82048 189948 82104
rect 70301 82046 189948 82048
rect 70301 82043 70367 82046
rect 189942 82044 189948 82046
rect 190012 82044 190018 82108
rect 193806 82044 193812 82108
rect 193876 82106 193882 82108
rect 269113 82106 269179 82109
rect 193876 82104 269179 82106
rect 193876 82048 269118 82104
rect 269174 82048 269179 82104
rect 193876 82046 269179 82048
rect 193876 82044 193882 82046
rect 269113 82043 269179 82046
rect 106181 81426 106247 81429
rect 226374 81426 226380 81428
rect 106181 81424 226380 81426
rect 106181 81368 106186 81424
rect 106242 81368 226380 81424
rect 106181 81366 226380 81368
rect 106181 81363 106247 81366
rect 226374 81364 226380 81366
rect 226444 81364 226450 81428
rect 68277 81290 68343 81293
rect 156689 81290 156755 81293
rect 68277 81288 156755 81290
rect 68277 81232 68282 81288
rect 68338 81232 156694 81288
rect 156750 81232 156755 81288
rect 68277 81230 156755 81232
rect 68277 81227 68343 81230
rect 156689 81227 156755 81230
rect 203701 81290 203767 81293
rect 284385 81290 284451 81293
rect 203701 81288 287070 81290
rect 203701 81232 203706 81288
rect 203762 81232 284390 81288
rect 284446 81232 287070 81288
rect 203701 81230 287070 81232
rect 203701 81227 203767 81230
rect 284385 81227 284451 81230
rect 77293 81154 77359 81157
rect 108297 81154 108363 81157
rect 77293 81152 108363 81154
rect 77293 81096 77298 81152
rect 77354 81096 108302 81152
rect 108358 81096 108363 81152
rect 77293 81094 108363 81096
rect 77293 81091 77359 81094
rect 108297 81091 108363 81094
rect 287010 80746 287070 81230
rect 582833 80746 582899 80749
rect 287010 80744 582899 80746
rect 287010 80688 582838 80744
rect 582894 80688 582899 80744
rect 287010 80686 582899 80688
rect 582833 80683 582899 80686
rect 89897 80066 89963 80069
rect 220169 80066 220235 80069
rect 89897 80064 220235 80066
rect 89897 80008 89902 80064
rect 89958 80008 220174 80064
rect 220230 80008 220235 80064
rect 89897 80006 220235 80008
rect 89897 80003 89963 80006
rect 220169 80003 220235 80006
rect 61377 79930 61443 79933
rect 97942 79930 97948 79932
rect 61377 79928 97948 79930
rect 61377 79872 61382 79928
rect 61438 79872 97948 79928
rect 61377 79870 97948 79872
rect 61377 79867 61443 79870
rect 97942 79868 97948 79870
rect 98012 79868 98018 79932
rect 181253 79930 181319 79933
rect 182081 79930 182147 79933
rect 210049 79930 210115 79933
rect 181253 79928 210115 79930
rect 181253 79872 181258 79928
rect 181314 79872 182086 79928
rect 182142 79872 210054 79928
rect 210110 79872 210115 79928
rect 181253 79870 210115 79872
rect 181253 79867 181319 79870
rect 182081 79867 182147 79870
rect 209730 79386 209790 79870
rect 210049 79867 210115 79870
rect 582925 79386 582991 79389
rect 209730 79384 582991 79386
rect 209730 79328 582930 79384
rect 582986 79328 582991 79384
rect 209730 79326 582991 79328
rect 582925 79323 582991 79326
rect 188981 78570 189047 78573
rect 284293 78570 284359 78573
rect 188981 78568 284359 78570
rect 188981 78512 188986 78568
rect 189042 78512 284298 78568
rect 284354 78512 284359 78568
rect 188981 78510 284359 78512
rect 188981 78507 189047 78510
rect 284293 78507 284359 78510
rect 86861 77890 86927 77893
rect 188286 77890 188292 77892
rect 86861 77888 188292 77890
rect 86861 77832 86866 77888
rect 86922 77832 188292 77888
rect 86861 77830 188292 77832
rect 86861 77827 86927 77830
rect 188286 77828 188292 77830
rect 188356 77828 188362 77892
rect 196566 77828 196572 77892
rect 196636 77890 196642 77892
rect 262213 77890 262279 77893
rect 196636 77888 262279 77890
rect 196636 77832 262218 77888
rect 262274 77832 262279 77888
rect 196636 77830 262279 77832
rect 196636 77828 196642 77830
rect 262213 77827 262279 77830
rect 101489 77210 101555 77213
rect 207657 77210 207723 77213
rect 101489 77208 207723 77210
rect 101489 77152 101494 77208
rect 101550 77152 207662 77208
rect 207718 77152 207723 77208
rect 101489 77150 207723 77152
rect 101489 77147 101555 77150
rect 207657 77147 207723 77150
rect 65977 77074 66043 77077
rect 123477 77074 123543 77077
rect 65977 77072 123543 77074
rect 65977 77016 65982 77072
rect 66038 77016 123482 77072
rect 123538 77016 123543 77072
rect 65977 77014 123543 77016
rect 65977 77011 66043 77014
rect 123477 77011 123543 77014
rect 178769 77074 178835 77077
rect 233233 77074 233299 77077
rect 178769 77072 233299 77074
rect 178769 77016 178774 77072
rect 178830 77016 233238 77072
rect 233294 77016 233299 77072
rect 178769 77014 233299 77016
rect 178769 77011 178835 77014
rect 233233 77011 233299 77014
rect 173249 75850 173315 75853
rect 229093 75850 229159 75853
rect 173249 75848 229159 75850
rect 173249 75792 173254 75848
rect 173310 75792 229098 75848
rect 229154 75792 229159 75848
rect 173249 75790 229159 75792
rect 173249 75787 173315 75790
rect 229093 75787 229159 75790
rect 177389 75714 177455 75717
rect 230565 75714 230631 75717
rect 177389 75712 230631 75714
rect 177389 75656 177394 75712
rect 177450 75656 230570 75712
rect 230626 75656 230631 75712
rect 177389 75654 230631 75656
rect 177389 75651 177455 75654
rect 230565 75651 230631 75654
rect 95141 75170 95207 75173
rect 104249 75170 104315 75173
rect 95141 75168 104315 75170
rect 95141 75112 95146 75168
rect 95202 75112 104254 75168
rect 104310 75112 104315 75168
rect 95141 75110 104315 75112
rect 95141 75107 95207 75110
rect 104249 75107 104315 75110
rect 98729 74490 98795 74493
rect 224902 74490 224908 74492
rect 98729 74488 224908 74490
rect 98729 74432 98734 74488
rect 98790 74432 224908 74488
rect 98729 74430 224908 74432
rect 98729 74427 98795 74430
rect 224902 74428 224908 74430
rect 224972 74428 224978 74492
rect 582373 72994 582439 72997
rect 583520 72994 584960 73084
rect 582373 72992 584960 72994
rect 582373 72936 582378 72992
rect 582434 72936 584960 72992
rect 582373 72934 584960 72936
rect 582373 72931 582439 72934
rect 583520 72844 584960 72934
rect 62021 72450 62087 72453
rect 180149 72450 180215 72453
rect 62021 72448 180215 72450
rect 62021 72392 62026 72448
rect 62082 72392 180154 72448
rect 180210 72392 180215 72448
rect 62021 72390 180215 72392
rect 62021 72387 62087 72390
rect 180149 72387 180215 72390
rect 194501 72450 194567 72453
rect 298093 72450 298159 72453
rect 194501 72448 298159 72450
rect 194501 72392 194506 72448
rect 194562 72392 298098 72448
rect 298154 72392 298159 72448
rect 194501 72390 298159 72392
rect 194501 72387 194567 72390
rect 298093 72387 298159 72390
rect -960 71634 480 71724
rect 3141 71634 3207 71637
rect -960 71632 3207 71634
rect -960 71576 3146 71632
rect 3202 71576 3207 71632
rect -960 71574 3207 71576
rect -960 71484 480 71574
rect 3141 71571 3207 71574
rect 582741 59666 582807 59669
rect 583520 59666 584960 59756
rect 582741 59664 584960 59666
rect 582741 59608 582746 59664
rect 582802 59608 584960 59664
rect 582741 59606 584960 59608
rect 582741 59603 582807 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3325 45522 3391 45525
rect -960 45520 3391 45522
rect -960 45464 3330 45520
rect 3386 45464 3391 45520
rect -960 45462 3391 45464
rect -960 45372 480 45462
rect 3325 45459 3391 45462
rect 37089 44842 37155 44845
rect 170254 44842 170260 44844
rect 37089 44840 170260 44842
rect 37089 44784 37094 44840
rect 37150 44784 170260 44840
rect 37089 44782 170260 44784
rect 37089 44779 37155 44782
rect 170254 44780 170260 44782
rect 170324 44780 170330 44844
rect 582925 33146 582991 33149
rect 583520 33146 584960 33236
rect 582925 33144 584960 33146
rect 582925 33088 582930 33144
rect 582986 33088 584960 33144
rect 582925 33086 584960 33088
rect 582925 33083 582991 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 206870 32404 206876 32468
rect 206940 32466 206946 32468
rect 318793 32466 318859 32469
rect 206940 32464 318859 32466
rect 206940 32408 318798 32464
rect 318854 32408 318859 32464
rect 206940 32406 318859 32408
rect 206940 32404 206946 32406
rect 318793 32403 318859 32406
rect 582649 19818 582715 19821
rect 583520 19818 584960 19908
rect 582649 19816 584960 19818
rect 582649 19760 582654 19816
rect 582710 19760 584960 19816
rect 582649 19758 584960 19760
rect 582649 19755 582715 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 582833 6626 582899 6629
rect 583520 6626 584960 6716
rect 582833 6624 584960 6626
rect -960 6490 480 6580
rect 582833 6568 582838 6624
rect 582894 6568 584960 6624
rect 582833 6566 584960 6568
rect 582833 6563 582899 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 300117 3634 300183 3637
rect 304349 3634 304415 3637
rect 300117 3632 304415 3634
rect 300117 3576 300122 3632
rect 300178 3576 304354 3632
rect 304410 3576 304415 3632
rect 300117 3574 304415 3576
rect 300117 3571 300183 3574
rect 304349 3571 304415 3574
rect 97441 3498 97507 3501
rect 130377 3498 130443 3501
rect 97441 3496 130443 3498
rect 97441 3440 97446 3496
rect 97502 3440 130382 3496
rect 130438 3440 130443 3496
rect 97441 3438 130443 3440
rect 97441 3435 97507 3438
rect 130377 3435 130443 3438
rect 302877 3498 302943 3501
rect 305545 3498 305611 3501
rect 302877 3496 305611 3498
rect 302877 3440 302882 3496
rect 302938 3440 305550 3496
rect 305606 3440 305611 3496
rect 302877 3438 305611 3440
rect 302877 3435 302943 3438
rect 305545 3435 305611 3438
rect 104525 3362 104591 3365
rect 148317 3362 148383 3365
rect 104525 3360 148383 3362
rect 104525 3304 104530 3360
rect 104586 3304 148322 3360
rect 148378 3304 148383 3360
rect 104525 3302 148383 3304
rect 104525 3299 104591 3302
rect 148317 3299 148383 3302
rect 286317 3362 286383 3365
rect 293677 3362 293743 3365
rect 286317 3360 293743 3362
rect 286317 3304 286322 3360
rect 286378 3304 293682 3360
rect 293738 3304 293743 3360
rect 286317 3302 293743 3304
rect 286317 3299 286383 3302
rect 293677 3299 293743 3302
<< via3 >>
rect 75868 596260 75932 596324
rect 83412 582388 83476 582452
rect 75684 581028 75748 581092
rect 71636 580756 71700 580820
rect 72924 580756 72988 580820
rect 79916 580816 79980 580820
rect 79916 580760 79930 580816
rect 79930 580760 79980 580816
rect 79916 580756 79980 580760
rect 88380 580756 88444 580820
rect 91692 580756 91756 580820
rect 104940 571372 105004 571436
rect 115060 569196 115124 569260
rect 69428 550836 69492 550900
rect 115980 550700 116044 550764
rect 96660 547028 96724 547092
rect 69428 543492 69492 543556
rect 75868 539548 75932 539612
rect 73292 537508 73356 537572
rect 91692 537508 91756 537572
rect 69796 537372 69860 537436
rect 106412 534788 106476 534852
rect 96660 534652 96724 534716
rect 79732 523636 79796 523700
rect 72740 520916 72804 520980
rect 96660 479436 96724 479500
rect 75684 476716 75748 476780
rect 107700 472500 107764 472564
rect 67772 468420 67836 468484
rect 69612 466576 69676 466580
rect 69612 466520 69662 466576
rect 69662 466520 69676 466576
rect 69612 466516 69676 466520
rect 72924 464340 72988 464404
rect 113220 464340 113284 464404
rect 262260 462300 262324 462364
rect 83412 460124 83476 460188
rect 97212 460124 97276 460188
rect 83596 459580 83660 459644
rect 99972 458764 100036 458828
rect 195836 458280 195900 458284
rect 195836 458224 195850 458280
rect 195850 458224 195900 458280
rect 195836 458220 195900 458224
rect 247724 456996 247788 457060
rect 252692 455636 252756 455700
rect 284340 455500 284404 455564
rect 276244 454140 276308 454204
rect 244780 454004 244844 454068
rect 197124 453052 197188 453116
rect 242020 452644 242084 452708
rect 254532 452644 254596 452708
rect 88380 449924 88444 449988
rect 241652 449924 241716 449988
rect 248460 449984 248524 449988
rect 248460 449928 248510 449984
rect 248510 449928 248524 449984
rect 248460 449924 248524 449928
rect 193444 449712 193508 449716
rect 193444 449656 193494 449712
rect 193494 449656 193508 449712
rect 193444 449652 193508 449656
rect 245700 449712 245764 449716
rect 245700 449656 245750 449712
rect 245750 449656 245764 449712
rect 245700 449652 245764 449656
rect 101260 448564 101324 448628
rect 66116 446388 66180 446452
rect 193444 445572 193508 445636
rect 69612 442988 69676 443052
rect 83596 439452 83660 439516
rect 107884 438092 107948 438156
rect 114324 436868 114388 436932
rect 262260 436928 262324 436932
rect 263364 436928 263428 436932
rect 262260 436872 262310 436928
rect 262310 436872 262324 436928
rect 263364 436872 263414 436928
rect 263414 436872 263428 436928
rect 262260 436868 262324 436872
rect 263364 436868 263428 436872
rect 94636 436188 94700 436252
rect 71820 436112 71884 436116
rect 71820 436056 71870 436112
rect 71870 436056 71884 436112
rect 71820 436052 71884 436056
rect 81020 436052 81084 436116
rect 83596 436052 83660 436116
rect 94452 436052 94516 436116
rect 73660 435372 73724 435436
rect 71636 434828 71700 434892
rect 67404 434556 67468 434620
rect 102732 434556 102796 434620
rect 69060 434284 69124 434348
rect 76420 434344 76484 434348
rect 76420 434288 76434 434344
rect 76434 434288 76484 434344
rect 76420 434284 76484 434288
rect 81940 434344 82004 434348
rect 81940 434288 81954 434344
rect 81954 434288 82004 434344
rect 81940 434284 82004 434288
rect 83044 434344 83108 434348
rect 83044 434288 83094 434344
rect 83094 434288 83108 434344
rect 83044 434284 83108 434288
rect 84700 434344 84764 434348
rect 84700 434288 84714 434344
rect 84714 434288 84764 434344
rect 84700 434284 84764 434288
rect 85804 434344 85868 434348
rect 85804 434288 85854 434344
rect 85854 434288 85868 434344
rect 85804 434284 85868 434288
rect 96292 434344 96356 434348
rect 96292 434288 96306 434344
rect 96306 434288 96356 434344
rect 96292 434284 96356 434288
rect 100524 434284 100588 434348
rect 92980 434148 93044 434212
rect 83228 434012 83292 434076
rect 67956 433876 68020 433940
rect 70900 433740 70964 433804
rect 74580 433604 74644 433668
rect 77340 433604 77404 433668
rect 87092 433604 87156 433668
rect 87460 433604 87524 433668
rect 89668 433664 89732 433668
rect 89668 433608 89682 433664
rect 89682 433608 89732 433664
rect 89668 433604 89732 433608
rect 90036 433664 90100 433668
rect 90036 433608 90086 433664
rect 90086 433608 90100 433664
rect 90036 433604 90100 433608
rect 91324 433664 91388 433668
rect 91324 433608 91338 433664
rect 91338 433608 91388 433664
rect 91324 433604 91388 433608
rect 91508 433664 91572 433668
rect 91508 433608 91558 433664
rect 91558 433608 91572 433664
rect 91508 433604 91572 433608
rect 92796 433604 92860 433668
rect 97948 433604 98012 433668
rect 98500 433604 98564 433668
rect 100708 433664 100772 433668
rect 100708 433608 100722 433664
rect 100722 433608 100772 433664
rect 100708 433604 100772 433608
rect 105492 433604 105556 433668
rect 108988 433664 109052 433668
rect 108988 433608 109038 433664
rect 109038 433608 109052 433664
rect 108988 433604 109052 433608
rect 281580 431156 281644 431220
rect 69428 429796 69492 429860
rect 112116 426532 112180 426596
rect 193812 423676 193876 423740
rect 67956 422180 68020 422244
rect 66300 417420 66364 417484
rect 177252 415924 177316 415988
rect 66300 412992 66364 412996
rect 66300 412936 66314 412992
rect 66314 412936 66364 412992
rect 66300 412932 66364 412936
rect 191604 412660 191668 412724
rect 66116 411844 66180 411908
rect 115060 409940 115124 410004
rect 67404 409668 67468 409732
rect 114324 405452 114388 405516
rect 66668 401644 66732 401708
rect 188844 400420 188908 400484
rect 256004 397972 256068 398036
rect 67772 397428 67836 397492
rect 113220 397156 113284 397220
rect 270540 396612 270604 396676
rect 193996 396476 194060 396540
rect 69428 393892 69492 393956
rect 112852 393484 112916 393548
rect 73476 390900 73540 390964
rect 107884 390688 107948 390692
rect 107884 390632 107934 390688
rect 107934 390632 107948 390688
rect 96660 390492 96724 390556
rect 101260 390492 101324 390556
rect 107884 390628 107948 390632
rect 112852 390628 112916 390692
rect 193996 390492 194060 390556
rect 99972 390356 100036 390420
rect 104940 390356 105004 390420
rect 106412 390356 106476 390420
rect 107700 390416 107764 390420
rect 107700 390360 107750 390416
rect 107750 390360 107764 390416
rect 107700 390356 107764 390360
rect 248460 389812 248524 389876
rect 72740 388996 72804 389060
rect 79732 388996 79796 389060
rect 80100 389056 80164 389060
rect 80100 389000 80114 389056
rect 80114 389000 80164 389056
rect 80100 388996 80164 389000
rect 97212 388860 97276 388924
rect 91324 387772 91388 387836
rect 269436 387500 269500 387564
rect 87460 386956 87524 387020
rect 81940 386140 82004 386204
rect 115980 386140 116044 386204
rect 100708 385596 100772 385660
rect 258396 385596 258460 385660
rect 90036 384236 90100 384300
rect 101260 384236 101324 384300
rect 94636 383692 94700 383756
rect 81020 382876 81084 382940
rect 195836 381516 195900 381580
rect 197124 380836 197188 380900
rect 274588 380156 274652 380220
rect 191604 379340 191668 379404
rect 266308 379204 266372 379268
rect 191604 378932 191668 378996
rect 96660 378660 96724 378724
rect 265756 377980 265820 378044
rect 255820 377300 255884 377364
rect 69612 375260 69676 375324
rect 188844 373900 188908 373964
rect 77340 373220 77404 373284
rect 252508 373220 252572 373284
rect 188844 372812 188908 372876
rect 193812 371860 193876 371924
rect 242020 371316 242084 371380
rect 66668 369684 66732 369748
rect 256004 369684 256068 369748
rect 273300 369004 273364 369068
rect 241652 366420 241716 366484
rect 252692 366284 252756 366348
rect 267780 363564 267844 363628
rect 245700 361660 245764 361724
rect 277164 359348 277228 359412
rect 258396 358668 258460 358732
rect 191604 346972 191668 347036
rect 250300 345612 250364 345676
rect 241652 344252 241716 344316
rect 269252 338676 269316 338740
rect 102732 329020 102796 329084
rect 254532 328340 254596 328404
rect 259500 323640 259564 323644
rect 259500 323584 259514 323640
rect 259514 323584 259564 323640
rect 259500 323580 259564 323584
rect 85804 322764 85868 322828
rect 84700 320044 84764 320108
rect 94452 319364 94516 319428
rect 105492 319364 105556 319428
rect 87092 318004 87156 318068
rect 97948 318004 98012 318068
rect 188476 317732 188540 317796
rect 267964 317596 268028 317660
rect 83044 317324 83108 317388
rect 84516 317324 84580 317388
rect 74580 316100 74644 316164
rect 258396 315284 258460 315348
rect 263548 311204 263612 311268
rect 280292 311068 280356 311132
rect 89668 309844 89732 309908
rect 96292 309708 96356 309772
rect 108988 309708 109052 309772
rect 260972 309708 261036 309772
rect 186820 308076 186884 308140
rect 166212 306580 166276 306644
rect 192524 306444 192588 306508
rect 100524 305220 100588 305284
rect 257292 305084 257356 305148
rect 258396 305084 258460 305148
rect 244780 304540 244844 304604
rect 100524 304132 100588 304196
rect 188292 303860 188356 303924
rect 189948 303724 190012 303788
rect 71820 303588 71884 303652
rect 197124 303588 197188 303652
rect 247724 303588 247788 303652
rect 259684 303588 259748 303652
rect 258396 302772 258460 302836
rect 192340 301412 192404 301476
rect 254532 301608 254596 301612
rect 254532 301552 254582 301608
rect 254582 301552 254596 301608
rect 254532 301548 254596 301552
rect 193444 301140 193508 301204
rect 193260 301064 193324 301068
rect 193260 301008 193310 301064
rect 193310 301008 193324 301064
rect 193260 301004 193324 301008
rect 241652 301004 241716 301068
rect 191604 300868 191668 300932
rect 194548 300868 194612 300932
rect 197308 300868 197372 300932
rect 250300 300188 250364 300252
rect 197308 300052 197372 300116
rect 188476 298692 188540 298756
rect 259684 298072 259748 298076
rect 259684 298016 259698 298072
rect 259698 298016 259748 298072
rect 259684 298012 259748 298016
rect 91508 297468 91572 297532
rect 191604 297468 191668 297532
rect 193812 297468 193876 297532
rect 193260 297332 193324 297396
rect 192340 294476 192404 294540
rect 191788 294340 191852 294404
rect 92796 293252 92860 293316
rect 98500 293116 98564 293180
rect 193444 293116 193508 293180
rect 83228 292572 83292 292636
rect 193444 292708 193508 292772
rect 263548 292496 263612 292500
rect 263548 292440 263562 292496
rect 263562 292440 263612 292496
rect 263548 292436 263612 292440
rect 191788 292300 191852 292364
rect 92980 291756 93044 291820
rect 86540 291076 86604 291140
rect 184060 290940 184124 291004
rect 191052 289988 191116 290052
rect 91508 289852 91572 289916
rect 88012 289716 88076 289780
rect 258396 289776 258460 289832
rect 258396 289768 258410 289776
rect 258410 289768 258460 289776
rect 259500 289580 259564 289644
rect 177252 289036 177316 289100
rect 192708 288900 192772 288964
rect 90956 288492 91020 288556
rect 177804 288492 177868 288556
rect 70900 288356 70964 288420
rect 192524 288356 192588 288420
rect 192340 287812 192404 287876
rect 66668 287676 66732 287740
rect 72924 286044 72988 286108
rect 95188 285908 95252 285972
rect 70900 285832 70964 285836
rect 70900 285776 70914 285832
rect 70914 285776 70964 285832
rect 70900 285772 70964 285776
rect 70900 285636 70964 285700
rect 258396 285016 258460 285020
rect 76420 284820 76484 284884
rect 258396 284960 258410 285016
rect 258410 284960 258460 285016
rect 258396 284956 258460 284960
rect 86724 283792 86788 283796
rect 86724 283736 86738 283792
rect 86738 283736 86788 283792
rect 86724 283732 86788 283736
rect 71636 283596 71700 283660
rect 68692 283460 68756 283524
rect 89484 283520 89548 283524
rect 89484 283464 89534 283520
rect 89534 283464 89548 283520
rect 89484 283460 89548 283464
rect 90036 283520 90100 283524
rect 90036 283464 90086 283520
rect 90086 283464 90100 283520
rect 90036 283460 90100 283464
rect 93900 283460 93964 283524
rect 194180 283324 194244 283388
rect 69244 283188 69308 283252
rect 83412 283248 83476 283252
rect 83412 283192 83462 283248
rect 83462 283192 83476 283248
rect 83412 283188 83476 283192
rect 84700 283188 84764 283252
rect 71636 283052 71700 283116
rect 73292 283052 73356 283116
rect 72372 282976 72436 282980
rect 72372 282920 72422 282976
rect 72422 282920 72436 282976
rect 72372 282916 72436 282920
rect 73476 282976 73540 282980
rect 73476 282920 73526 282976
rect 73526 282920 73540 282976
rect 73476 282916 73540 282920
rect 263548 282976 263612 282980
rect 263548 282920 263562 282976
rect 263562 282920 263612 282976
rect 263548 282916 263612 282920
rect 69060 282780 69124 282844
rect 67956 280468 68020 280532
rect 166212 280060 166276 280124
rect 111748 278156 111812 278220
rect 257292 278020 257356 278084
rect 98500 277476 98564 277540
rect 101260 276932 101324 276996
rect 69244 275980 69308 276044
rect 101260 275300 101324 275364
rect 258580 275164 258644 275228
rect 99972 270404 100036 270468
rect 98132 267820 98196 267884
rect 148180 265508 148244 265572
rect 260972 264420 261036 264484
rect 260972 264284 261036 264348
rect 262260 264148 262324 264212
rect 284340 264148 284404 264212
rect 269252 263332 269316 263396
rect 270540 262788 270604 262852
rect 265756 262652 265820 262716
rect 263548 262244 263612 262308
rect 280292 262168 280356 262172
rect 280292 262112 280306 262168
rect 280306 262112 280356 262168
rect 280292 262108 280356 262112
rect 263180 261564 263244 261628
rect 269068 260748 269132 260812
rect 273300 260748 273364 260812
rect 258396 260476 258460 260540
rect 263364 260068 263428 260132
rect 265756 260068 265820 260132
rect 262260 259932 262324 259996
rect 285628 259584 285692 259588
rect 285628 259528 285678 259584
rect 285678 259528 285692 259584
rect 285628 259524 285692 259528
rect 269068 259388 269132 259452
rect 273300 259388 273364 259452
rect 274588 259388 274652 259452
rect 191236 258708 191300 258772
rect 267780 258164 267844 258228
rect 255820 257892 255884 257956
rect 259684 257892 259748 257956
rect 254532 257484 254596 257548
rect 267780 257408 267844 257412
rect 267780 257352 267794 257408
rect 267794 257352 267844 257408
rect 267780 257348 267844 257352
rect 66668 256668 66732 256732
rect 66116 255308 66180 255372
rect 177252 255308 177316 255372
rect 276428 255368 276492 255372
rect 276428 255312 276442 255368
rect 276442 255312 276492 255368
rect 276428 255308 276492 255312
rect 269436 255172 269500 255236
rect 270540 255172 270604 255236
rect 184980 253948 185044 254012
rect 252876 253948 252940 254012
rect 100708 252452 100772 252516
rect 266492 252588 266556 252652
rect 69060 250548 69124 250612
rect 101260 250412 101324 250476
rect 170260 248372 170324 248436
rect 258396 247692 258460 247756
rect 184060 247556 184124 247620
rect 66668 247012 66732 247076
rect 266308 246196 266372 246260
rect 276244 245516 276308 245580
rect 184060 244564 184124 244628
rect 184244 244428 184308 244492
rect 69428 244292 69492 244356
rect 267964 244156 268028 244220
rect 253612 243612 253676 243676
rect 102732 243476 102796 243540
rect 193444 242796 193508 242860
rect 281580 242252 281644 242316
rect 70900 241768 70964 241772
rect 70900 241712 70950 241768
rect 70950 241712 70964 241768
rect 70900 241708 70964 241712
rect 84516 241708 84580 241772
rect 86540 241768 86604 241772
rect 86540 241712 86590 241768
rect 86590 241712 86604 241768
rect 86540 241708 86604 241712
rect 90956 241708 91020 241772
rect 91508 241768 91572 241772
rect 91508 241712 91558 241768
rect 91558 241712 91572 241768
rect 91508 241708 91572 241712
rect 88012 241572 88076 241636
rect 195836 242040 195900 242044
rect 195836 241984 195850 242040
rect 195850 241984 195900 242040
rect 195836 241980 195900 241984
rect 248460 242040 248524 242044
rect 248460 241984 248510 242040
rect 248510 241984 248524 242040
rect 248460 241980 248524 241984
rect 67956 241436 68020 241500
rect 277164 241436 277228 241500
rect 258396 240212 258460 240276
rect 277164 240212 277228 240276
rect 68876 240076 68940 240140
rect 71452 240136 71516 240140
rect 71452 240080 71466 240136
rect 71466 240080 71516 240136
rect 71452 240076 71516 240080
rect 72372 240076 72436 240140
rect 72924 240136 72988 240140
rect 72924 240080 72974 240136
rect 72974 240080 72988 240136
rect 72924 240076 72988 240080
rect 73292 240076 73356 240140
rect 90956 240136 91020 240140
rect 90956 240080 90970 240136
rect 90970 240080 91020 240136
rect 90956 240076 91020 240080
rect 97764 240076 97828 240140
rect 72740 239940 72804 240004
rect 72556 239804 72620 239868
rect 88012 239804 88076 239868
rect 192340 239804 192404 239868
rect 96660 239396 96724 239460
rect 259684 239396 259748 239460
rect 84516 238716 84580 238780
rect 96660 238716 96724 238780
rect 200620 238036 200684 238100
rect 93716 237356 93780 237420
rect 208348 236540 208412 236604
rect 69612 235860 69676 235924
rect 258396 235860 258460 235924
rect 193812 235180 193876 235244
rect 248460 235180 248524 235244
rect 97580 233956 97644 234020
rect 99972 233956 100036 234020
rect 192708 233820 192772 233884
rect 207060 233820 207124 233884
rect 207060 233004 207124 233068
rect 191236 231780 191300 231844
rect 187004 231100 187068 231164
rect 276428 231100 276492 231164
rect 263548 228924 263612 228988
rect 69060 227564 69124 227628
rect 267780 227564 267844 227628
rect 93900 227020 93964 227084
rect 69060 226884 69124 226948
rect 90036 226340 90100 226404
rect 265756 225524 265820 225588
rect 66668 224844 66732 224908
rect 102732 224708 102796 224772
rect 177804 224708 177868 224772
rect 194548 221444 194612 221508
rect 95188 220900 95252 220964
rect 270540 220084 270604 220148
rect 269068 219268 269132 219332
rect 184244 218588 184308 218652
rect 269068 218044 269132 218108
rect 197124 217364 197188 217428
rect 202092 214644 202156 214708
rect 260972 214644 261036 214708
rect 273300 214508 273364 214572
rect 72740 213828 72804 213892
rect 71452 211788 71516 211852
rect 97764 210292 97828 210356
rect 210372 208932 210436 208996
rect 97212 205668 97276 205732
rect 266492 204852 266556 204916
rect 184980 203492 185044 203556
rect 195836 202268 195900 202332
rect 253060 202132 253124 202196
rect 186820 199276 186884 199340
rect 187004 196556 187068 196620
rect 86540 190980 86604 191044
rect 215340 189076 215404 189140
rect 184060 186900 184124 186964
rect 262260 186900 262324 186964
rect 148180 182820 148244 182884
rect 69612 180780 69676 180844
rect 211660 175884 211724 175948
rect 89484 175340 89548 175404
rect 90956 169764 91020 169828
rect 86724 169084 86788 169148
rect 83412 169008 83476 169012
rect 83412 168952 83462 169008
rect 83462 168952 83476 169008
rect 83412 168948 83476 168952
rect 86724 168404 86788 168468
rect 96660 167724 96724 167788
rect 222332 167724 222396 167788
rect 227668 167588 227732 167652
rect 68692 165548 68756 165612
rect 93532 161468 93596 161532
rect 68140 160788 68204 160852
rect 191052 160652 191116 160716
rect 194364 157932 194428 157996
rect 71636 153036 71700 153100
rect 71636 152084 71700 152148
rect 224908 149636 224972 149700
rect 285628 148412 285692 148476
rect 259500 146916 259564 146980
rect 97948 146372 98012 146436
rect 226380 146236 226444 146300
rect 226564 145012 226628 145076
rect 196572 143380 196636 143444
rect 73476 142292 73540 142356
rect 196572 142292 196636 142356
rect 224356 142156 224420 142220
rect 193076 141068 193140 141132
rect 69796 140932 69860 140996
rect 73476 140796 73540 140860
rect 196572 140388 196636 140452
rect 193444 140116 193508 140180
rect 206876 140388 206940 140452
rect 225276 140388 225340 140452
rect 222332 140116 222396 140180
rect 226564 139844 226628 139908
rect 193076 139028 193140 139092
rect 192708 138212 192772 138276
rect 84700 138000 84764 138004
rect 84700 137944 84750 138000
rect 84750 137944 84764 138000
rect 84700 137940 84764 137944
rect 193444 137940 193508 138004
rect 225276 137260 225340 137324
rect 90956 136716 91020 136780
rect 93532 136716 93596 136780
rect 65932 135900 65996 135964
rect 95188 133996 95252 134060
rect 69428 133452 69492 133516
rect 224356 131684 224420 131748
rect 98500 129236 98564 129300
rect 68140 128828 68204 128892
rect 192340 127604 192404 127668
rect 191052 125700 191116 125764
rect 193260 125700 193324 125764
rect 97948 125428 98012 125492
rect 69428 124884 69492 124948
rect 224908 121348 224972 121412
rect 226380 119444 226444 119508
rect 65932 118356 65996 118420
rect 224908 108020 224972 108084
rect 66116 106388 66180 106452
rect 100708 105844 100772 105908
rect 193812 104484 193876 104548
rect 194180 104076 194244 104140
rect 191052 99996 191116 100060
rect 94820 98500 94884 98564
rect 226380 98772 226444 98836
rect 66668 97956 66732 98020
rect 224540 97412 224604 97476
rect 94820 95508 94884 95572
rect 69428 95236 69492 95300
rect 186820 95236 186884 95300
rect 224724 94692 224788 94756
rect 69244 94420 69308 94484
rect 192340 93740 192404 93804
rect 202092 93332 202156 93396
rect 224724 93392 224788 93396
rect 224724 93336 224774 93392
rect 224774 93336 224788 93392
rect 224724 93332 224788 93336
rect 227668 93196 227732 93260
rect 210372 92984 210436 92988
rect 210372 92928 210422 92984
rect 210422 92928 210436 92984
rect 97212 92788 97276 92852
rect 210372 92924 210436 92928
rect 200620 92788 200684 92852
rect 208348 92848 208412 92852
rect 208348 92792 208398 92848
rect 208398 92792 208412 92848
rect 208348 92788 208412 92792
rect 224540 92788 224604 92852
rect 68876 92652 68940 92716
rect 71452 92652 71516 92716
rect 93716 92652 93780 92716
rect 193444 92652 193508 92716
rect 191052 92516 191116 92580
rect 72556 92380 72620 92444
rect 95188 92380 95252 92444
rect 207060 92380 207124 92444
rect 211660 92380 211724 92444
rect 72740 91020 72804 91084
rect 69244 90884 69308 90948
rect 96660 90400 96724 90404
rect 96660 90344 96710 90400
rect 96710 90344 96724 90400
rect 96660 90340 96724 90344
rect 215340 90264 215404 90268
rect 215340 90208 215354 90264
rect 215354 90208 215404 90264
rect 215340 90204 215404 90208
rect 66668 89388 66732 89452
rect 94636 89388 94700 89452
rect 192708 83404 192772 83468
rect 69612 82588 69676 82652
rect 94452 82588 94516 82652
rect 189948 82044 190012 82108
rect 193812 82044 193876 82108
rect 226380 81364 226444 81428
rect 97948 79868 98012 79932
rect 188292 77828 188356 77892
rect 196572 77828 196636 77892
rect 224908 74428 224972 74492
rect 170260 44780 170324 44844
rect 206876 32404 206940 32468
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 583166 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 583166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 75867 596324 75933 596325
rect 75867 596260 75868 596324
rect 75932 596260 75933 596324
rect 75867 596259 75933 596260
rect 75683 581092 75749 581093
rect 75683 581028 75684 581092
rect 75748 581028 75749 581092
rect 75683 581027 75749 581028
rect 71635 580820 71701 580821
rect 71635 580756 71636 580820
rect 71700 580756 71701 580820
rect 71635 580755 71701 580756
rect 72923 580820 72989 580821
rect 72923 580756 72924 580820
rect 72988 580756 72989 580820
rect 72923 580755 72989 580756
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 69427 550900 69493 550901
rect 69427 550836 69428 550900
rect 69492 550836 69493 550900
rect 69427 550835 69493 550836
rect 69430 547890 69490 550835
rect 69430 547830 69858 547890
rect 69427 543556 69493 543557
rect 69427 543492 69428 543556
rect 69492 543492 69493 543556
rect 69427 543491 69493 543492
rect 69430 538230 69490 543491
rect 69430 538170 69674 538230
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 67771 468484 67837 468485
rect 67771 468420 67772 468484
rect 67836 468420 67837 468484
rect 67771 468419 67837 468420
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66115 446452 66181 446453
rect 66115 446388 66116 446452
rect 66180 446388 66181 446452
rect 66115 446387 66181 446388
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66118 411909 66178 446387
rect 66954 436356 67574 464058
rect 67403 434620 67469 434621
rect 67403 434556 67404 434620
rect 67468 434556 67469 434620
rect 67403 434555 67469 434556
rect 66299 417484 66365 417485
rect 66299 417420 66300 417484
rect 66364 417420 66365 417484
rect 66299 417419 66365 417420
rect 66302 412997 66362 417419
rect 66299 412996 66365 412997
rect 66299 412932 66300 412996
rect 66364 412932 66365 412996
rect 66299 412931 66365 412932
rect 66115 411908 66181 411909
rect 66115 411844 66116 411908
rect 66180 411844 66181 411908
rect 66115 411843 66181 411844
rect 67406 409733 67466 434555
rect 67403 409732 67469 409733
rect 67403 409668 67404 409732
rect 67468 409668 67469 409732
rect 67403 409667 67469 409668
rect 66667 401708 66733 401709
rect 66667 401644 66668 401708
rect 66732 401644 66733 401708
rect 66667 401643 66733 401644
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 66670 369749 66730 401643
rect 67774 397493 67834 468419
rect 69614 466581 69674 538170
rect 69798 537437 69858 547830
rect 69795 537436 69861 537437
rect 69795 537372 69796 537436
rect 69860 537372 69861 537436
rect 69795 537371 69861 537372
rect 69611 466580 69677 466581
rect 69611 466516 69612 466580
rect 69676 466516 69677 466580
rect 69611 466515 69677 466516
rect 69611 443052 69677 443053
rect 69611 442988 69612 443052
rect 69676 442988 69677 443052
rect 69611 442987 69677 442988
rect 69059 434348 69125 434349
rect 69059 434284 69060 434348
rect 69124 434284 69125 434348
rect 69059 434283 69125 434284
rect 67955 433940 68021 433941
rect 67955 433876 67956 433940
rect 68020 433876 68021 433940
rect 67955 433875 68021 433876
rect 67958 422245 68018 433875
rect 67955 422244 68021 422245
rect 67955 422180 67956 422244
rect 68020 422180 68021 422244
rect 67955 422179 68021 422180
rect 67771 397492 67837 397493
rect 67771 397428 67772 397492
rect 67836 397428 67837 397492
rect 67771 397427 67837 397428
rect 66667 369748 66733 369749
rect 66667 369684 66668 369748
rect 66732 369684 66733 369748
rect 66667 369683 66733 369684
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 66954 356614 67574 388356
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66667 287740 66733 287741
rect 66667 287676 66668 287740
rect 66732 287676 66733 287740
rect 66667 287675 66733 287676
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 66670 256733 66730 287675
rect 66954 285592 67574 320058
rect 68691 283524 68757 283525
rect 68691 283460 68692 283524
rect 68756 283460 68757 283524
rect 68691 283459 68757 283460
rect 67955 280532 68021 280533
rect 67955 280468 67956 280532
rect 68020 280468 68021 280532
rect 67955 280467 68021 280468
rect 66667 256732 66733 256733
rect 66667 256668 66668 256732
rect 66732 256668 66733 256732
rect 66667 256667 66733 256668
rect 66115 255372 66181 255373
rect 66115 255308 66116 255372
rect 66180 255308 66181 255372
rect 66115 255307 66181 255308
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 65931 135964 65997 135965
rect 65931 135900 65932 135964
rect 65996 135900 65997 135964
rect 65931 135899 65997 135900
rect 65934 118421 65994 135899
rect 65931 118420 65997 118421
rect 65931 118356 65932 118420
rect 65996 118356 65997 118420
rect 65931 118355 65997 118356
rect 66118 106453 66178 255307
rect 66667 247076 66733 247077
rect 66667 247012 66668 247076
rect 66732 247012 66733 247076
rect 66667 247011 66733 247012
rect 66670 224909 66730 247011
rect 67958 241501 68018 280467
rect 67955 241500 68021 241501
rect 67955 241436 67956 241500
rect 68020 241436 68021 241500
rect 67955 241435 68021 241436
rect 66667 224908 66733 224909
rect 66667 224844 66668 224908
rect 66732 224844 66733 224908
rect 66667 224843 66733 224844
rect 66115 106452 66181 106453
rect 66115 106388 66116 106452
rect 66180 106388 66181 106452
rect 66115 106387 66181 106388
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 66670 98021 66730 224843
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 68694 165613 68754 283459
rect 69062 282845 69122 434283
rect 69614 431970 69674 442987
rect 71638 434893 71698 580755
rect 72739 520980 72805 520981
rect 72739 520916 72740 520980
rect 72804 520916 72805 520980
rect 72739 520915 72805 520916
rect 71819 436116 71885 436117
rect 71819 436052 71820 436116
rect 71884 436052 71885 436116
rect 71819 436051 71885 436052
rect 71635 434892 71701 434893
rect 71635 434828 71636 434892
rect 71700 434828 71701 434892
rect 71635 434827 71701 434828
rect 70899 433804 70965 433805
rect 70899 433740 70900 433804
rect 70964 433740 70965 433804
rect 70899 433739 70965 433740
rect 69430 431910 69674 431970
rect 69430 429861 69490 431910
rect 69427 429860 69493 429861
rect 69427 429796 69428 429860
rect 69492 429796 69493 429860
rect 69427 429795 69493 429796
rect 69427 393956 69493 393957
rect 69427 393892 69428 393956
rect 69492 393892 69493 393956
rect 69427 393891 69493 393892
rect 69430 393330 69490 393891
rect 69430 393270 69674 393330
rect 69614 375325 69674 393270
rect 69611 375324 69677 375325
rect 69611 375260 69612 375324
rect 69676 375260 69677 375324
rect 69611 375259 69677 375260
rect 70902 288421 70962 433739
rect 71822 303653 71882 436051
rect 72742 389061 72802 520915
rect 72926 464405 72986 580755
rect 73679 543454 73999 543486
rect 73679 543218 73721 543454
rect 73957 543218 73999 543454
rect 73679 543134 73999 543218
rect 73679 542898 73721 543134
rect 73957 542898 73999 543134
rect 73679 542866 73999 542898
rect 73291 537572 73357 537573
rect 73291 537508 73292 537572
rect 73356 537508 73357 537572
rect 73291 537507 73357 537508
rect 72923 464404 72989 464405
rect 72923 464340 72924 464404
rect 72988 464340 72989 464404
rect 72923 464339 72989 464340
rect 73294 441630 73354 537507
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 75686 476781 75746 581027
rect 75870 539613 75930 596259
rect 77514 583166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 583166 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 583166 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 583166 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 583166 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 83411 582452 83477 582453
rect 83411 582388 83412 582452
rect 83476 582388 83477 582452
rect 83411 582387 83477 582388
rect 79915 580820 79981 580821
rect 79915 580756 79916 580820
rect 79980 580756 79981 580820
rect 79915 580755 79981 580756
rect 77644 561454 77964 561486
rect 77644 561218 77686 561454
rect 77922 561218 77964 561454
rect 77644 561134 77964 561218
rect 77644 560898 77686 561134
rect 77922 560898 77964 561134
rect 77644 560866 77964 560898
rect 75867 539612 75933 539613
rect 75867 539548 75868 539612
rect 75932 539548 75933 539612
rect 75867 539547 75933 539548
rect 77514 511174 78134 537166
rect 79731 523700 79797 523701
rect 79731 523636 79732 523700
rect 79796 523636 79797 523700
rect 79731 523635 79797 523636
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 75683 476780 75749 476781
rect 75683 476716 75684 476780
rect 75748 476716 75749 476780
rect 75683 476715 75749 476716
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73294 441570 73538 441630
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 73478 390965 73538 441570
rect 73794 436356 74414 470898
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 436356 78134 438618
rect 73659 435436 73725 435437
rect 73659 435372 73660 435436
rect 73724 435372 73725 435436
rect 73659 435371 73725 435372
rect 73662 402990 73722 435371
rect 76419 434348 76485 434349
rect 76419 434284 76420 434348
rect 76484 434284 76485 434348
rect 76419 434283 76485 434284
rect 74579 433668 74645 433669
rect 74579 433604 74580 433668
rect 74644 433604 74645 433668
rect 74579 433603 74645 433604
rect 73662 402930 73906 402990
rect 73475 390964 73541 390965
rect 73475 390900 73476 390964
rect 73540 390900 73541 390964
rect 73475 390899 73541 390900
rect 73846 389190 73906 402930
rect 73478 389130 73906 389190
rect 72739 389060 72805 389061
rect 72739 388996 72740 389060
rect 72804 388996 72805 389060
rect 72739 388995 72805 388996
rect 71819 303652 71885 303653
rect 71819 303588 71820 303652
rect 71884 303588 71885 303652
rect 71819 303587 71885 303588
rect 70899 288420 70965 288421
rect 70899 288356 70900 288420
rect 70964 288356 70965 288420
rect 70899 288355 70965 288356
rect 70902 285837 70962 288355
rect 72923 286108 72989 286109
rect 72923 286044 72924 286108
rect 72988 286044 72989 286108
rect 72923 286043 72989 286044
rect 70899 285836 70965 285837
rect 70899 285772 70900 285836
rect 70964 285772 70965 285836
rect 70899 285771 70965 285772
rect 70899 285700 70965 285701
rect 70899 285636 70900 285700
rect 70964 285636 70965 285700
rect 70899 285635 70965 285636
rect 69243 283252 69309 283253
rect 69243 283188 69244 283252
rect 69308 283188 69309 283252
rect 69243 283187 69309 283188
rect 69059 282844 69125 282845
rect 69059 282780 69060 282844
rect 69124 282780 69125 282844
rect 69059 282779 69125 282780
rect 69246 276045 69306 283187
rect 69243 276044 69309 276045
rect 69243 275980 69244 276044
rect 69308 275980 69309 276044
rect 69243 275979 69309 275980
rect 69059 250612 69125 250613
rect 69059 250548 69060 250612
rect 69124 250548 69125 250612
rect 69059 250547 69125 250548
rect 68875 240140 68941 240141
rect 68875 240076 68876 240140
rect 68940 240076 68941 240140
rect 68875 240075 68941 240076
rect 68691 165612 68757 165613
rect 68691 165548 68692 165612
rect 68756 165548 68757 165612
rect 68691 165547 68757 165548
rect 68139 160852 68205 160853
rect 68139 160788 68140 160852
rect 68204 160788 68205 160852
rect 68139 160787 68205 160788
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 136782 67574 140058
rect 68142 128893 68202 160787
rect 68139 128892 68205 128893
rect 68139 128828 68140 128892
rect 68204 128828 68205 128892
rect 68139 128827 68205 128828
rect 66667 98020 66733 98021
rect 66667 97956 66668 98020
rect 66732 97956 66733 98020
rect 66667 97955 66733 97956
rect 66670 89453 66730 97955
rect 68878 92717 68938 240075
rect 69062 227629 69122 250547
rect 69427 244356 69493 244357
rect 69427 244292 69428 244356
rect 69492 244292 69493 244356
rect 69427 244291 69493 244292
rect 69430 238770 69490 244291
rect 70902 241773 70962 285635
rect 71635 283660 71701 283661
rect 71635 283596 71636 283660
rect 71700 283596 71701 283660
rect 71635 283595 71701 283596
rect 71638 283117 71698 283595
rect 71635 283116 71701 283117
rect 71635 283052 71636 283116
rect 71700 283052 71701 283116
rect 71635 283051 71701 283052
rect 70899 241772 70965 241773
rect 70899 241708 70900 241772
rect 70964 241708 70965 241772
rect 70899 241707 70965 241708
rect 71451 240140 71517 240141
rect 71451 240076 71452 240140
rect 71516 240076 71517 240140
rect 71451 240075 71517 240076
rect 69430 238710 69674 238770
rect 69614 235925 69674 238710
rect 69611 235924 69677 235925
rect 69611 235860 69612 235924
rect 69676 235860 69677 235924
rect 69611 235859 69677 235860
rect 69059 227628 69125 227629
rect 69059 227564 69060 227628
rect 69124 227564 69125 227628
rect 69059 227563 69125 227564
rect 69062 226949 69122 227563
rect 69059 226948 69125 226949
rect 69059 226884 69060 226948
rect 69124 226884 69125 226948
rect 69059 226883 69125 226884
rect 71454 211853 71514 240075
rect 71451 211852 71517 211853
rect 71451 211788 71452 211852
rect 71516 211788 71517 211852
rect 71451 211787 71517 211788
rect 69611 180844 69677 180845
rect 69611 180780 69612 180844
rect 69676 180780 69677 180844
rect 69611 180779 69677 180780
rect 69614 142170 69674 180779
rect 69430 142110 69674 142170
rect 69430 133517 69490 142110
rect 69795 140996 69861 140997
rect 69795 140932 69796 140996
rect 69860 140932 69861 140996
rect 69795 140931 69861 140932
rect 69427 133516 69493 133517
rect 69427 133452 69428 133516
rect 69492 133452 69493 133516
rect 69427 133451 69493 133452
rect 69798 132510 69858 140931
rect 69430 132450 69858 132510
rect 69430 124949 69490 132450
rect 69427 124948 69493 124949
rect 69427 124884 69428 124948
rect 69492 124884 69493 124948
rect 69427 124883 69493 124884
rect 69427 95300 69493 95301
rect 69427 95236 69428 95300
rect 69492 95236 69493 95300
rect 69427 95235 69493 95236
rect 69243 94484 69309 94485
rect 69243 94420 69244 94484
rect 69308 94420 69309 94484
rect 69243 94419 69309 94420
rect 68875 92716 68941 92717
rect 68875 92652 68876 92716
rect 68940 92652 68941 92716
rect 68875 92651 68941 92652
rect 69246 90949 69306 94419
rect 69430 93870 69490 95235
rect 69430 93810 69674 93870
rect 69243 90948 69309 90949
rect 69243 90884 69244 90948
rect 69308 90884 69309 90948
rect 69243 90883 69309 90884
rect 66667 89452 66733 89453
rect 66667 89388 66668 89452
rect 66732 89388 66733 89452
rect 66667 89387 66733 89388
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 90782
rect 69614 82653 69674 93810
rect 71454 92717 71514 211787
rect 71638 153101 71698 283051
rect 72371 282980 72437 282981
rect 72371 282916 72372 282980
rect 72436 282916 72437 282980
rect 72371 282915 72437 282916
rect 72374 240141 72434 282915
rect 72926 240141 72986 286043
rect 73291 283116 73357 283117
rect 73291 283052 73292 283116
rect 73356 283052 73357 283116
rect 73291 283051 73357 283052
rect 73294 240141 73354 283051
rect 73478 282981 73538 389130
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 74582 316165 74642 433603
rect 74579 316164 74645 316165
rect 74579 316100 74580 316164
rect 74644 316100 74645 316164
rect 74579 316099 74645 316100
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 285592 74414 290898
rect 76422 284885 76482 434283
rect 77339 433668 77405 433669
rect 77339 433604 77340 433668
rect 77404 433604 77405 433668
rect 77339 433603 77405 433604
rect 77342 373285 77402 433603
rect 79734 389061 79794 523635
rect 79918 437610 79978 580755
rect 81609 543454 81929 543486
rect 81609 543218 81651 543454
rect 81887 543218 81929 543454
rect 81609 543134 81929 543218
rect 81609 542898 81651 543134
rect 81887 542898 81929 543134
rect 81609 542866 81929 542898
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 83414 460189 83474 582387
rect 88379 580820 88445 580821
rect 88379 580756 88380 580820
rect 88444 580756 88445 580820
rect 88379 580755 88445 580756
rect 91691 580820 91757 580821
rect 91691 580756 91692 580820
rect 91756 580756 91757 580820
rect 91691 580755 91757 580756
rect 85575 561454 85895 561486
rect 85575 561218 85617 561454
rect 85853 561218 85895 561454
rect 85575 561134 85895 561218
rect 85575 560898 85617 561134
rect 85853 560898 85895 561134
rect 85575 560866 85895 560898
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 83411 460188 83477 460189
rect 83411 460124 83412 460188
rect 83476 460124 83477 460188
rect 83411 460123 83477 460124
rect 83595 459644 83661 459645
rect 83595 459580 83596 459644
rect 83660 459580 83661 459644
rect 83595 459579 83661 459580
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 79918 437550 80162 437610
rect 80102 389061 80162 437550
rect 81234 436356 81854 442338
rect 83598 439517 83658 459579
rect 84954 446614 85574 482058
rect 88382 449989 88442 580755
rect 89540 543454 89860 543486
rect 89540 543218 89582 543454
rect 89818 543218 89860 543454
rect 89540 543134 89860 543218
rect 89540 542898 89582 543134
rect 89818 542898 89860 543134
rect 89540 542866 89860 542898
rect 91694 537573 91754 580755
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 96659 547092 96725 547093
rect 96659 547028 96660 547092
rect 96724 547028 96725 547092
rect 96659 547027 96725 547028
rect 91691 537572 91757 537573
rect 91691 537508 91692 537572
rect 91756 537508 91757 537572
rect 91691 537507 91757 537508
rect 91794 525454 92414 537166
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 88379 449988 88445 449989
rect 88379 449924 88380 449988
rect 88444 449924 88445 449988
rect 88379 449923 88445 449924
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 83595 439516 83661 439517
rect 83595 439452 83596 439516
rect 83660 439452 83661 439516
rect 83595 439451 83661 439452
rect 83598 436117 83658 439451
rect 84954 436356 85574 446058
rect 91794 436356 92414 452898
rect 95514 529174 96134 537166
rect 96662 534717 96722 547027
rect 96659 534716 96725 534717
rect 96659 534652 96660 534716
rect 96724 534652 96725 534716
rect 96659 534651 96725 534652
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 96659 479500 96725 479501
rect 96659 479436 96660 479500
rect 96724 479436 96725 479500
rect 96659 479435 96725 479436
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 436356 96134 456618
rect 94635 436252 94701 436253
rect 94635 436188 94636 436252
rect 94700 436188 94701 436252
rect 94635 436187 94701 436188
rect 81019 436116 81085 436117
rect 81019 436052 81020 436116
rect 81084 436052 81085 436116
rect 81019 436051 81085 436052
rect 83595 436116 83661 436117
rect 83595 436052 83596 436116
rect 83660 436052 83661 436116
rect 83595 436051 83661 436052
rect 94451 436116 94517 436117
rect 94451 436052 94452 436116
rect 94516 436052 94517 436116
rect 94451 436051 94517 436052
rect 79731 389060 79797 389061
rect 79731 388996 79732 389060
rect 79796 388996 79797 389060
rect 79731 388995 79797 388996
rect 80099 389060 80165 389061
rect 80099 388996 80100 389060
rect 80164 388996 80165 389060
rect 80099 388995 80165 388996
rect 77339 373284 77405 373285
rect 77339 373220 77340 373284
rect 77404 373220 77405 373284
rect 77339 373219 77405 373220
rect 77514 367174 78134 388356
rect 81022 382941 81082 436051
rect 81939 434348 82005 434349
rect 81939 434284 81940 434348
rect 82004 434284 82005 434348
rect 81939 434283 82005 434284
rect 83043 434348 83109 434349
rect 83043 434284 83044 434348
rect 83108 434284 83109 434348
rect 83043 434283 83109 434284
rect 84699 434348 84765 434349
rect 84699 434284 84700 434348
rect 84764 434284 84765 434348
rect 84699 434283 84765 434284
rect 85803 434348 85869 434349
rect 85803 434284 85804 434348
rect 85868 434284 85869 434348
rect 85803 434283 85869 434284
rect 81019 382940 81085 382941
rect 81019 382876 81020 382940
rect 81084 382876 81085 382940
rect 81019 382875 81085 382876
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285592 78134 294618
rect 81234 370894 81854 388356
rect 81942 386205 82002 434283
rect 81939 386204 82005 386205
rect 81939 386140 81940 386204
rect 82004 386140 82005 386204
rect 81939 386139 82005 386140
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 83046 317389 83106 434283
rect 83227 434076 83293 434077
rect 83227 434012 83228 434076
rect 83292 434012 83293 434076
rect 83227 434011 83293 434012
rect 83043 317388 83109 317389
rect 83043 317324 83044 317388
rect 83108 317324 83109 317388
rect 83043 317323 83109 317324
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 285592 81854 298338
rect 83230 292637 83290 434011
rect 84702 320109 84762 434283
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84699 320108 84765 320109
rect 84699 320044 84700 320108
rect 84764 320044 84765 320108
rect 84699 320043 84765 320044
rect 84515 317388 84581 317389
rect 84515 317324 84516 317388
rect 84580 317324 84581 317388
rect 84515 317323 84581 317324
rect 83227 292636 83293 292637
rect 83227 292572 83228 292636
rect 83292 292572 83293 292636
rect 83227 292571 83293 292572
rect 76419 284884 76485 284885
rect 76419 284820 76420 284884
rect 76484 284820 76485 284884
rect 76419 284819 76485 284820
rect 83411 283252 83477 283253
rect 83411 283188 83412 283252
rect 83476 283188 83477 283252
rect 83411 283187 83477 283188
rect 73475 282980 73541 282981
rect 73475 282916 73476 282980
rect 73540 282916 73541 282980
rect 73475 282915 73541 282916
rect 72371 240140 72437 240141
rect 72371 240076 72372 240140
rect 72436 240076 72437 240140
rect 72371 240075 72437 240076
rect 72923 240140 72989 240141
rect 72923 240076 72924 240140
rect 72988 240076 72989 240140
rect 72923 240075 72989 240076
rect 73291 240140 73357 240141
rect 73291 240076 73292 240140
rect 73356 240076 73357 240140
rect 73291 240075 73357 240076
rect 72739 240004 72805 240005
rect 72739 239940 72740 240004
rect 72804 239940 72805 240004
rect 72739 239939 72805 239940
rect 72555 239868 72621 239869
rect 72555 239804 72556 239868
rect 72620 239804 72621 239868
rect 72555 239803 72621 239804
rect 71635 153100 71701 153101
rect 71635 153036 71636 153100
rect 71700 153036 71701 153100
rect 71635 153035 71701 153036
rect 71638 152149 71698 153035
rect 71635 152148 71701 152149
rect 71635 152084 71636 152148
rect 71700 152084 71701 152148
rect 71635 152083 71701 152084
rect 71451 92716 71517 92717
rect 71451 92652 71452 92716
rect 71516 92652 71517 92716
rect 71451 92651 71517 92652
rect 72558 92445 72618 239803
rect 72742 213893 72802 239939
rect 72739 213892 72805 213893
rect 72739 213828 72740 213892
rect 72804 213828 72805 213892
rect 72739 213827 72805 213828
rect 72555 92444 72621 92445
rect 72555 92380 72556 92444
rect 72620 92380 72621 92444
rect 72555 92379 72621 92380
rect 72742 91085 72802 213827
rect 73478 142357 73538 282915
rect 78977 273454 79297 273486
rect 78977 273218 79019 273454
rect 79255 273218 79297 273454
rect 78977 273134 79297 273218
rect 78977 272898 79019 273134
rect 79255 272898 79297 273134
rect 78977 272866 79297 272898
rect 74345 255454 74665 255486
rect 74345 255218 74387 255454
rect 74623 255218 74665 255454
rect 74345 255134 74665 255218
rect 74345 254898 74387 255134
rect 74623 254898 74665 255134
rect 74345 254866 74665 254898
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73475 142356 73541 142357
rect 73475 142292 73476 142356
rect 73540 142292 73541 142356
rect 73475 142291 73541 142292
rect 73478 140861 73538 142291
rect 73475 140860 73541 140861
rect 73475 140796 73476 140860
rect 73540 140796 73541 140860
rect 73475 140795 73541 140796
rect 73794 136782 74414 146898
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 136782 78134 150618
rect 81234 226894 81854 239592
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 83414 169013 83474 283187
rect 83609 255454 83929 255486
rect 83609 255218 83651 255454
rect 83887 255218 83929 255454
rect 83609 255134 83929 255218
rect 83609 254898 83651 255134
rect 83887 254898 83929 255134
rect 83609 254866 83929 254898
rect 84518 241773 84578 317323
rect 84954 302614 85574 338058
rect 85806 322829 85866 434283
rect 92979 434212 93045 434213
rect 92979 434148 92980 434212
rect 93044 434148 93045 434212
rect 92979 434147 93045 434148
rect 87091 433668 87157 433669
rect 87091 433604 87092 433668
rect 87156 433604 87157 433668
rect 87091 433603 87157 433604
rect 87459 433668 87525 433669
rect 87459 433604 87460 433668
rect 87524 433604 87525 433668
rect 87459 433603 87525 433604
rect 89667 433668 89733 433669
rect 89667 433604 89668 433668
rect 89732 433604 89733 433668
rect 89667 433603 89733 433604
rect 90035 433668 90101 433669
rect 90035 433604 90036 433668
rect 90100 433604 90101 433668
rect 90035 433603 90101 433604
rect 91323 433668 91389 433669
rect 91323 433604 91324 433668
rect 91388 433604 91389 433668
rect 91323 433603 91389 433604
rect 91507 433668 91573 433669
rect 91507 433604 91508 433668
rect 91572 433604 91573 433668
rect 91507 433603 91573 433604
rect 92795 433668 92861 433669
rect 92795 433604 92796 433668
rect 92860 433604 92861 433668
rect 92795 433603 92861 433604
rect 85803 322828 85869 322829
rect 85803 322764 85804 322828
rect 85868 322764 85869 322828
rect 85803 322763 85869 322764
rect 87094 318069 87154 433603
rect 87462 387021 87522 433603
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 87459 387020 87525 387021
rect 87459 386956 87460 387020
rect 87524 386956 87525 387020
rect 87459 386955 87525 386956
rect 87091 318068 87157 318069
rect 87091 318004 87092 318068
rect 87156 318004 87157 318068
rect 87091 318003 87157 318004
rect 89670 309909 89730 433603
rect 90038 384301 90098 433603
rect 91326 387837 91386 433603
rect 91323 387836 91389 387837
rect 91323 387772 91324 387836
rect 91388 387772 91389 387836
rect 91323 387771 91389 387772
rect 90035 384300 90101 384301
rect 90035 384236 90036 384300
rect 90100 384236 90101 384300
rect 90035 384235 90101 384236
rect 89667 309908 89733 309909
rect 89667 309844 89668 309908
rect 89732 309844 89733 309908
rect 89667 309843 89733 309844
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 285592 85574 302058
rect 91510 297533 91570 433603
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91507 297532 91573 297533
rect 91507 297468 91508 297532
rect 91572 297468 91573 297532
rect 91507 297467 91573 297468
rect 86539 291140 86605 291141
rect 86539 291076 86540 291140
rect 86604 291076 86605 291140
rect 86539 291075 86605 291076
rect 84699 283252 84765 283253
rect 84699 283188 84700 283252
rect 84764 283188 84765 283252
rect 84699 283187 84765 283188
rect 84515 241772 84581 241773
rect 84515 241708 84516 241772
rect 84580 241708 84581 241772
rect 84515 241707 84581 241708
rect 84518 238781 84578 241707
rect 84515 238780 84581 238781
rect 84515 238716 84516 238780
rect 84580 238716 84581 238780
rect 84515 238715 84581 238716
rect 83411 169012 83477 169013
rect 83411 168948 83412 169012
rect 83476 168948 83477 169012
rect 83411 168947 83477 168948
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 136782 81854 154338
rect 84702 138005 84762 283187
rect 86542 241773 86602 291075
rect 91507 289916 91573 289917
rect 91507 289852 91508 289916
rect 91572 289852 91573 289916
rect 91507 289851 91573 289852
rect 88011 289780 88077 289781
rect 88011 289716 88012 289780
rect 88076 289716 88077 289780
rect 88011 289715 88077 289716
rect 86723 283796 86789 283797
rect 86723 283732 86724 283796
rect 86788 283732 86789 283796
rect 86723 283731 86789 283732
rect 86539 241772 86605 241773
rect 86539 241708 86540 241772
rect 86604 241708 86605 241772
rect 86539 241707 86605 241708
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 86542 191045 86602 241707
rect 86539 191044 86605 191045
rect 86539 190980 86540 191044
rect 86604 190980 86605 191044
rect 86539 190979 86605 190980
rect 86726 169149 86786 283731
rect 88014 241637 88074 289715
rect 90955 288556 91021 288557
rect 90955 288492 90956 288556
rect 91020 288492 91021 288556
rect 90955 288491 91021 288492
rect 89483 283524 89549 283525
rect 89483 283460 89484 283524
rect 89548 283460 89549 283524
rect 89483 283459 89549 283460
rect 90035 283524 90101 283525
rect 90035 283460 90036 283524
rect 90100 283460 90101 283524
rect 90035 283459 90101 283460
rect 88241 273454 88561 273486
rect 88241 273218 88283 273454
rect 88519 273218 88561 273454
rect 88241 273134 88561 273218
rect 88241 272898 88283 273134
rect 88519 272898 88561 273134
rect 88241 272866 88561 272898
rect 88011 241636 88077 241637
rect 88011 241572 88012 241636
rect 88076 241572 88077 241636
rect 88011 241571 88077 241572
rect 88014 239869 88074 241571
rect 88011 239868 88077 239869
rect 88011 239804 88012 239868
rect 88076 239804 88077 239868
rect 88011 239803 88077 239804
rect 89486 175405 89546 283459
rect 90038 226405 90098 283459
rect 90958 241773 91018 288491
rect 91510 241773 91570 289851
rect 91794 285592 92414 308898
rect 92798 293317 92858 433603
rect 92795 293316 92861 293317
rect 92795 293252 92796 293316
rect 92860 293252 92861 293316
rect 92795 293251 92861 293252
rect 92982 291821 93042 434147
rect 94454 319429 94514 436051
rect 94638 383757 94698 436187
rect 96291 434348 96357 434349
rect 96291 434284 96292 434348
rect 96356 434284 96357 434348
rect 96291 434283 96357 434284
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 94635 383756 94701 383757
rect 94635 383692 94636 383756
rect 94700 383692 94701 383756
rect 94635 383691 94701 383692
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 94451 319428 94517 319429
rect 94451 319364 94452 319428
rect 94516 319364 94517 319428
rect 94451 319363 94517 319364
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 92979 291820 93045 291821
rect 92979 291756 92980 291820
rect 93044 291756 93045 291820
rect 92979 291755 93045 291756
rect 95187 285972 95253 285973
rect 95187 285908 95188 285972
rect 95252 285970 95253 285972
rect 95252 285910 95434 285970
rect 95252 285908 95253 285910
rect 95187 285907 95253 285908
rect 93899 283524 93965 283525
rect 93899 283460 93900 283524
rect 93964 283460 93965 283524
rect 93899 283459 93965 283460
rect 92873 255454 93193 255486
rect 92873 255218 92915 255454
rect 93151 255218 93193 255454
rect 92873 255134 93193 255218
rect 92873 254898 92915 255134
rect 93151 254898 93193 255134
rect 92873 254866 93193 254898
rect 90955 241772 91021 241773
rect 90955 241708 90956 241772
rect 91020 241708 91021 241772
rect 90955 241707 91021 241708
rect 91507 241772 91573 241773
rect 91507 241708 91508 241772
rect 91572 241708 91573 241772
rect 91507 241707 91573 241708
rect 90958 240141 91018 241707
rect 90955 240140 91021 240141
rect 90955 240076 90956 240140
rect 91020 240076 91021 240140
rect 90955 240075 91021 240076
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 93715 237420 93781 237421
rect 93715 237356 93716 237420
rect 93780 237356 93781 237420
rect 93715 237355 93781 237356
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 90035 226404 90101 226405
rect 90035 226340 90036 226404
rect 90100 226340 90101 226404
rect 90035 226339 90101 226340
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 89483 175404 89549 175405
rect 89483 175340 89484 175404
rect 89548 175340 89549 175404
rect 89483 175339 89549 175340
rect 90955 169828 91021 169829
rect 90955 169764 90956 169828
rect 91020 169764 91021 169828
rect 90955 169763 91021 169764
rect 86723 169148 86789 169149
rect 86723 169084 86724 169148
rect 86788 169084 86789 169148
rect 86723 169083 86789 169084
rect 86726 168469 86786 169083
rect 86723 168468 86789 168469
rect 86723 168404 86724 168468
rect 86788 168404 86789 168468
rect 86723 168403 86789 168404
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84699 138004 84765 138005
rect 84699 137940 84700 138004
rect 84764 137940 84765 138004
rect 84699 137939 84765 137940
rect 84954 136782 85574 158058
rect 90958 136781 91018 169763
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 136782 92414 164898
rect 93531 161532 93597 161533
rect 93531 161468 93532 161532
rect 93596 161468 93597 161532
rect 93531 161467 93597 161468
rect 93534 136781 93594 161467
rect 90955 136780 91021 136781
rect 90955 136716 90956 136780
rect 91020 136716 91021 136780
rect 90955 136715 91021 136716
rect 93531 136780 93597 136781
rect 93531 136716 93532 136780
rect 93596 136716 93597 136780
rect 93531 136715 93597 136716
rect 77644 129454 77964 129486
rect 77644 129218 77686 129454
rect 77922 129218 77964 129454
rect 77644 129134 77964 129218
rect 77644 128898 77686 129134
rect 77922 128898 77964 129134
rect 77644 128866 77964 128898
rect 85575 129454 85895 129486
rect 85575 129218 85617 129454
rect 85853 129218 85895 129454
rect 85575 129134 85895 129218
rect 85575 128898 85617 129134
rect 85853 128898 85895 129134
rect 85575 128866 85895 128898
rect 73679 111454 73999 111486
rect 73679 111218 73721 111454
rect 73957 111218 73999 111454
rect 73679 111134 73999 111218
rect 73679 110898 73721 111134
rect 73957 110898 73999 111134
rect 73679 110866 73999 110898
rect 81609 111454 81929 111486
rect 81609 111218 81651 111454
rect 81887 111218 81929 111454
rect 81609 111134 81929 111218
rect 81609 110898 81651 111134
rect 81887 110898 81929 111134
rect 81609 110866 81929 110898
rect 89540 111454 89860 111486
rect 89540 111218 89582 111454
rect 89818 111218 89860 111454
rect 89540 111134 89860 111218
rect 89540 110898 89582 111134
rect 89818 110898 89860 111134
rect 89540 110866 89860 110898
rect 93718 92717 93778 237355
rect 93902 227085 93962 283459
rect 95374 229110 95434 285910
rect 95514 285592 96134 312618
rect 96294 309773 96354 434283
rect 96662 390557 96722 479435
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 97211 460188 97277 460189
rect 97211 460124 97212 460188
rect 97276 460124 97277 460188
rect 97211 460123 97277 460124
rect 96659 390556 96725 390557
rect 96659 390492 96660 390556
rect 96724 390492 96725 390556
rect 96659 390491 96725 390492
rect 97214 388925 97274 460123
rect 99234 436356 99854 460338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 104939 571436 105005 571437
rect 104939 571372 104940 571436
rect 105004 571372 105005 571436
rect 104939 571371 105005 571372
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 99971 458828 100037 458829
rect 99971 458764 99972 458828
rect 100036 458764 100037 458828
rect 99971 458763 100037 458764
rect 97947 433668 98013 433669
rect 97947 433604 97948 433668
rect 98012 433604 98013 433668
rect 97947 433603 98013 433604
rect 98499 433668 98565 433669
rect 98499 433604 98500 433668
rect 98564 433604 98565 433668
rect 98499 433603 98565 433604
rect 97211 388924 97277 388925
rect 97211 388860 97212 388924
rect 97276 388860 97277 388924
rect 97211 388859 97277 388860
rect 96659 378724 96725 378725
rect 96659 378660 96660 378724
rect 96724 378660 96725 378724
rect 96659 378659 96725 378660
rect 96291 309772 96357 309773
rect 96291 309708 96292 309772
rect 96356 309708 96357 309772
rect 96291 309707 96357 309708
rect 95190 229050 95434 229110
rect 93899 227084 93965 227085
rect 93899 227020 93900 227084
rect 93964 227020 93965 227084
rect 93899 227019 93965 227020
rect 95190 220965 95250 229050
rect 95187 220964 95253 220965
rect 95187 220900 95188 220964
rect 95252 220900 95253 220964
rect 95187 220899 95253 220900
rect 95514 205174 96134 239592
rect 96662 239461 96722 378659
rect 97950 318069 98010 433603
rect 97947 318068 98013 318069
rect 97947 318004 97948 318068
rect 98012 318004 98013 318068
rect 97947 318003 98013 318004
rect 98502 293181 98562 433603
rect 99974 390421 100034 458763
rect 101259 448628 101325 448629
rect 101259 448564 101260 448628
rect 101324 448564 101325 448628
rect 101259 448563 101325 448564
rect 100523 434348 100589 434349
rect 100523 434284 100524 434348
rect 100588 434284 100589 434348
rect 100523 434283 100589 434284
rect 99971 390420 100037 390421
rect 99971 390356 99972 390420
rect 100036 390356 100037 390420
rect 99971 390355 100037 390356
rect 99234 352894 99854 388356
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 98499 293180 98565 293181
rect 98499 293116 98500 293180
rect 98564 293116 98565 293180
rect 98499 293115 98565 293116
rect 99234 285592 99854 316338
rect 100526 305285 100586 434283
rect 100707 433668 100773 433669
rect 100707 433604 100708 433668
rect 100772 433604 100773 433668
rect 100707 433603 100773 433604
rect 100710 385661 100770 433603
rect 101262 390557 101322 448563
rect 102954 436356 103574 464058
rect 102731 434620 102797 434621
rect 102731 434556 102732 434620
rect 102796 434556 102797 434620
rect 102731 434555 102797 434556
rect 101259 390556 101325 390557
rect 101259 390492 101260 390556
rect 101324 390492 101325 390556
rect 101259 390491 101325 390492
rect 100707 385660 100773 385661
rect 100707 385596 100708 385660
rect 100772 385596 100773 385660
rect 100707 385595 100773 385596
rect 101259 384300 101325 384301
rect 101259 384236 101260 384300
rect 101324 384236 101325 384300
rect 101259 384235 101325 384236
rect 100523 305284 100589 305285
rect 100523 305220 100524 305284
rect 100588 305220 100589 305284
rect 100523 305219 100589 305220
rect 100526 304197 100586 305219
rect 100523 304196 100589 304197
rect 100523 304132 100524 304196
rect 100588 304132 100589 304196
rect 100523 304131 100589 304132
rect 98499 277540 98565 277541
rect 98499 277476 98500 277540
rect 98564 277476 98565 277540
rect 98499 277475 98565 277476
rect 98131 267884 98197 267885
rect 98131 267820 98132 267884
rect 98196 267820 98197 267884
rect 98131 267819 98197 267820
rect 98134 258090 98194 267819
rect 97950 258030 98194 258090
rect 97763 240140 97829 240141
rect 97763 240076 97764 240140
rect 97828 240076 97829 240140
rect 97763 240075 97829 240076
rect 96659 239460 96725 239461
rect 96659 239396 96660 239460
rect 96724 239396 96725 239460
rect 96659 239395 96725 239396
rect 96662 238781 96722 239395
rect 96659 238780 96725 238781
rect 96659 238716 96660 238780
rect 96724 238716 96725 238780
rect 96659 238715 96725 238716
rect 97579 234020 97645 234021
rect 97579 233956 97580 234020
rect 97644 233956 97645 234020
rect 97579 233955 97645 233956
rect 97582 209790 97642 233955
rect 97766 210357 97826 240075
rect 97763 210356 97829 210357
rect 97763 210292 97764 210356
rect 97828 210292 97829 210356
rect 97763 210291 97829 210292
rect 97214 209730 97642 209790
rect 97214 205733 97274 209730
rect 97211 205732 97277 205733
rect 97211 205668 97212 205732
rect 97276 205668 97277 205732
rect 97211 205667 97277 205668
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 136782 96134 168618
rect 96659 167788 96725 167789
rect 96659 167724 96660 167788
rect 96724 167724 96725 167788
rect 96659 167723 96725 167724
rect 95187 134060 95253 134061
rect 95187 133996 95188 134060
rect 95252 133996 95253 134060
rect 95187 133995 95253 133996
rect 94819 98564 94885 98565
rect 94819 98500 94820 98564
rect 94884 98500 94885 98564
rect 94819 98499 94885 98500
rect 94822 96250 94882 98499
rect 94638 96190 94882 96250
rect 93715 92716 93781 92717
rect 93715 92652 93716 92716
rect 93780 92652 93781 92716
rect 93715 92651 93781 92652
rect 72739 91084 72805 91085
rect 72739 91020 72740 91084
rect 72804 91020 72805 91084
rect 72739 91019 72805 91020
rect 69611 82652 69677 82653
rect 69611 82588 69612 82652
rect 69676 82588 69677 82652
rect 69611 82587 69677 82588
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 90782
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 90782
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 90782
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 90782
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 90782
rect 94638 89453 94698 96190
rect 94819 95572 94885 95573
rect 94819 95508 94820 95572
rect 94884 95508 94885 95572
rect 94819 95507 94885 95508
rect 94635 89452 94701 89453
rect 94635 89388 94636 89452
rect 94700 89388 94701 89452
rect 94635 89387 94701 89388
rect 94822 84210 94882 95507
rect 95190 92445 95250 133995
rect 95187 92444 95253 92445
rect 95187 92380 95188 92444
rect 95252 92380 95253 92444
rect 95187 92379 95253 92380
rect 94454 84150 94882 84210
rect 94454 82653 94514 84150
rect 94451 82652 94517 82653
rect 94451 82588 94452 82652
rect 94516 82588 94517 82652
rect 94451 82587 94517 82588
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 90782
rect 96662 90405 96722 167723
rect 97214 92853 97274 205667
rect 97950 146437 98010 258030
rect 97947 146436 98013 146437
rect 97947 146372 97948 146436
rect 98012 146372 98013 146436
rect 97947 146371 98013 146372
rect 98502 129301 98562 277475
rect 101262 276997 101322 384235
rect 102734 329085 102794 434555
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 104942 390421 105002 571371
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 106411 534852 106477 534853
rect 106411 534788 106412 534852
rect 106476 534788 106477 534852
rect 106411 534787 106477 534788
rect 105491 433668 105557 433669
rect 105491 433604 105492 433668
rect 105556 433604 105557 433668
rect 105491 433603 105557 433604
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102731 329084 102797 329085
rect 102731 329020 102732 329084
rect 102796 329020 102797 329084
rect 102731 329019 102797 329020
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 105494 319429 105554 433603
rect 106414 390421 106474 534787
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 107699 472564 107765 472565
rect 107699 472500 107700 472564
rect 107764 472500 107765 472564
rect 107699 472499 107765 472500
rect 107702 390421 107762 472499
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 107883 438156 107949 438157
rect 107883 438092 107884 438156
rect 107948 438092 107949 438156
rect 107883 438091 107949 438092
rect 107886 390693 107946 438091
rect 109794 436356 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 115059 569260 115125 569261
rect 115059 569196 115060 569260
rect 115124 569196 115125 569260
rect 115059 569195 115125 569196
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113219 464404 113285 464405
rect 113219 464340 113220 464404
rect 113284 464340 113285 464404
rect 113219 464339 113285 464340
rect 108987 433668 109053 433669
rect 108987 433604 108988 433668
rect 109052 433604 109053 433668
rect 108987 433603 109053 433604
rect 107883 390692 107949 390693
rect 107883 390628 107884 390692
rect 107948 390628 107949 390692
rect 107883 390627 107949 390628
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 107699 390420 107765 390421
rect 107699 390356 107700 390420
rect 107764 390356 107765 390420
rect 107699 390355 107765 390356
rect 105491 319428 105557 319429
rect 105491 319364 105492 319428
rect 105556 319364 105557 319428
rect 105491 319363 105557 319364
rect 108990 309773 109050 433603
rect 112115 426596 112181 426597
rect 112115 426532 112116 426596
rect 112180 426532 112181 426596
rect 112115 426531 112181 426532
rect 112118 412650 112178 426531
rect 111750 412590 112178 412650
rect 109794 363454 110414 388356
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 108987 309772 109053 309773
rect 108987 309708 108988 309772
rect 109052 309708 109053 309772
rect 108987 309707 109053 309708
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 101259 276996 101325 276997
rect 101259 276932 101260 276996
rect 101324 276932 101325 276996
rect 101259 276931 101325 276932
rect 101259 275364 101325 275365
rect 101259 275300 101260 275364
rect 101324 275300 101325 275364
rect 101259 275299 101325 275300
rect 99971 270468 100037 270469
rect 99971 270404 99972 270468
rect 100036 270404 100037 270468
rect 99971 270403 100037 270404
rect 99234 208894 99854 239592
rect 99974 234021 100034 270403
rect 100707 252516 100773 252517
rect 100707 252452 100708 252516
rect 100772 252452 100773 252516
rect 100707 252451 100773 252452
rect 99971 234020 100037 234021
rect 99971 233956 99972 234020
rect 100036 233956 100037 234020
rect 99971 233955 100037 233956
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 98499 129300 98565 129301
rect 98499 129236 98500 129300
rect 98564 129236 98565 129300
rect 98499 129235 98565 129236
rect 97947 125492 98013 125493
rect 97947 125428 97948 125492
rect 98012 125428 98013 125492
rect 97947 125427 98013 125428
rect 97211 92852 97277 92853
rect 97211 92788 97212 92852
rect 97276 92788 97277 92852
rect 97211 92787 97277 92788
rect 96659 90404 96725 90405
rect 96659 90340 96660 90404
rect 96724 90340 96725 90404
rect 96659 90339 96725 90340
rect 97950 79933 98010 125427
rect 99234 100894 99854 136338
rect 100710 105909 100770 252451
rect 101262 250477 101322 275299
rect 101259 250476 101325 250477
rect 101259 250412 101260 250476
rect 101324 250412 101325 250476
rect 101259 250411 101325 250412
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102731 243540 102797 243541
rect 102731 243476 102732 243540
rect 102796 243476 102797 243540
rect 102731 243475 102797 243476
rect 102734 224773 102794 243475
rect 102731 224772 102797 224773
rect 102731 224708 102732 224772
rect 102796 224708 102797 224772
rect 102731 224707 102797 224708
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 100707 105908 100773 105909
rect 100707 105844 100708 105908
rect 100772 105844 100773 105908
rect 100707 105843 100773 105844
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 97947 79932 98013 79933
rect 97947 79868 97948 79932
rect 98012 79868 98013 79932
rect 97947 79867 98013 79868
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 111750 278221 111810 412590
rect 113222 397221 113282 464339
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 436356 114134 438618
rect 114323 436932 114389 436933
rect 114323 436868 114324 436932
rect 114388 436868 114389 436932
rect 114323 436867 114389 436868
rect 114326 405517 114386 436867
rect 115062 410005 115122 569195
rect 117234 550894 117854 586338
rect 115979 550764 116045 550765
rect 115979 550700 115980 550764
rect 116044 550700 116045 550764
rect 115979 550699 116045 550700
rect 115059 410004 115125 410005
rect 115059 409940 115060 410004
rect 115124 409940 115125 410004
rect 115059 409939 115125 409940
rect 114323 405516 114389 405517
rect 114323 405452 114324 405516
rect 114388 405452 114389 405516
rect 114323 405451 114389 405452
rect 113219 397220 113285 397221
rect 113219 397156 113220 397220
rect 113284 397156 113285 397220
rect 113219 397155 113285 397156
rect 112851 393548 112917 393549
rect 112851 393484 112852 393548
rect 112916 393484 112917 393548
rect 112851 393483 112917 393484
rect 112854 390693 112914 393483
rect 112851 390692 112917 390693
rect 112851 390628 112852 390692
rect 112916 390628 112917 390692
rect 112851 390627 112917 390628
rect 113514 367174 114134 388356
rect 115982 386205 116042 550699
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 115979 386204 116045 386205
rect 115979 386140 115980 386204
rect 116044 386140 116045 386204
rect 115979 386139 116045 386140
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 111747 278220 111813 278221
rect 111747 278156 111748 278220
rect 111812 278156 111813 278220
rect 111747 278155 111813 278156
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 148179 265572 148245 265573
rect 148179 265508 148180 265572
rect 148244 265508 148245 265572
rect 148179 265507 148245 265508
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 148182 182885 148242 265507
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 182884 148245 182885
rect 148179 182820 148180 182884
rect 148244 182820 148245 182884
rect 148179 182819 148245 182820
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 166211 306644 166277 306645
rect 166211 306580 166212 306644
rect 166276 306580 166277 306644
rect 166211 306579 166277 306580
rect 166214 280125 166274 306579
rect 166211 280124 166277 280125
rect 166211 280060 166212 280124
rect 166276 280060 166277 280124
rect 166211 280059 166277 280060
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 170259 248436 170325 248437
rect 170259 248372 170260 248436
rect 170324 248372 170325 248436
rect 170259 248371 170325 248372
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 170262 44845 170322 248371
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 170259 44844 170325 44845
rect 170259 44780 170260 44844
rect 170324 44780 170325 44844
rect 170259 44779 170325 44780
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 177251 415988 177317 415989
rect 177251 415924 177252 415988
rect 177316 415924 177317 415988
rect 177251 415923 177317 415924
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 177254 289101 177314 415923
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 452356 193574 482058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 195835 458284 195901 458285
rect 195835 458220 195836 458284
rect 195900 458220 195901 458284
rect 195835 458219 195901 458220
rect 193443 449716 193509 449717
rect 193443 449652 193444 449716
rect 193508 449652 193509 449716
rect 193443 449651 193509 449652
rect 193446 445637 193506 449651
rect 193443 445636 193509 445637
rect 193443 445572 193444 445636
rect 193508 445572 193509 445636
rect 193443 445571 193509 445572
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 193811 423740 193877 423741
rect 193811 423676 193812 423740
rect 193876 423676 193877 423740
rect 193811 423675 193877 423676
rect 191603 412724 191669 412725
rect 191603 412660 191604 412724
rect 191668 412660 191669 412724
rect 191603 412659 191669 412660
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 188843 400484 188909 400485
rect 188843 400420 188844 400484
rect 188908 400420 188909 400484
rect 188843 400419 188909 400420
rect 188846 373965 188906 400419
rect 188843 373964 188909 373965
rect 188843 373900 188844 373964
rect 188908 373900 188909 373964
rect 188843 373899 188909 373900
rect 188846 372877 188906 373899
rect 188843 372876 188909 372877
rect 188843 372812 188844 372876
rect 188908 372812 188909 372876
rect 188843 372811 188909 372812
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 189234 370894 189854 406338
rect 191606 379405 191666 412659
rect 191603 379404 191669 379405
rect 191603 379340 191604 379404
rect 191668 379340 191669 379404
rect 191603 379339 191669 379340
rect 191606 378997 191666 379339
rect 191603 378996 191669 378997
rect 191603 378932 191604 378996
rect 191668 378932 191669 378996
rect 191603 378931 191669 378932
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 192954 374614 193574 388356
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 191603 347036 191669 347037
rect 191603 346972 191604 347036
rect 191668 346972 191669 347036
rect 191603 346971 191669 346972
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 188475 317796 188541 317797
rect 188475 317732 188476 317796
rect 188540 317732 188541 317796
rect 188475 317731 188541 317732
rect 186819 308140 186885 308141
rect 186819 308076 186820 308140
rect 186884 308076 186885 308140
rect 186819 308075 186885 308076
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 184059 291004 184125 291005
rect 184059 290940 184060 291004
rect 184124 290940 184125 291004
rect 184059 290939 184125 290940
rect 177251 289100 177317 289101
rect 177251 289036 177252 289100
rect 177316 289036 177317 289100
rect 177251 289035 177317 289036
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 177254 255373 177314 289035
rect 177803 288556 177869 288557
rect 177803 288492 177804 288556
rect 177868 288492 177869 288556
rect 177803 288491 177869 288492
rect 177251 255372 177317 255373
rect 177251 255308 177252 255372
rect 177316 255308 177317 255372
rect 177251 255307 177317 255308
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 177806 224773 177866 288491
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 177803 224772 177869 224773
rect 177803 224708 177804 224772
rect 177868 224708 177869 224772
rect 177803 224707 177869 224708
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 219454 182414 254898
rect 184062 247621 184122 290939
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 184979 254012 185045 254013
rect 184979 253948 184980 254012
rect 185044 253948 185045 254012
rect 184979 253947 185045 253948
rect 184059 247620 184125 247621
rect 184059 247556 184060 247620
rect 184124 247556 184125 247620
rect 184059 247555 184125 247556
rect 184059 244628 184125 244629
rect 184059 244564 184060 244628
rect 184124 244564 184125 244628
rect 184059 244563 184125 244564
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 184062 186965 184122 244563
rect 184243 244492 184309 244493
rect 184243 244428 184244 244492
rect 184308 244428 184309 244492
rect 184243 244427 184309 244428
rect 184246 218653 184306 244427
rect 184243 218652 184309 218653
rect 184243 218588 184244 218652
rect 184308 218588 184309 218652
rect 184243 218587 184309 218588
rect 184982 203557 185042 253947
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 184979 203556 185045 203557
rect 184979 203492 184980 203556
rect 185044 203492 185045 203556
rect 184979 203491 185045 203492
rect 185514 187174 186134 222618
rect 186822 199341 186882 308075
rect 188291 303924 188357 303925
rect 188291 303860 188292 303924
rect 188356 303860 188357 303924
rect 188291 303859 188357 303860
rect 187003 231164 187069 231165
rect 187003 231100 187004 231164
rect 187068 231100 187069 231164
rect 187003 231099 187069 231100
rect 186819 199340 186885 199341
rect 186819 199276 186820 199340
rect 186884 199276 186885 199340
rect 186819 199275 186885 199276
rect 187006 196621 187066 231099
rect 187003 196620 187069 196621
rect 187003 196556 187004 196620
rect 187068 196556 187069 196620
rect 187003 196555 187069 196556
rect 184059 186964 184125 186965
rect 184059 186900 184060 186964
rect 184124 186900 184125 186964
rect 184059 186899 184125 186900
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 187006 180810 187066 196555
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 186822 180750 187066 180810
rect 186822 95301 186882 180750
rect 186819 95300 186885 95301
rect 186819 95236 186820 95300
rect 186884 95236 186885 95300
rect 186819 95235 186885 95236
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 188294 77893 188354 303859
rect 188478 298757 188538 317731
rect 189234 298894 189854 334338
rect 191606 306390 191666 346971
rect 192954 338614 193574 374058
rect 193814 371925 193874 423675
rect 193995 396540 194061 396541
rect 193995 396476 193996 396540
rect 194060 396476 194061 396540
rect 193995 396475 194061 396476
rect 193998 390557 194058 396475
rect 193995 390556 194061 390557
rect 193995 390492 193996 390556
rect 194060 390492 194061 390556
rect 193995 390491 194061 390492
rect 195838 381581 195898 458219
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 197123 453116 197189 453117
rect 197123 453052 197124 453116
rect 197188 453052 197189 453116
rect 197123 453051 197189 453052
rect 195835 381580 195901 381581
rect 195835 381516 195836 381580
rect 195900 381516 195901 381580
rect 195835 381515 195901 381516
rect 197126 380901 197186 453051
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 452356 200414 452898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 452356 204134 456618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 452356 207854 460338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 452356 211574 464058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 452356 218414 470898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 452356 222134 474618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 452356 225854 478338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 452356 229574 482058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 452356 236414 452898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 452356 240134 456618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 242019 452708 242085 452709
rect 242019 452644 242020 452708
rect 242084 452644 242085 452708
rect 242019 452643 242085 452644
rect 241651 449988 241717 449989
rect 241651 449924 241652 449988
rect 241716 449924 241717 449988
rect 241651 449923 241717 449924
rect 197776 435454 198096 435486
rect 197776 435218 197818 435454
rect 198054 435218 198096 435454
rect 197776 435134 198096 435218
rect 197776 434898 197818 435134
rect 198054 434898 198096 435134
rect 197776 434866 198096 434898
rect 228496 435454 228816 435486
rect 228496 435218 228538 435454
rect 228774 435218 228816 435454
rect 228496 435134 228816 435218
rect 228496 434898 228538 435134
rect 228774 434898 228816 435134
rect 228496 434866 228816 434898
rect 213136 417454 213456 417486
rect 213136 417218 213178 417454
rect 213414 417218 213456 417454
rect 213136 417134 213456 417218
rect 213136 416898 213178 417134
rect 213414 416898 213456 417134
rect 213136 416866 213456 416898
rect 197776 399454 198096 399486
rect 197776 399218 197818 399454
rect 198054 399218 198096 399454
rect 197776 399134 198096 399218
rect 197776 398898 197818 399134
rect 198054 398898 198096 399134
rect 197776 398866 198096 398898
rect 228496 399454 228816 399486
rect 228496 399218 228538 399454
rect 228774 399218 228816 399454
rect 228496 399134 228816 399218
rect 228496 398898 228538 399134
rect 228774 398898 228816 399134
rect 228496 398866 228816 398898
rect 199794 381454 200414 388356
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 197123 380900 197189 380901
rect 197123 380836 197124 380900
rect 197188 380836 197189 380900
rect 197123 380835 197189 380836
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 193811 371924 193877 371925
rect 193811 371860 193812 371924
rect 193876 371860 193877 371924
rect 193811 371859 193877 371860
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192523 306508 192589 306509
rect 192523 306444 192524 306508
rect 192588 306444 192589 306508
rect 192523 306443 192589 306444
rect 191606 306330 191850 306390
rect 189947 303788 190013 303789
rect 189947 303724 189948 303788
rect 190012 303724 190013 303788
rect 189947 303723 190013 303724
rect 188475 298756 188541 298757
rect 188475 298692 188476 298756
rect 188540 298692 188541 298756
rect 188475 298691 188541 298692
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 188291 77892 188357 77893
rect 188291 77828 188292 77892
rect 188356 77828 188357 77892
rect 188291 77827 188357 77828
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 82338
rect 189950 82109 190010 303723
rect 191603 300932 191669 300933
rect 191603 300868 191604 300932
rect 191668 300868 191669 300932
rect 191603 300867 191669 300868
rect 191606 297533 191666 300867
rect 191603 297532 191669 297533
rect 191603 297468 191604 297532
rect 191668 297468 191669 297532
rect 191603 297467 191669 297468
rect 191790 294405 191850 306330
rect 192339 301476 192405 301477
rect 192339 301412 192340 301476
rect 192404 301412 192405 301476
rect 192339 301411 192405 301412
rect 192342 294541 192402 301411
rect 192339 294540 192405 294541
rect 192339 294476 192340 294540
rect 192404 294476 192405 294540
rect 192339 294475 192405 294476
rect 191787 294404 191853 294405
rect 191787 294340 191788 294404
rect 191852 294340 191853 294404
rect 191787 294339 191853 294340
rect 191790 292365 191850 294339
rect 191787 292364 191853 292365
rect 191787 292300 191788 292364
rect 191852 292300 191853 292364
rect 191787 292299 191853 292300
rect 191051 290052 191117 290053
rect 191051 289988 191052 290052
rect 191116 289988 191117 290052
rect 191051 289987 191117 289988
rect 191054 160717 191114 289987
rect 192526 288421 192586 306443
rect 192954 303592 193574 338058
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 197123 303652 197189 303653
rect 197123 303588 197124 303652
rect 197188 303588 197189 303652
rect 199794 303592 200414 308898
rect 203514 385174 204134 388356
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 303592 204134 312618
rect 207234 352894 207854 388356
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 303592 207854 316338
rect 210954 356614 211574 388356
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 303592 211574 320058
rect 217794 363454 218414 388356
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 303592 218414 326898
rect 221514 367174 222134 388356
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 303592 222134 330618
rect 225234 370894 225854 388356
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 303592 225854 334338
rect 228954 374614 229574 388356
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 303592 229574 338058
rect 235794 381454 236414 388356
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 303592 236414 308898
rect 239514 385174 240134 388356
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 241654 366485 241714 449923
rect 242022 371381 242082 452643
rect 243234 452356 243854 460338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 244779 454068 244845 454069
rect 244779 454004 244780 454068
rect 244844 454004 244845 454068
rect 244779 454003 244845 454004
rect 243856 417454 244176 417486
rect 243856 417218 243898 417454
rect 244134 417218 244176 417454
rect 243856 417134 244176 417218
rect 243856 416898 243898 417134
rect 244134 416898 244176 417134
rect 243856 416866 244176 416898
rect 242019 371380 242085 371381
rect 242019 371316 242020 371380
rect 242084 371316 242085 371380
rect 242019 371315 242085 371316
rect 241651 366484 241717 366485
rect 241651 366420 241652 366484
rect 241716 366420 241717 366484
rect 241651 366419 241717 366420
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 243234 352894 243854 388356
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 241651 344316 241717 344317
rect 241651 344252 241652 344316
rect 241716 344252 241717 344316
rect 241651 344251 241717 344252
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 303592 240134 312618
rect 197123 303587 197189 303588
rect 193443 301204 193509 301205
rect 193443 301140 193444 301204
rect 193508 301140 193509 301204
rect 193443 301139 193509 301140
rect 193259 301068 193325 301069
rect 193259 301004 193260 301068
rect 193324 301004 193325 301068
rect 193259 301003 193325 301004
rect 193262 297397 193322 301003
rect 193259 297396 193325 297397
rect 193259 297332 193260 297396
rect 193324 297332 193325 297396
rect 193259 297331 193325 297332
rect 193446 293181 193506 301139
rect 194547 300932 194613 300933
rect 194547 300868 194548 300932
rect 194612 300868 194613 300932
rect 194547 300867 194613 300868
rect 193811 297532 193877 297533
rect 193811 297468 193812 297532
rect 193876 297468 193877 297532
rect 193811 297467 193877 297468
rect 193443 293180 193509 293181
rect 193443 293116 193444 293180
rect 193508 293116 193509 293180
rect 193443 293115 193509 293116
rect 193443 292772 193509 292773
rect 193443 292708 193444 292772
rect 193508 292708 193509 292772
rect 193443 292707 193509 292708
rect 192707 288964 192773 288965
rect 192707 288900 192708 288964
rect 192772 288900 192773 288964
rect 192707 288899 192773 288900
rect 192523 288420 192589 288421
rect 192523 288356 192524 288420
rect 192588 288356 192589 288420
rect 192523 288355 192589 288356
rect 192339 287876 192405 287877
rect 192339 287812 192340 287876
rect 192404 287812 192405 287876
rect 192339 287811 192405 287812
rect 191235 258772 191301 258773
rect 191235 258708 191236 258772
rect 191300 258708 191301 258772
rect 191235 258707 191301 258708
rect 191238 231845 191298 258707
rect 192342 239869 192402 287811
rect 192339 239868 192405 239869
rect 192339 239804 192340 239868
rect 192404 239804 192405 239868
rect 192339 239803 192405 239804
rect 192710 233885 192770 288899
rect 193446 242861 193506 292707
rect 193443 242860 193509 242861
rect 193443 242796 193444 242860
rect 193508 242796 193509 242860
rect 193443 242795 193509 242796
rect 192707 233884 192773 233885
rect 192707 233820 192708 233884
rect 192772 233820 192773 233884
rect 192707 233819 192773 233820
rect 191235 231844 191301 231845
rect 191235 231780 191236 231844
rect 191300 231780 191301 231844
rect 191235 231779 191301 231780
rect 192954 230614 193574 239592
rect 193814 235245 193874 297467
rect 194550 289830 194610 300867
rect 193998 289770 194610 289830
rect 193998 280170 194058 289770
rect 194179 283388 194245 283389
rect 194179 283324 194180 283388
rect 194244 283324 194245 283388
rect 194179 283323 194245 283324
rect 194182 281890 194242 283323
rect 197126 281890 197186 303587
rect 241654 301069 241714 344251
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 303592 243854 316338
rect 244782 304605 244842 454003
rect 246954 452356 247574 464058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 247723 457060 247789 457061
rect 247723 456996 247724 457060
rect 247788 456996 247789 457060
rect 247723 456995 247789 456996
rect 245699 449716 245765 449717
rect 245699 449652 245700 449716
rect 245764 449652 245765 449716
rect 245699 449651 245765 449652
rect 245702 361725 245762 449651
rect 245699 361724 245765 361725
rect 245699 361660 245700 361724
rect 245764 361660 245765 361724
rect 245699 361659 245765 361660
rect 246954 356614 247574 388356
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 244779 304604 244845 304605
rect 244779 304540 244780 304604
rect 244844 304540 244845 304604
rect 244779 304539 244845 304540
rect 246954 303592 247574 320058
rect 247726 303653 247786 456995
rect 252691 455700 252757 455701
rect 252691 455636 252692 455700
rect 252756 455636 252757 455700
rect 252691 455635 252757 455636
rect 248459 449988 248525 449989
rect 248459 449924 248460 449988
rect 248524 449924 248525 449988
rect 248459 449923 248525 449924
rect 248462 389877 248522 449923
rect 248459 389876 248525 389877
rect 248459 389812 248460 389876
rect 248524 389812 248525 389876
rect 248459 389811 248525 389812
rect 252507 373284 252573 373285
rect 252507 373220 252508 373284
rect 252572 373220 252573 373284
rect 252507 373219 252573 373220
rect 250299 345676 250365 345677
rect 250299 345612 250300 345676
rect 250364 345612 250365 345676
rect 250299 345611 250365 345612
rect 247723 303652 247789 303653
rect 247723 303588 247724 303652
rect 247788 303588 247789 303652
rect 247723 303587 247789 303588
rect 241651 301068 241717 301069
rect 241651 301004 241652 301068
rect 241716 301004 241717 301068
rect 241651 301003 241717 301004
rect 197307 300932 197373 300933
rect 197307 300868 197308 300932
rect 197372 300868 197373 300932
rect 197307 300867 197373 300868
rect 197310 300117 197370 300867
rect 250302 300253 250362 345611
rect 250299 300252 250365 300253
rect 250299 300188 250300 300252
rect 250364 300188 250365 300252
rect 250299 300187 250365 300188
rect 197307 300116 197373 300117
rect 197307 300052 197308 300116
rect 197372 300052 197373 300116
rect 197307 300051 197373 300052
rect 197776 291454 198096 291486
rect 197776 291218 197818 291454
rect 198054 291218 198096 291454
rect 197776 291134 198096 291218
rect 197776 290898 197818 291134
rect 198054 290898 198096 291134
rect 197776 290866 198096 290898
rect 228496 291454 228816 291486
rect 228496 291218 228538 291454
rect 228774 291218 228816 291454
rect 228496 291134 228816 291218
rect 228496 290898 228538 291134
rect 228774 290898 228816 291134
rect 228496 290866 228816 290898
rect 194182 281830 197186 281890
rect 193998 280110 194794 280170
rect 194734 273270 194794 280110
rect 194550 273210 194794 273270
rect 193811 235244 193877 235245
rect 193811 235180 193812 235244
rect 193876 235180 193877 235244
rect 193811 235179 193877 235180
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 194550 221509 194610 273210
rect 195835 242044 195901 242045
rect 195835 241980 195836 242044
rect 195900 241980 195901 242044
rect 195835 241979 195901 241980
rect 194547 221508 194613 221509
rect 194547 221444 194548 221508
rect 194612 221444 194613 221508
rect 194547 221443 194613 221444
rect 195838 202333 195898 241979
rect 197126 217429 197186 281830
rect 213136 273454 213456 273486
rect 213136 273218 213178 273454
rect 213414 273218 213456 273454
rect 213136 273134 213456 273218
rect 213136 272898 213178 273134
rect 213414 272898 213456 273134
rect 213136 272866 213456 272898
rect 243856 273454 244176 273486
rect 243856 273218 243898 273454
rect 244134 273218 244176 273454
rect 243856 273134 244176 273218
rect 243856 272898 243898 273134
rect 244134 272898 244176 273134
rect 243856 272866 244176 272898
rect 252510 267750 252570 373219
rect 252694 366349 252754 455635
rect 253794 452356 254414 470898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 254531 452708 254597 452709
rect 254531 452644 254532 452708
rect 254596 452644 254597 452708
rect 254531 452643 254597 452644
rect 252691 366348 252757 366349
rect 252691 366284 252692 366348
rect 252756 366284 252757 366348
rect 252691 366283 252757 366284
rect 253794 363454 254414 388356
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 254534 328405 254594 452643
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 256003 398036 256069 398037
rect 256003 397972 256004 398036
rect 256068 397972 256069 398036
rect 256003 397971 256069 397972
rect 255819 377364 255885 377365
rect 255819 377300 255820 377364
rect 255884 377300 255885 377364
rect 255819 377299 255885 377300
rect 254531 328404 254597 328405
rect 254531 328340 254532 328404
rect 254596 328340 254597 328404
rect 254531 328339 254597 328340
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 303592 254414 326898
rect 254531 301612 254597 301613
rect 254531 301548 254532 301612
rect 254596 301548 254597 301612
rect 254531 301547 254597 301548
rect 252510 267690 252938 267750
rect 197776 255454 198096 255486
rect 197776 255218 197818 255454
rect 198054 255218 198096 255454
rect 197776 255134 198096 255218
rect 197776 254898 197818 255134
rect 198054 254898 198096 255134
rect 197776 254866 198096 254898
rect 228496 255454 228816 255486
rect 228496 255218 228538 255454
rect 228774 255218 228816 255454
rect 228496 255134 228816 255218
rect 228496 254898 228538 255134
rect 228774 254898 228816 255134
rect 228496 254866 228816 254898
rect 252878 254013 252938 267690
rect 254534 257549 254594 301547
rect 255822 257957 255882 377299
rect 256006 369749 256066 397971
rect 256003 369748 256069 369749
rect 256003 369684 256004 369748
rect 256068 369684 256069 369748
rect 256003 369683 256069 369684
rect 257514 367174 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 262259 462364 262325 462365
rect 262259 462300 262260 462364
rect 262324 462300 262325 462364
rect 262259 462299 262325 462300
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 262262 436933 262322 462299
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 262259 436932 262325 436933
rect 262259 436868 262260 436932
rect 262324 436868 262325 436932
rect 262259 436867 262325 436868
rect 263363 436932 263429 436933
rect 263363 436868 263364 436932
rect 263428 436868 263429 436932
rect 263363 436867 263429 436868
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 258395 385660 258461 385661
rect 258395 385596 258396 385660
rect 258460 385596 258461 385660
rect 258395 385595 258461 385596
rect 258398 374010 258458 385595
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257291 305148 257357 305149
rect 257291 305084 257292 305148
rect 257356 305084 257357 305148
rect 257291 305083 257357 305084
rect 257294 278085 257354 305083
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257291 278084 257357 278085
rect 257291 278020 257292 278084
rect 257356 278020 257357 278084
rect 257291 278019 257357 278020
rect 257514 259174 258134 294618
rect 258214 373950 258458 374010
rect 258214 358730 258274 373950
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 258395 358732 258461 358733
rect 258395 358730 258396 358732
rect 258214 358670 258396 358730
rect 258214 285290 258274 358670
rect 258395 358668 258396 358670
rect 258460 358668 258461 358732
rect 258395 358667 258461 358668
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 259499 323644 259565 323645
rect 259499 323580 259500 323644
rect 259564 323580 259565 323644
rect 259499 323579 259565 323580
rect 258395 315348 258461 315349
rect 258395 315284 258396 315348
rect 258460 315284 258461 315348
rect 258395 315283 258461 315284
rect 258398 305149 258458 315283
rect 258395 305148 258461 305149
rect 258395 305084 258396 305148
rect 258460 305084 258461 305148
rect 258395 305083 258461 305084
rect 258395 302836 258461 302837
rect 258395 302772 258396 302836
rect 258460 302772 258461 302836
rect 258395 302771 258461 302772
rect 258398 289833 258458 302771
rect 258395 289832 258461 289833
rect 258395 289768 258396 289832
rect 258460 289768 258461 289832
rect 258395 289767 258461 289768
rect 259502 289645 259562 323579
rect 260971 309772 261037 309773
rect 260971 309708 260972 309772
rect 261036 309708 261037 309772
rect 260971 309707 261037 309708
rect 259683 303652 259749 303653
rect 259683 303588 259684 303652
rect 259748 303588 259749 303652
rect 259683 303587 259749 303588
rect 259686 298077 259746 303587
rect 259683 298076 259749 298077
rect 259683 298012 259684 298076
rect 259748 298012 259749 298076
rect 259683 298011 259749 298012
rect 259499 289644 259565 289645
rect 259499 289580 259500 289644
rect 259564 289580 259565 289644
rect 259499 289579 259565 289580
rect 258214 285230 258642 285290
rect 258395 285020 258461 285021
rect 258395 284956 258396 285020
rect 258460 284956 258461 285020
rect 258395 284955 258461 284956
rect 258398 263610 258458 284955
rect 258582 275229 258642 285230
rect 258579 275228 258645 275229
rect 258579 275164 258580 275228
rect 258644 275164 258645 275228
rect 258579 275163 258645 275164
rect 258398 263550 258826 263610
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 255819 257956 255885 257957
rect 255819 257892 255820 257956
rect 255884 257892 255885 257956
rect 255819 257891 255885 257892
rect 254531 257548 254597 257549
rect 254531 257484 254532 257548
rect 254596 257484 254597 257548
rect 254531 257483 254597 257484
rect 252875 254012 252941 254013
rect 252875 253948 252876 254012
rect 252940 253948 252941 254012
rect 252875 253947 252941 253948
rect 253611 243676 253677 243677
rect 253611 243612 253612 243676
rect 253676 243612 253677 243676
rect 253611 243611 253677 243612
rect 248459 242044 248525 242045
rect 248459 241980 248460 242044
rect 248524 241980 248525 242044
rect 248459 241979 248525 241980
rect 199794 237454 200414 239592
rect 200619 238100 200685 238101
rect 200619 238036 200620 238100
rect 200684 238036 200685 238100
rect 200619 238035 200685 238036
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 197123 217428 197189 217429
rect 197123 217364 197124 217428
rect 197188 217364 197189 217428
rect 197123 217363 197189 217364
rect 195835 202332 195901 202333
rect 195835 202268 195836 202332
rect 195900 202268 195901 202332
rect 195835 202267 195901 202268
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 191051 160716 191117 160717
rect 191051 160652 191052 160716
rect 191116 160652 191117 160716
rect 191051 160651 191117 160652
rect 191054 125765 191114 160651
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 143035 193574 158058
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 194363 157996 194429 157997
rect 194363 157932 194364 157996
rect 194428 157932 194429 157996
rect 194363 157931 194429 157932
rect 193075 141132 193141 141133
rect 193075 141068 193076 141132
rect 193140 141068 193141 141132
rect 193075 141067 193141 141068
rect 193078 139093 193138 141067
rect 193443 140180 193509 140181
rect 193443 140116 193444 140180
rect 193508 140116 193509 140180
rect 193443 140115 193509 140116
rect 193075 139092 193141 139093
rect 193075 139028 193076 139092
rect 193140 139028 193141 139092
rect 193075 139027 193141 139028
rect 192707 138276 192773 138277
rect 192707 138212 192708 138276
rect 192772 138212 192773 138276
rect 192707 138211 192773 138212
rect 192339 127668 192405 127669
rect 192339 127604 192340 127668
rect 192404 127604 192405 127668
rect 192339 127603 192405 127604
rect 191051 125764 191117 125765
rect 191051 125700 191052 125764
rect 191116 125700 191117 125764
rect 191051 125699 191117 125700
rect 191051 100060 191117 100061
rect 191051 99996 191052 100060
rect 191116 99996 191117 100060
rect 191051 99995 191117 99996
rect 191054 92581 191114 99995
rect 192342 93805 192402 127603
rect 192339 93804 192405 93805
rect 192339 93740 192340 93804
rect 192404 93740 192405 93804
rect 192339 93739 192405 93740
rect 191051 92580 191117 92581
rect 191051 92516 191052 92580
rect 191116 92516 191117 92580
rect 191051 92515 191117 92516
rect 192710 83469 192770 138211
rect 193446 138005 193506 140115
rect 193443 138004 193509 138005
rect 193443 137940 193444 138004
rect 193508 137940 193509 138004
rect 193443 137939 193509 137940
rect 193259 125764 193325 125765
rect 193259 125700 193260 125764
rect 193324 125700 193325 125764
rect 193259 125699 193325 125700
rect 193262 113190 193322 125699
rect 194366 113190 194426 157931
rect 196571 143444 196637 143445
rect 196571 143380 196572 143444
rect 196636 143380 196637 143444
rect 196571 143379 196637 143380
rect 196574 142357 196634 143379
rect 199794 143035 200414 164898
rect 196571 142356 196637 142357
rect 196571 142292 196572 142356
rect 196636 142292 196637 142356
rect 196571 142291 196637 142292
rect 196574 140453 196634 142291
rect 196571 140452 196637 140453
rect 196571 140388 196572 140452
rect 196636 140388 196637 140452
rect 196571 140387 196637 140388
rect 193262 113130 193506 113190
rect 193446 92717 193506 113130
rect 194182 113130 194426 113190
rect 193811 104548 193877 104549
rect 193811 104484 193812 104548
rect 193876 104484 193877 104548
rect 193811 104483 193877 104484
rect 193443 92716 193509 92717
rect 193443 92652 193444 92716
rect 193508 92652 193509 92716
rect 193443 92651 193509 92652
rect 192954 86614 193574 90782
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192707 83468 192773 83469
rect 192707 83404 192708 83468
rect 192772 83404 192773 83468
rect 192707 83403 192773 83404
rect 189947 82108 190013 82109
rect 189947 82044 189948 82108
rect 190012 82044 190013 82108
rect 189947 82043 190013 82044
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 86058
rect 193814 82109 193874 104483
rect 194182 104141 194242 113130
rect 194179 104140 194245 104141
rect 194179 104076 194180 104140
rect 194244 104076 194245 104140
rect 194179 104075 194245 104076
rect 193811 82108 193877 82109
rect 193811 82044 193812 82108
rect 193876 82044 193877 82108
rect 193811 82043 193877 82044
rect 196574 77893 196634 140387
rect 199388 111454 199708 111486
rect 199388 111218 199430 111454
rect 199666 111218 199708 111454
rect 199388 111134 199708 111218
rect 199388 110898 199430 111134
rect 199666 110898 199708 111134
rect 199388 110866 199708 110898
rect 200622 92853 200682 238035
rect 202091 214708 202157 214709
rect 202091 214644 202092 214708
rect 202156 214644 202157 214708
rect 202091 214643 202157 214644
rect 202094 93397 202154 214643
rect 203514 205174 204134 239592
rect 207059 233884 207125 233885
rect 207059 233820 207060 233884
rect 207124 233820 207125 233884
rect 207059 233819 207125 233820
rect 207062 233069 207122 233819
rect 207059 233068 207125 233069
rect 207059 233004 207060 233068
rect 207124 233004 207125 233068
rect 207059 233003 207125 233004
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 143035 204134 168618
rect 206875 140452 206941 140453
rect 206875 140388 206876 140452
rect 206940 140388 206941 140452
rect 206875 140387 206941 140388
rect 204264 129454 204584 129486
rect 204264 129218 204306 129454
rect 204542 129218 204584 129454
rect 204264 129134 204584 129218
rect 204264 128898 204306 129134
rect 204542 128898 204584 129134
rect 204264 128866 204584 128898
rect 202091 93396 202157 93397
rect 202091 93332 202092 93396
rect 202156 93332 202157 93396
rect 202091 93331 202157 93332
rect 200619 92852 200685 92853
rect 200619 92788 200620 92852
rect 200684 92788 200685 92852
rect 200619 92787 200685 92788
rect 196571 77892 196637 77893
rect 196571 77828 196572 77892
rect 196636 77828 196637 77892
rect 196571 77827 196637 77828
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 90782
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 90782
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 206878 32469 206938 140387
rect 207062 92445 207122 233003
rect 207234 208894 207854 239592
rect 208347 236604 208413 236605
rect 208347 236540 208348 236604
rect 208412 236540 208413 236604
rect 208347 236539 208413 236540
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 143035 207854 172338
rect 208350 92853 208410 236539
rect 210954 212614 211574 239592
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210371 208996 210437 208997
rect 210371 208932 210372 208996
rect 210436 208932 210437 208996
rect 210371 208931 210437 208932
rect 209140 111454 209460 111486
rect 209140 111218 209182 111454
rect 209418 111218 209460 111454
rect 209140 111134 209460 111218
rect 209140 110898 209182 111134
rect 209418 110898 209460 111134
rect 209140 110866 209460 110898
rect 210374 92989 210434 208931
rect 210954 176614 211574 212058
rect 217794 219454 218414 239592
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 215339 189140 215405 189141
rect 215339 189076 215340 189140
rect 215404 189076 215405 189140
rect 215339 189075 215405 189076
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 143035 211574 176058
rect 211659 175948 211725 175949
rect 211659 175884 211660 175948
rect 211724 175884 211725 175948
rect 211659 175883 211725 175884
rect 210371 92988 210437 92989
rect 210371 92924 210372 92988
rect 210436 92924 210437 92988
rect 210371 92923 210437 92924
rect 208347 92852 208413 92853
rect 208347 92788 208348 92852
rect 208412 92788 208413 92852
rect 208347 92787 208413 92788
rect 211662 92445 211722 175883
rect 214016 129454 214336 129486
rect 214016 129218 214058 129454
rect 214294 129218 214336 129454
rect 214016 129134 214336 129218
rect 214016 128898 214058 129134
rect 214294 128898 214336 129134
rect 214016 128866 214336 128898
rect 207059 92444 207125 92445
rect 207059 92380 207060 92444
rect 207124 92380 207125 92444
rect 207059 92379 207125 92380
rect 211659 92444 211725 92445
rect 211659 92380 211660 92444
rect 211724 92380 211725 92444
rect 211659 92379 211725 92380
rect 207234 64894 207854 90782
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 206875 32468 206941 32469
rect 206875 32404 206876 32468
rect 206940 32404 206941 32468
rect 206875 32403 206941 32404
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 68614 211574 90782
rect 215342 90269 215402 189075
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 143035 218414 146898
rect 221514 223174 222134 239592
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 225234 226894 225854 239592
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 222331 167788 222397 167789
rect 222331 167724 222332 167788
rect 222396 167724 222397 167788
rect 222331 167723 222397 167724
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 143035 222134 150618
rect 222334 140181 222394 167723
rect 225234 154894 225854 190338
rect 228954 230614 229574 239592
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 227667 167652 227733 167653
rect 227667 167588 227668 167652
rect 227732 167588 227733 167652
rect 227667 167587 227733 167588
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 224907 149700 224973 149701
rect 224907 149636 224908 149700
rect 224972 149636 224973 149700
rect 224907 149635 224973 149636
rect 224355 142220 224421 142221
rect 224355 142156 224356 142220
rect 224420 142156 224421 142220
rect 224355 142155 224421 142156
rect 222331 140180 222397 140181
rect 222331 140116 222332 140180
rect 222396 140116 222397 140180
rect 222331 140115 222397 140116
rect 224358 131749 224418 142155
rect 224355 131748 224421 131749
rect 224355 131684 224356 131748
rect 224420 131684 224421 131748
rect 224355 131683 224421 131684
rect 224910 121413 224970 149635
rect 225234 143035 225854 154338
rect 226379 146300 226445 146301
rect 226379 146236 226380 146300
rect 226444 146236 226445 146300
rect 226379 146235 226445 146236
rect 225275 140452 225341 140453
rect 225275 140388 225276 140452
rect 225340 140388 225341 140452
rect 225275 140387 225341 140388
rect 225278 137325 225338 140387
rect 225275 137324 225341 137325
rect 225275 137260 225276 137324
rect 225340 137260 225341 137324
rect 225275 137259 225341 137260
rect 224907 121412 224973 121413
rect 224907 121348 224908 121412
rect 224972 121348 224973 121412
rect 224907 121347 224973 121348
rect 226382 119509 226442 146235
rect 226563 145076 226629 145077
rect 226563 145012 226564 145076
rect 226628 145012 226629 145076
rect 226563 145011 226629 145012
rect 226566 139909 226626 145011
rect 226563 139908 226629 139909
rect 226563 139844 226564 139908
rect 226628 139844 226629 139908
rect 226563 139843 226629 139844
rect 226379 119508 226445 119509
rect 226379 119444 226380 119508
rect 226444 119444 226445 119508
rect 226379 119443 226445 119444
rect 218892 111454 219212 111486
rect 218892 111218 218934 111454
rect 219170 111218 219212 111454
rect 218892 111134 219212 111218
rect 218892 110898 218934 111134
rect 219170 110898 219212 111134
rect 218892 110866 219212 110898
rect 224907 108084 224973 108085
rect 224907 108020 224908 108084
rect 224972 108020 224973 108084
rect 224907 108019 224973 108020
rect 224539 97476 224605 97477
rect 224539 97412 224540 97476
rect 224604 97412 224605 97476
rect 224539 97411 224605 97412
rect 224542 92853 224602 97411
rect 224723 94756 224789 94757
rect 224723 94692 224724 94756
rect 224788 94692 224789 94756
rect 224723 94691 224789 94692
rect 224726 93397 224786 94691
rect 224723 93396 224789 93397
rect 224723 93332 224724 93396
rect 224788 93332 224789 93396
rect 224723 93331 224789 93332
rect 224539 92852 224605 92853
rect 224539 92788 224540 92852
rect 224604 92788 224605 92852
rect 224539 92787 224605 92788
rect 215339 90268 215405 90269
rect 215339 90204 215340 90268
rect 215404 90204 215405 90268
rect 215339 90203 215405 90204
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 90782
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 90782
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 224910 74493 224970 108019
rect 226379 98836 226445 98837
rect 226379 98772 226380 98836
rect 226444 98772 226445 98836
rect 226379 98771 226445 98772
rect 225234 82894 225854 90782
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 224907 74492 224973 74493
rect 224907 74428 224908 74492
rect 224972 74428 224973 74492
rect 224907 74427 224973 74428
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 82338
rect 226382 81429 226442 98771
rect 227670 93261 227730 167587
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 227667 93260 227733 93261
rect 227667 93196 227668 93260
rect 227732 93196 227733 93260
rect 227667 93195 227733 93196
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 226379 81428 226445 81429
rect 226379 81364 226380 81428
rect 226444 81364 226445 81428
rect 226379 81363 226445 81364
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 237454 236414 239592
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 205174 240134 239592
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 208894 243854 239592
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 212614 247574 239592
rect 248462 235245 248522 241979
rect 253614 238770 253674 243611
rect 253062 238710 253674 238770
rect 248459 235244 248525 235245
rect 248459 235180 248460 235244
rect 248524 235180 248525 235244
rect 248459 235179 248525 235180
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 253062 202197 253122 238710
rect 253794 219454 254414 239592
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253059 202196 253125 202197
rect 253059 202132 253060 202196
rect 253124 202132 253125 202196
rect 253059 202131 253125 202132
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 223174 258134 258618
rect 258214 260750 258458 260810
rect 258214 238770 258274 260750
rect 258398 260541 258458 260750
rect 258395 260540 258461 260541
rect 258395 260476 258396 260540
rect 258460 260476 258461 260540
rect 258395 260475 258461 260476
rect 258766 258770 258826 263550
rect 258398 258710 258826 258770
rect 258398 247757 258458 258710
rect 258395 247756 258461 247757
rect 258395 247692 258396 247756
rect 258460 247692 258461 247756
rect 258395 247691 258461 247692
rect 258398 240277 258458 247691
rect 258395 240276 258461 240277
rect 258395 240212 258396 240276
rect 258460 240212 258461 240276
rect 258395 240211 258461 240212
rect 258214 238710 258458 238770
rect 258398 235925 258458 238710
rect 258395 235924 258461 235925
rect 258395 235860 258396 235924
rect 258460 235860 258461 235924
rect 258395 235859 258461 235860
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 259502 146981 259562 289579
rect 260974 264485 261034 309707
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 260971 264484 261037 264485
rect 260971 264420 260972 264484
rect 261036 264420 261037 264484
rect 260971 264419 261037 264420
rect 260971 264348 261037 264349
rect 260971 264284 260972 264348
rect 261036 264284 261037 264348
rect 260971 264283 261037 264284
rect 259683 257956 259749 257957
rect 259683 257892 259684 257956
rect 259748 257892 259749 257956
rect 259683 257891 259749 257892
rect 259686 239461 259746 257891
rect 259683 239460 259749 239461
rect 259683 239396 259684 239460
rect 259748 239396 259749 239460
rect 259683 239395 259749 239396
rect 260974 214709 261034 264283
rect 261234 262894 261854 298338
rect 262259 264212 262325 264213
rect 262259 264148 262260 264212
rect 262324 264148 262325 264212
rect 262259 264147 262325 264148
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 262262 259997 262322 264147
rect 263179 261628 263245 261629
rect 263179 261564 263180 261628
rect 263244 261564 263245 261628
rect 263179 261563 263245 261564
rect 262259 259996 262325 259997
rect 262259 259932 262260 259996
rect 262324 259932 262325 259996
rect 262259 259931 262325 259932
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 260971 214708 261037 214709
rect 260971 214644 260972 214708
rect 261036 214644 261037 214708
rect 260971 214643 261037 214644
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 262262 186965 262322 259931
rect 263182 253950 263242 261563
rect 263366 260133 263426 436867
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 270539 396676 270605 396677
rect 270539 396612 270540 396676
rect 270604 396612 270605 396676
rect 270539 396611 270605 396612
rect 269435 387564 269501 387565
rect 269435 387500 269436 387564
rect 269500 387500 269501 387564
rect 269435 387499 269501 387500
rect 266307 379268 266373 379269
rect 266307 379204 266308 379268
rect 266372 379204 266373 379268
rect 266307 379203 266373 379204
rect 265755 378044 265821 378045
rect 265755 377980 265756 378044
rect 265820 377980 265821 378044
rect 265755 377979 265821 377980
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 263547 311268 263613 311269
rect 263547 311204 263548 311268
rect 263612 311204 263613 311268
rect 263547 311203 263613 311204
rect 263550 292501 263610 311203
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 263547 292500 263613 292501
rect 263547 292436 263548 292500
rect 263612 292436 263613 292500
rect 263547 292435 263613 292436
rect 263547 282980 263613 282981
rect 263547 282916 263548 282980
rect 263612 282916 263613 282980
rect 263547 282915 263613 282916
rect 263550 262309 263610 282915
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 263547 262308 263613 262309
rect 263547 262244 263548 262308
rect 263612 262244 263613 262308
rect 263547 262243 263613 262244
rect 263363 260132 263429 260133
rect 263363 260068 263364 260132
rect 263428 260068 263429 260132
rect 263363 260067 263429 260068
rect 263182 253890 263426 253950
rect 263366 244290 263426 253890
rect 263366 244230 263610 244290
rect 263550 228989 263610 244230
rect 264954 230614 265574 266058
rect 265758 262717 265818 377979
rect 265755 262716 265821 262717
rect 265755 262652 265756 262716
rect 265820 262652 265821 262716
rect 265755 262651 265821 262652
rect 265755 260132 265821 260133
rect 265755 260068 265756 260132
rect 265820 260068 265821 260132
rect 265755 260067 265821 260068
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 263547 228988 263613 228989
rect 263547 228924 263548 228988
rect 263612 228924 263613 228988
rect 263547 228923 263613 228924
rect 264954 194614 265574 230058
rect 265758 225589 265818 260067
rect 266310 246261 266370 379203
rect 267779 363628 267845 363629
rect 267779 363564 267780 363628
rect 267844 363564 267845 363628
rect 267779 363563 267845 363564
rect 267782 258229 267842 363563
rect 269251 338740 269317 338741
rect 269251 338676 269252 338740
rect 269316 338676 269317 338740
rect 269251 338675 269317 338676
rect 267963 317660 268029 317661
rect 267963 317596 267964 317660
rect 268028 317596 268029 317660
rect 267963 317595 268029 317596
rect 267779 258228 267845 258229
rect 267779 258164 267780 258228
rect 267844 258164 267845 258228
rect 267779 258163 267845 258164
rect 267779 257412 267845 257413
rect 267779 257348 267780 257412
rect 267844 257348 267845 257412
rect 267779 257347 267845 257348
rect 266491 252652 266557 252653
rect 266491 252588 266492 252652
rect 266556 252588 266557 252652
rect 266491 252587 266557 252588
rect 266307 246260 266373 246261
rect 266307 246196 266308 246260
rect 266372 246196 266373 246260
rect 266307 246195 266373 246196
rect 265755 225588 265821 225589
rect 265755 225524 265756 225588
rect 265820 225524 265821 225588
rect 265755 225523 265821 225524
rect 266494 204917 266554 252587
rect 267782 227629 267842 257347
rect 267966 244221 268026 317595
rect 269254 263397 269314 338675
rect 269251 263396 269317 263397
rect 269251 263332 269252 263396
rect 269316 263332 269317 263396
rect 269251 263331 269317 263332
rect 269067 260812 269133 260813
rect 269067 260748 269068 260812
rect 269132 260748 269133 260812
rect 269067 260747 269133 260748
rect 269070 259453 269130 260747
rect 269067 259452 269133 259453
rect 269067 259388 269068 259452
rect 269132 259388 269133 259452
rect 269067 259387 269133 259388
rect 267963 244220 268029 244221
rect 267963 244156 267964 244220
rect 268028 244156 268029 244220
rect 267963 244155 268029 244156
rect 267779 227628 267845 227629
rect 267779 227564 267780 227628
rect 267844 227564 267845 227628
rect 267779 227563 267845 227564
rect 269070 219333 269130 259387
rect 269438 255237 269498 387499
rect 270542 262853 270602 396611
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 276243 454204 276309 454205
rect 276243 454140 276244 454204
rect 276308 454140 276309 454204
rect 276243 454139 276309 454140
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 274587 380220 274653 380221
rect 274587 380156 274588 380220
rect 274652 380156 274653 380220
rect 274587 380155 274653 380156
rect 273299 369068 273365 369069
rect 273299 369004 273300 369068
rect 273364 369004 273365 369068
rect 273299 369003 273365 369004
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 270539 262852 270605 262853
rect 270539 262788 270540 262852
rect 270604 262788 270605 262852
rect 270539 262787 270605 262788
rect 269435 255236 269501 255237
rect 269435 255172 269436 255236
rect 269500 255172 269501 255236
rect 269435 255171 269501 255172
rect 270539 255236 270605 255237
rect 270539 255172 270540 255236
rect 270604 255172 270605 255236
rect 270539 255171 270605 255172
rect 270542 220149 270602 255171
rect 271794 237454 272414 272898
rect 273302 260813 273362 369003
rect 273299 260812 273365 260813
rect 273299 260748 273300 260812
rect 273364 260748 273365 260812
rect 273299 260747 273365 260748
rect 274590 259453 274650 380155
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 273299 259452 273365 259453
rect 273299 259388 273300 259452
rect 273364 259388 273365 259452
rect 273299 259387 273365 259388
rect 274587 259452 274653 259453
rect 274587 259388 274588 259452
rect 274652 259388 274653 259452
rect 274587 259387 274653 259388
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 270539 220148 270605 220149
rect 270539 220084 270540 220148
rect 270604 220084 270605 220148
rect 270539 220083 270605 220084
rect 269067 219332 269133 219333
rect 269067 219268 269068 219332
rect 269132 219268 269133 219332
rect 269067 219267 269133 219268
rect 269070 218109 269130 219267
rect 269067 218108 269133 218109
rect 269067 218044 269068 218108
rect 269132 218044 269133 218108
rect 269067 218043 269133 218044
rect 266491 204916 266557 204917
rect 266491 204852 266492 204916
rect 266556 204852 266557 204916
rect 266491 204851 266557 204852
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 262259 186964 262325 186965
rect 262259 186900 262260 186964
rect 262324 186900 262325 186964
rect 262259 186899 262325 186900
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 259499 146980 259565 146981
rect 259499 146916 259500 146980
rect 259564 146916 259565 146980
rect 259499 146915 259565 146916
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 201454 272414 236898
rect 273302 214573 273362 259387
rect 275514 241174 276134 276618
rect 276246 245581 276306 454139
rect 279234 424894 279854 460338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 281579 431220 281645 431221
rect 281579 431156 281580 431220
rect 281644 431156 281645 431220
rect 281579 431155 281645 431156
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 277163 359412 277229 359413
rect 277163 359348 277164 359412
rect 277228 359348 277229 359412
rect 277163 359347 277229 359348
rect 276427 255372 276493 255373
rect 276427 255308 276428 255372
rect 276492 255308 276493 255372
rect 276427 255307 276493 255308
rect 276243 245580 276309 245581
rect 276243 245516 276244 245580
rect 276308 245516 276309 245580
rect 276243 245515 276309 245516
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 273299 214572 273365 214573
rect 273299 214508 273300 214572
rect 273364 214508 273365 214572
rect 273299 214507 273365 214508
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 205174 276134 240618
rect 276430 231165 276490 255307
rect 277166 241501 277226 359347
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 280291 311132 280357 311133
rect 280291 311068 280292 311132
rect 280356 311068 280357 311132
rect 280291 311067 280357 311068
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 280294 262173 280354 311067
rect 280291 262172 280357 262173
rect 280291 262108 280292 262172
rect 280356 262108 280357 262172
rect 280291 262107 280357 262108
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 277163 241500 277229 241501
rect 277163 241436 277164 241500
rect 277228 241436 277229 241500
rect 277163 241435 277229 241436
rect 277166 240277 277226 241435
rect 277163 240276 277229 240277
rect 277163 240212 277164 240276
rect 277228 240212 277229 240276
rect 277163 240211 277229 240212
rect 276427 231164 276493 231165
rect 276427 231100 276428 231164
rect 276492 231100 276493 231164
rect 276427 231099 276493 231100
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 208894 279854 244338
rect 281582 242317 281642 431155
rect 282954 428614 283574 464058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 284339 455564 284405 455565
rect 284339 455500 284340 455564
rect 284404 455500 284405 455564
rect 284339 455499 284405 455500
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 284342 264213 284402 455499
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 284339 264212 284405 264213
rect 284339 264148 284340 264212
rect 284404 264148 284405 264212
rect 284339 264147 284405 264148
rect 285627 259588 285693 259589
rect 285627 259524 285628 259588
rect 285692 259524 285693 259588
rect 285627 259523 285693 259524
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 281579 242316 281645 242317
rect 281579 242252 281580 242316
rect 281644 242252 281645 242316
rect 281579 242251 281645 242252
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 285630 148477 285690 259523
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 285627 148476 285693 148477
rect 285627 148412 285628 148476
rect 285692 148412 285693 148476
rect 285627 148411 285693 148412
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 73721 543218 73957 543454
rect 73721 542898 73957 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 77686 561218 77922 561454
rect 77686 560898 77922 561134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 81651 543218 81887 543454
rect 81651 542898 81887 543134
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 85617 561218 85853 561454
rect 85617 560898 85853 561134
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 89582 543218 89818 543454
rect 89582 542898 89818 543134
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 79019 273218 79255 273454
rect 79019 272898 79255 273134
rect 74387 255218 74623 255454
rect 74387 254898 74623 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 83651 255218 83887 255454
rect 83651 254898 83887 255134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 88283 273218 88519 273454
rect 88283 272898 88519 273134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 92915 255218 93151 255454
rect 92915 254898 93151 255134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 77686 129218 77922 129454
rect 77686 128898 77922 129134
rect 85617 129218 85853 129454
rect 85617 128898 85853 129134
rect 73721 111218 73957 111454
rect 73721 110898 73957 111134
rect 81651 111218 81887 111454
rect 81651 110898 81887 111134
rect 89582 111218 89818 111454
rect 89582 110898 89818 111134
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 197818 435218 198054 435454
rect 197818 434898 198054 435134
rect 228538 435218 228774 435454
rect 228538 434898 228774 435134
rect 213178 417218 213414 417454
rect 213178 416898 213414 417134
rect 197818 399218 198054 399454
rect 197818 398898 198054 399134
rect 228538 399218 228774 399454
rect 228538 398898 228774 399134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 243898 417218 244134 417454
rect 243898 416898 244134 417134
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 197818 291218 198054 291454
rect 197818 290898 198054 291134
rect 228538 291218 228774 291454
rect 228538 290898 228774 291134
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 213178 273218 213414 273454
rect 213178 272898 213414 273134
rect 243898 273218 244134 273454
rect 243898 272898 244134 273134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 197818 255218 198054 255454
rect 197818 254898 198054 255134
rect 228538 255218 228774 255454
rect 228538 254898 228774 255134
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 199430 111218 199666 111454
rect 199430 110898 199666 111134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 204306 129218 204542 129454
rect 204306 128898 204542 129134
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 209182 111218 209418 111454
rect 209182 110898 209418 111134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 214058 129218 214294 129454
rect 214058 128898 214294 129134
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 218934 111218 219170 111454
rect 218934 110898 219170 111134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 77686 561454
rect 77922 561218 85617 561454
rect 85853 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 77686 561134
rect 77922 560898 85617 561134
rect 85853 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73721 543454
rect 73957 543218 81651 543454
rect 81887 543218 89582 543454
rect 89818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73721 543134
rect 73957 542898 81651 543134
rect 81887 542898 89582 543134
rect 89818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 197818 435454
rect 198054 435218 228538 435454
rect 228774 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 197818 435134
rect 198054 434898 228538 435134
rect 228774 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 213178 417454
rect 213414 417218 243898 417454
rect 244134 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 213178 417134
rect 213414 416898 243898 417134
rect 244134 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 197818 399454
rect 198054 399218 228538 399454
rect 228774 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 197818 399134
rect 198054 398898 228538 399134
rect 228774 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 197818 291454
rect 198054 291218 228538 291454
rect 228774 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 197818 291134
rect 198054 290898 228538 291134
rect 228774 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 79019 273454
rect 79255 273218 88283 273454
rect 88519 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 213178 273454
rect 213414 273218 243898 273454
rect 244134 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 79019 273134
rect 79255 272898 88283 273134
rect 88519 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 213178 273134
rect 213414 272898 243898 273134
rect 244134 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74387 255454
rect 74623 255218 83651 255454
rect 83887 255218 92915 255454
rect 93151 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 197818 255454
rect 198054 255218 228538 255454
rect 228774 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74387 255134
rect 74623 254898 83651 255134
rect 83887 254898 92915 255134
rect 93151 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 197818 255134
rect 198054 254898 228538 255134
rect 228774 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 77686 129454
rect 77922 129218 85617 129454
rect 85853 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 204306 129454
rect 204542 129218 214058 129454
rect 214294 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 77686 129134
rect 77922 128898 85617 129134
rect 85853 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 204306 129134
rect 204542 128898 214058 129134
rect 214294 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73721 111454
rect 73957 111218 81651 111454
rect 81887 111218 89582 111454
rect 89818 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 199430 111454
rect 199666 111218 209182 111454
rect 209418 111218 218934 111454
rect 219170 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73721 111134
rect 73957 110898 81651 111134
rect 81887 110898 89582 111134
rect 89818 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 199430 111134
rect 199666 110898 209182 111134
rect 209418 110898 218934 111134
rect 219170 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use zube_wrapped_project  zube_wrapped_project_5
timestamp 1635348390
transform 1 0 193568 0 1 241592
box 0 0 60000 60000
use wrapped_ws2812  wrapped_ws2812_4
timestamp 1635348390
transform 1 0 193568 0 1 92782
box 0 0 31475 48253
use wrapped_vga_clock  wrapped_vga_clock_2
timestamp 1635348390
transform 1 0 68770 0 1 390356
box 0 0 44000 44000
use wrapped_tpm2137  wrapped_tpm2137_3
timestamp 1635348390
transform 1 0 68770 0 1 539166
box 0 0 26000 42000
use wrapped_rgb_mixer  wrapped_rgb_mixer_0
timestamp 1635348390
transform 1 0 68770 0 1 92782
box 0 0 26000 42000
use wrapped_hack_soc  wrapped_hack_soc_6
timestamp 1635348390
transform 1 0 193568 0 1 390356
box 0 0 60000 60000
use wrapped_frequency_counter  wrapped_frequency_counter_1
timestamp 1635348390
transform 1 0 68770 0 1 241592
box 0 0 30000 42000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 136782 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 143035 218414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 303592 218414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 303592 254414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 436356 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 583166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 436356 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 452356 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 452356 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 136782 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 143035 222134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 303592 222134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 436356 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 583166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 436356 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 452356 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 136782 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 143035 225854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 303592 225854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 436356 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 583166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 452356 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 136782 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 143035 193574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 303592 193574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 303592 229574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 436356 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 583166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 452356 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 452356 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 90782 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 143035 207854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 303592 207854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 303592 243854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 436356 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 452356 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 452356 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 136782 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 143035 211574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 303592 211574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 303592 247574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 436356 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 583166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 436356 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 452356 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 452356 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 136782 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 143035 200414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 303592 200414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 303592 236414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 436356 92414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 583166 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 452356 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 452356 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 136782 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 143035 204134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 303592 204134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 303592 240134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 436356 96134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 583166 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 452356 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 452356 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
