magic
tech sky130A
magscale 1 2
timestamp 1635173914
<< metal1 >>
rect 70210 703264 70216 703316
rect 70268 703304 70274 703316
rect 154114 703304 154120 703316
rect 70268 703276 154120 703304
rect 70268 703264 70274 703276
rect 154114 703264 154120 703276
rect 154172 703264 154178 703316
rect 89714 703196 89720 703248
rect 89772 703236 89778 703248
rect 235166 703236 235172 703248
rect 89772 703208 235172 703236
rect 89772 703196 89778 703208
rect 235166 703196 235172 703208
rect 235224 703196 235230 703248
rect 119338 703128 119344 703180
rect 119396 703168 119402 703180
rect 218974 703168 218980 703180
rect 119396 703140 218980 703168
rect 119396 703128 119402 703140
rect 218974 703128 218980 703140
rect 219032 703128 219038 703180
rect 271138 703128 271144 703180
rect 271196 703168 271202 703180
rect 397454 703168 397460 703180
rect 271196 703140 397460 703168
rect 271196 703128 271202 703140
rect 397454 703128 397460 703140
rect 397512 703128 397518 703180
rect 67634 703060 67640 703112
rect 67692 703100 67698 703112
rect 170306 703100 170312 703112
rect 67692 703072 170312 703100
rect 67692 703060 67698 703072
rect 170306 703060 170312 703072
rect 170364 703060 170370 703112
rect 276658 703060 276664 703112
rect 276716 703100 276722 703112
rect 413646 703100 413652 703112
rect 276716 703072 413652 703100
rect 276716 703060 276722 703072
rect 413646 703060 413652 703072
rect 413704 703060 413710 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 84102 702992 84108 703044
rect 84160 703032 84166 703044
rect 202782 703032 202788 703044
rect 84160 703004 202788 703032
rect 84160 702992 84166 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 268378 702992 268384 703044
rect 268436 703032 268442 703044
rect 462314 703032 462320 703044
rect 268436 703004 462320 703032
rect 268436 702992 268442 703004
rect 462314 702992 462320 703004
rect 462372 702992 462378 703044
rect 101490 702924 101496 702976
rect 101548 702964 101554 702976
rect 300118 702964 300124 702976
rect 101548 702936 300124 702964
rect 101548 702924 101554 702936
rect 300118 702924 300124 702936
rect 300176 702924 300182 702976
rect 61930 702856 61936 702908
rect 61988 702896 61994 702908
rect 364978 702896 364984 702908
rect 61988 702868 364984 702896
rect 61988 702856 61994 702868
rect 364978 702856 364984 702868
rect 365036 702856 365042 702908
rect 116578 702788 116584 702840
rect 116636 702828 116642 702840
rect 429838 702828 429844 702840
rect 116636 702800 429844 702828
rect 116636 702788 116642 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 24302 702720 24308 702772
rect 24360 702760 24366 702772
rect 86218 702760 86224 702772
rect 24360 702732 86224 702760
rect 24360 702720 24366 702732
rect 86218 702720 86224 702732
rect 86276 702720 86282 702772
rect 99282 702720 99288 702772
rect 99340 702760 99346 702772
rect 478506 702760 478512 702772
rect 99340 702732 478512 702760
rect 99340 702720 99346 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 79962 702652 79968 702704
rect 80020 702692 80026 702704
rect 494790 702692 494796 702704
rect 80020 702664 494796 702692
rect 80020 702652 80026 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 8110 702584 8116 702636
rect 8168 702624 8174 702636
rect 96614 702624 96620 702636
rect 8168 702596 96620 702624
rect 8168 702584 8174 702596
rect 96614 702584 96620 702596
rect 96672 702584 96678 702636
rect 106918 702584 106924 702636
rect 106976 702624 106982 702636
rect 527174 702624 527180 702636
rect 106976 702596 527180 702624
rect 106976 702584 106982 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 57882 702516 57888 702568
rect 57940 702556 57946 702568
rect 582466 702556 582472 702568
rect 57940 702528 582472 702556
rect 57940 702516 57946 702528
rect 582466 702516 582472 702528
rect 582524 702516 582530 702568
rect 66162 702448 66168 702500
rect 66220 702488 66226 702500
rect 559650 702488 559656 702500
rect 66220 702460 559656 702488
rect 66220 702448 66226 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 71682 700272 71688 700324
rect 71740 700312 71746 700324
rect 105446 700312 105452 700324
rect 71740 700284 105452 700312
rect 71740 700272 71746 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 269758 700272 269764 700324
rect 269816 700312 269822 700324
rect 283834 700312 283840 700324
rect 269816 700284 283840 700312
rect 269816 700272 269822 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 286318 700272 286324 700324
rect 286376 700312 286382 700324
rect 332502 700312 332508 700324
rect 286376 700284 332508 700312
rect 286376 700272 286382 700284
rect 332502 700272 332508 700284
rect 332560 700272 332566 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 18598 683176 18604 683188
rect 3476 683148 18604 683176
rect 3476 683136 3482 683148
rect 18598 683136 18604 683148
rect 18656 683136 18662 683188
rect 2774 671032 2780 671084
rect 2832 671072 2838 671084
rect 4798 671072 4804 671084
rect 2832 671044 4804 671072
rect 2832 671032 2838 671044
rect 4798 671032 4804 671044
rect 4856 671032 4862 671084
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 74534 656928 74540 656940
rect 3476 656900 74540 656928
rect 3476 656888 3482 656900
rect 74534 656888 74540 656900
rect 74592 656888 74598 656940
rect 309778 643084 309784 643136
rect 309836 643124 309842 643136
rect 580166 643124 580172 643136
rect 309836 643096 580172 643124
rect 309836 643084 309842 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 39298 618304 39304 618316
rect 3568 618276 39304 618304
rect 3568 618264 3574 618276
rect 39298 618264 39304 618276
rect 39356 618264 39362 618316
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 94774 605860 94780 605872
rect 3568 605832 94780 605860
rect 3568 605820 3574 605832
rect 94774 605820 94780 605832
rect 94832 605820 94838 605872
rect 83458 590656 83464 590708
rect 83516 590696 83522 590708
rect 84102 590696 84108 590708
rect 83516 590668 84108 590696
rect 83516 590656 83522 590668
rect 84102 590656 84108 590668
rect 84160 590696 84166 590708
rect 132586 590696 132592 590708
rect 84160 590668 132592 590696
rect 84160 590656 84166 590668
rect 132586 590656 132592 590668
rect 132644 590656 132650 590708
rect 307018 590656 307024 590708
rect 307076 590696 307082 590708
rect 579798 590696 579804 590708
rect 307076 590668 579804 590696
rect 307076 590656 307082 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 40034 589908 40040 589960
rect 40092 589948 40098 589960
rect 96706 589948 96712 589960
rect 40092 589920 96712 589948
rect 40092 589908 40098 589920
rect 96706 589908 96712 589920
rect 96764 589908 96770 589960
rect 67726 587120 67732 587172
rect 67784 587160 67790 587172
rect 71682 587160 71688 587172
rect 67784 587132 71688 587160
rect 67784 587120 67790 587132
rect 71682 587120 71688 587132
rect 71740 587160 71746 587172
rect 125594 587160 125600 587172
rect 71740 587132 125600 587160
rect 71740 587120 71746 587132
rect 125594 587120 125600 587132
rect 125652 587120 125658 587172
rect 78122 585760 78128 585812
rect 78180 585800 78186 585812
rect 88334 585800 88340 585812
rect 78180 585772 88340 585800
rect 78180 585760 78186 585772
rect 88334 585760 88340 585772
rect 88392 585760 88398 585812
rect 121730 585760 121736 585812
rect 121788 585800 121794 585812
rect 582558 585800 582564 585812
rect 121788 585772 582564 585800
rect 121788 585760 121794 585772
rect 582558 585760 582564 585772
rect 582616 585760 582622 585812
rect 55122 585148 55128 585200
rect 55180 585188 55186 585200
rect 79318 585188 79324 585200
rect 55180 585160 79324 585188
rect 55180 585148 55186 585160
rect 79318 585148 79324 585160
rect 79376 585148 79382 585200
rect 87506 585148 87512 585200
rect 87564 585188 87570 585200
rect 121454 585188 121460 585200
rect 87564 585160 121460 585188
rect 87564 585148 87570 585160
rect 121454 585148 121460 585160
rect 121512 585188 121518 585200
rect 121730 585188 121736 585200
rect 121512 585160 121736 585188
rect 121512 585148 121518 585160
rect 121730 585148 121736 585160
rect 121788 585148 121794 585200
rect 76282 583788 76288 583840
rect 76340 583828 76346 583840
rect 107654 583828 107660 583840
rect 76340 583800 107660 583828
rect 76340 583788 76346 583800
rect 107654 583788 107660 583800
rect 107712 583788 107718 583840
rect 44082 583720 44088 583772
rect 44140 583760 44146 583772
rect 92474 583760 92480 583772
rect 44140 583732 92480 583760
rect 44140 583720 44146 583732
rect 92474 583720 92480 583732
rect 92532 583720 92538 583772
rect 77202 583108 77208 583160
rect 77260 583148 77266 583160
rect 79962 583148 79968 583160
rect 77260 583120 79968 583148
rect 77260 583108 77266 583120
rect 79962 583108 79968 583120
rect 80020 583108 80026 583160
rect 81802 582564 81808 582616
rect 81860 582604 81866 582616
rect 83458 582604 83464 582616
rect 81860 582576 83464 582604
rect 81860 582564 81866 582576
rect 83458 582564 83464 582576
rect 83516 582564 83522 582616
rect 62022 582428 62028 582480
rect 62080 582468 62086 582480
rect 73798 582468 73804 582480
rect 62080 582440 73804 582468
rect 62080 582428 62086 582440
rect 73798 582428 73804 582440
rect 73856 582428 73862 582480
rect 90266 582428 90272 582480
rect 90324 582468 90330 582480
rect 95878 582468 95884 582480
rect 90324 582440 95884 582468
rect 90324 582428 90330 582440
rect 95878 582428 95884 582440
rect 95936 582428 95942 582480
rect 50982 582360 50988 582412
rect 51040 582400 51046 582412
rect 69934 582400 69940 582412
rect 51040 582372 69940 582400
rect 51040 582360 51046 582372
rect 69934 582360 69940 582372
rect 69992 582360 69998 582412
rect 73522 582360 73528 582412
rect 73580 582400 73586 582412
rect 110414 582400 110420 582412
rect 73580 582372 110420 582400
rect 73580 582360 73586 582372
rect 110414 582360 110420 582372
rect 110472 582360 110478 582412
rect 69658 581068 69664 581120
rect 69716 581108 69722 581120
rect 80238 581108 80244 581120
rect 69716 581080 80244 581108
rect 69716 581068 69722 581080
rect 80238 581068 80244 581080
rect 80296 581068 80302 581120
rect 86586 581068 86592 581120
rect 86644 581108 86650 581120
rect 126974 581108 126980 581120
rect 86644 581080 126980 581108
rect 86644 581068 86650 581080
rect 126974 581068 126980 581080
rect 127032 581068 127038 581120
rect 43990 581000 43996 581052
rect 44048 581040 44054 581052
rect 89806 581040 89812 581052
rect 44048 581012 89812 581040
rect 44048 581000 44054 581012
rect 89806 581000 89812 581012
rect 89864 581040 89870 581052
rect 90542 581040 90548 581052
rect 89864 581012 90548 581040
rect 89864 581000 89870 581012
rect 90542 581000 90548 581012
rect 90600 581000 90606 581052
rect 93762 581000 93768 581052
rect 93820 581040 93826 581052
rect 105538 581040 105544 581052
rect 93820 581012 105544 581040
rect 93820 581000 93826 581012
rect 105538 581000 105544 581012
rect 105596 581000 105602 581052
rect 69658 580700 69664 580712
rect 64846 580672 69664 580700
rect 46842 580252 46848 580304
rect 46900 580292 46906 580304
rect 64846 580292 64874 580672
rect 69658 580660 69664 580672
rect 69716 580660 69722 580712
rect 85482 580660 85488 580712
rect 85540 580700 85546 580712
rect 85540 580672 93854 580700
rect 85540 580660 85546 580672
rect 46900 580264 64874 580292
rect 46900 580252 46906 580264
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 46842 579680 46848 579692
rect 3384 579652 46848 579680
rect 3384 579640 3390 579652
rect 46842 579640 46848 579652
rect 46900 579640 46906 579692
rect 64690 579640 64696 579692
rect 64748 579680 64754 579692
rect 66530 579680 66536 579692
rect 64748 579652 66536 579680
rect 64748 579640 64754 579652
rect 66530 579640 66536 579652
rect 66588 579640 66594 579692
rect 93826 579680 93854 580672
rect 113358 579680 113364 579692
rect 93826 579652 113364 579680
rect 113358 579640 113364 579652
rect 113416 579640 113422 579692
rect 94774 579572 94780 579624
rect 94832 579612 94838 579624
rect 96798 579612 96804 579624
rect 94832 579584 96804 579612
rect 94832 579572 94838 579584
rect 96798 579572 96804 579584
rect 96856 579572 96862 579624
rect 97534 576852 97540 576904
rect 97592 576892 97598 576904
rect 118694 576892 118700 576904
rect 97592 576864 118700 576892
rect 97592 576852 97598 576864
rect 118694 576852 118700 576864
rect 118752 576852 118758 576904
rect 97902 576716 97908 576768
rect 97960 576756 97966 576768
rect 99190 576756 99196 576768
rect 97960 576728 99196 576756
rect 97960 576716 97966 576728
rect 99190 576716 99196 576728
rect 99248 576756 99254 576768
rect 101490 576756 101496 576768
rect 99248 576728 101496 576756
rect 99248 576716 99254 576728
rect 101490 576716 101496 576728
rect 101548 576716 101554 576768
rect 3418 576104 3424 576156
rect 3476 576144 3482 576156
rect 33134 576144 33140 576156
rect 3476 576116 33140 576144
rect 3476 576104 3482 576116
rect 33134 576104 33140 576116
rect 33192 576104 33198 576156
rect 33134 575492 33140 575544
rect 33192 575532 33198 575544
rect 34422 575532 34428 575544
rect 33192 575504 34428 575532
rect 33192 575492 33198 575504
rect 34422 575492 34428 575504
rect 34480 575532 34486 575544
rect 66438 575532 66444 575544
rect 34480 575504 66444 575532
rect 34480 575492 34486 575504
rect 66438 575492 66444 575504
rect 66496 575492 66502 575544
rect 97626 575424 97632 575476
rect 97684 575464 97690 575476
rect 106918 575464 106924 575476
rect 97684 575436 106924 575464
rect 97684 575424 97690 575436
rect 106918 575424 106924 575436
rect 106976 575424 106982 575476
rect 97442 572704 97448 572756
rect 97500 572744 97506 572756
rect 100846 572744 100852 572756
rect 97500 572716 100852 572744
rect 97500 572704 97506 572716
rect 100846 572704 100852 572716
rect 100904 572704 100910 572756
rect 99282 571956 99288 572008
rect 99340 571996 99346 572008
rect 106918 571996 106924 572008
rect 99340 571968 106924 571996
rect 99340 571956 99346 571968
rect 106918 571956 106924 571968
rect 106976 571956 106982 572008
rect 64782 571344 64788 571396
rect 64840 571384 64846 571396
rect 66714 571384 66720 571396
rect 64840 571356 66720 571384
rect 64840 571344 64846 571356
rect 66714 571344 66720 571356
rect 66772 571344 66778 571396
rect 97074 571344 97080 571396
rect 97132 571384 97138 571396
rect 100018 571384 100024 571396
rect 97132 571356 100024 571384
rect 97132 571344 97138 571356
rect 100018 571344 100024 571356
rect 100076 571344 100082 571396
rect 56502 570596 56508 570648
rect 56560 570636 56566 570648
rect 66622 570636 66628 570648
rect 56560 570608 66628 570636
rect 56560 570596 56566 570608
rect 66622 570596 66628 570608
rect 66680 570596 66686 570648
rect 97902 570596 97908 570648
rect 97960 570636 97966 570648
rect 103422 570636 103428 570648
rect 97960 570608 103428 570636
rect 97960 570596 97966 570608
rect 103422 570596 103428 570608
rect 103480 570636 103486 570648
rect 582650 570636 582656 570648
rect 103480 570608 582656 570636
rect 103480 570596 103486 570608
rect 582650 570596 582656 570608
rect 582708 570596 582714 570648
rect 103422 569236 103428 569288
rect 103480 569276 103486 569288
rect 114646 569276 114652 569288
rect 103480 569248 114652 569276
rect 103480 569236 103486 569248
rect 114646 569236 114652 569248
rect 114704 569236 114710 569288
rect 97902 569168 97908 569220
rect 97960 569208 97966 569220
rect 133874 569208 133880 569220
rect 97960 569180 133880 569208
rect 97960 569168 97966 569180
rect 133874 569168 133880 569180
rect 133932 569168 133938 569220
rect 95878 567808 95884 567860
rect 95936 567848 95942 567860
rect 103514 567848 103520 567860
rect 95936 567820 103520 567848
rect 95936 567808 95942 567820
rect 103514 567808 103520 567820
rect 103572 567808 103578 567860
rect 49602 565836 49608 565888
rect 49660 565876 49666 565888
rect 67634 565876 67640 565888
rect 49660 565848 67640 565876
rect 49660 565836 49666 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 63402 564408 63408 564460
rect 63460 564448 63466 564460
rect 66806 564448 66812 564460
rect 63460 564420 66812 564448
rect 63460 564408 63466 564420
rect 66806 564408 66812 564420
rect 66864 564408 66870 564460
rect 52362 564340 52368 564392
rect 52420 564380 52426 564392
rect 57882 564380 57888 564392
rect 52420 564352 57888 564380
rect 52420 564340 52426 564352
rect 57882 564340 57888 564352
rect 57940 564380 57946 564392
rect 66530 564380 66536 564392
rect 57940 564352 66536 564380
rect 57940 564340 57946 564352
rect 66530 564340 66536 564352
rect 66588 564340 66594 564392
rect 35802 561688 35808 561740
rect 35860 561728 35866 561740
rect 66806 561728 66812 561740
rect 35860 561700 66812 561728
rect 35860 561688 35866 561700
rect 66806 561688 66812 561700
rect 66864 561688 66870 561740
rect 96798 561688 96804 561740
rect 96856 561728 96862 561740
rect 128354 561728 128360 561740
rect 96856 561700 128360 561728
rect 96856 561688 96862 561700
rect 128354 561688 128360 561700
rect 128412 561688 128418 561740
rect 48222 560260 48228 560312
rect 48280 560300 48286 560312
rect 66806 560300 66812 560312
rect 48280 560272 66812 560300
rect 48280 560260 48286 560272
rect 66806 560260 66812 560272
rect 66864 560260 66870 560312
rect 60642 558900 60648 558952
rect 60700 558940 60706 558952
rect 66806 558940 66812 558952
rect 60700 558912 66812 558940
rect 60700 558900 60706 558912
rect 66806 558900 66812 558912
rect 66864 558900 66870 558952
rect 96798 558900 96804 558952
rect 96856 558940 96862 558952
rect 114554 558940 114560 558952
rect 96856 558912 114560 558940
rect 96856 558900 96862 558912
rect 114554 558900 114560 558912
rect 114612 558900 114618 558952
rect 97166 558696 97172 558748
rect 97224 558736 97230 558748
rect 100754 558736 100760 558748
rect 97224 558708 100760 558736
rect 97224 558696 97230 558708
rect 100754 558696 100760 558708
rect 100812 558696 100818 558748
rect 53650 557540 53656 557592
rect 53708 557580 53714 557592
rect 66806 557580 66812 557592
rect 53708 557552 66812 557580
rect 53708 557540 53714 557552
rect 66806 557540 66812 557552
rect 66864 557540 66870 557592
rect 57882 554752 57888 554804
rect 57940 554792 57946 554804
rect 66714 554792 66720 554804
rect 57940 554764 66720 554792
rect 57940 554752 57946 554764
rect 66714 554752 66720 554764
rect 66772 554752 66778 554804
rect 3510 554004 3516 554056
rect 3568 554044 3574 554056
rect 21358 554044 21364 554056
rect 3568 554016 21364 554044
rect 3568 554004 3574 554016
rect 21358 554004 21364 554016
rect 21416 554004 21422 554056
rect 57238 553392 57244 553444
rect 57296 553432 57302 553444
rect 66806 553432 66812 553444
rect 57296 553404 66812 553432
rect 57296 553392 57302 553404
rect 66806 553392 66812 553404
rect 66864 553392 66870 553444
rect 96982 552032 96988 552084
rect 97040 552072 97046 552084
rect 111794 552072 111800 552084
rect 97040 552044 111800 552072
rect 97040 552032 97046 552044
rect 111794 552032 111800 552044
rect 111852 552032 111858 552084
rect 97902 550604 97908 550656
rect 97960 550644 97966 550656
rect 115934 550644 115940 550656
rect 97960 550616 115940 550644
rect 97960 550604 97966 550616
rect 115934 550604 115940 550616
rect 115992 550604 115998 550656
rect 97074 549312 97080 549364
rect 97132 549352 97138 549364
rect 100110 549352 100116 549364
rect 97132 549324 100116 549352
rect 97132 549312 97138 549324
rect 100110 549312 100116 549324
rect 100168 549312 100174 549364
rect 41322 549244 41328 549296
rect 41380 549284 41386 549296
rect 66806 549284 66812 549296
rect 41380 549256 66812 549284
rect 41380 549244 41386 549256
rect 66806 549244 66812 549256
rect 66864 549244 66870 549296
rect 50890 546456 50896 546508
rect 50948 546496 50954 546508
rect 66530 546496 66536 546508
rect 50948 546468 66536 546496
rect 50948 546456 50954 546468
rect 66530 546456 66536 546468
rect 66588 546456 66594 546508
rect 65978 545096 65984 545148
rect 66036 545136 66042 545148
rect 66162 545136 66168 545148
rect 66036 545108 66168 545136
rect 66036 545096 66042 545108
rect 66162 545096 66168 545108
rect 66220 545096 66226 545148
rect 55030 544348 55036 544400
rect 55088 544388 55094 544400
rect 61930 544388 61936 544400
rect 55088 544360 61936 544388
rect 55088 544348 55094 544360
rect 61930 544348 61936 544360
rect 61988 544388 61994 544400
rect 66346 544388 66352 544400
rect 61988 544360 66352 544388
rect 61988 544348 61994 544360
rect 66346 544348 66352 544360
rect 66404 544348 66410 544400
rect 97350 543736 97356 543788
rect 97408 543776 97414 543788
rect 108298 543776 108304 543788
rect 97408 543748 108304 543776
rect 97408 543736 97414 543748
rect 108298 543736 108304 543748
rect 108356 543736 108362 543788
rect 18598 542988 18604 543040
rect 18656 543028 18662 543040
rect 66162 543028 66168 543040
rect 18656 543000 66168 543028
rect 18656 542988 18662 543000
rect 66162 542988 66168 543000
rect 66220 543028 66226 543040
rect 66622 543028 66628 543040
rect 66220 543000 66628 543028
rect 66220 542988 66226 543000
rect 66622 542988 66628 543000
rect 66680 542988 66686 543040
rect 95142 540880 95148 540932
rect 95200 540920 95206 540932
rect 95510 540920 95516 540932
rect 95200 540892 95516 540920
rect 95200 540880 95206 540892
rect 95510 540880 95516 540892
rect 95568 540880 95574 540932
rect 67450 539860 67456 539912
rect 67508 539900 67514 539912
rect 71774 539900 71780 539912
rect 67508 539872 71780 539900
rect 67508 539860 67514 539872
rect 71774 539860 71780 539872
rect 71832 539860 71838 539912
rect 87598 539792 87604 539844
rect 87656 539832 87662 539844
rect 93854 539832 93860 539844
rect 87656 539804 93860 539832
rect 87656 539792 87662 539804
rect 93854 539792 93860 539804
rect 93912 539792 93918 539844
rect 48130 539588 48136 539640
rect 48188 539628 48194 539640
rect 66622 539628 66628 539640
rect 48188 539600 66628 539628
rect 48188 539588 48194 539600
rect 66622 539588 66628 539600
rect 66680 539588 66686 539640
rect 75178 538840 75184 538892
rect 75236 538880 75242 538892
rect 96890 538880 96896 538892
rect 75236 538852 96896 538880
rect 75236 538840 75242 538852
rect 96890 538840 96896 538852
rect 96948 538840 96954 538892
rect 3418 538228 3424 538280
rect 3476 538268 3482 538280
rect 70946 538268 70952 538280
rect 3476 538240 70952 538268
rect 3476 538228 3482 538240
rect 70946 538228 70952 538240
rect 71004 538228 71010 538280
rect 89714 538228 89720 538280
rect 89772 538268 89778 538280
rect 90174 538268 90180 538280
rect 89772 538240 90180 538268
rect 89772 538228 89778 538240
rect 90174 538228 90180 538240
rect 90232 538268 90238 538280
rect 136634 538268 136640 538280
rect 90232 538240 136640 538268
rect 90232 538228 90238 538240
rect 136634 538228 136640 538240
rect 136692 538228 136698 538280
rect 70946 537548 70952 537600
rect 71004 537588 71010 537600
rect 79318 537588 79324 537600
rect 71004 537560 79324 537588
rect 71004 537548 71010 537560
rect 79318 537548 79324 537560
rect 79376 537548 79382 537600
rect 4798 537480 4804 537532
rect 4856 537520 4862 537532
rect 96614 537520 96620 537532
rect 4856 537492 96620 537520
rect 4856 537480 4862 537492
rect 96614 537480 96620 537492
rect 96672 537480 96678 537532
rect 304258 536800 304264 536852
rect 304316 536840 304322 536852
rect 580166 536840 580172 536852
rect 304316 536812 580172 536840
rect 304316 536800 304322 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 39298 536732 39304 536784
rect 39356 536772 39362 536784
rect 73430 536772 73436 536784
rect 39356 536744 73436 536772
rect 39356 536732 39362 536744
rect 73430 536732 73436 536744
rect 73488 536772 73494 536784
rect 76558 536772 76564 536784
rect 73488 536744 76564 536772
rect 73488 536732 73494 536744
rect 76558 536732 76564 536744
rect 76616 536732 76622 536784
rect 78306 536596 78312 536648
rect 78364 536636 78370 536648
rect 82170 536636 82176 536648
rect 78364 536608 82176 536636
rect 78364 536596 78370 536608
rect 82170 536596 82176 536608
rect 82228 536596 82234 536648
rect 21358 536052 21364 536104
rect 21416 536092 21422 536104
rect 39850 536092 39856 536104
rect 21416 536064 39856 536092
rect 21416 536052 21422 536064
rect 39850 536052 39856 536064
rect 39908 536092 39914 536104
rect 69382 536092 69388 536104
rect 39908 536064 69388 536092
rect 39908 536052 39914 536064
rect 69382 536052 69388 536064
rect 69440 536052 69446 536104
rect 86678 536052 86684 536104
rect 86736 536092 86742 536104
rect 91002 536092 91008 536104
rect 86736 536064 91008 536092
rect 86736 536052 86742 536064
rect 91002 536052 91008 536064
rect 91060 536092 91066 536104
rect 119338 536092 119344 536104
rect 91060 536064 119344 536092
rect 91060 536052 91066 536064
rect 119338 536052 119344 536064
rect 119396 536052 119402 536104
rect 80146 535780 80152 535832
rect 80204 535820 80210 535832
rect 81342 535820 81348 535832
rect 80204 535792 81348 535820
rect 80204 535780 80210 535792
rect 81342 535780 81348 535792
rect 81400 535780 81406 535832
rect 82078 535440 82084 535492
rect 82136 535480 82142 535492
rect 86218 535480 86224 535492
rect 82136 535452 86224 535480
rect 82136 535440 82142 535452
rect 86218 535440 86224 535452
rect 86276 535440 86282 535492
rect 90358 535440 90364 535492
rect 90416 535480 90422 535492
rect 91830 535480 91836 535492
rect 90416 535452 91836 535480
rect 90416 535440 90422 535452
rect 91830 535440 91836 535452
rect 91888 535440 91894 535492
rect 3418 534080 3424 534132
rect 3476 534120 3482 534132
rect 94498 534120 94504 534132
rect 3476 534092 94504 534120
rect 3476 534080 3482 534092
rect 94498 534080 94504 534092
rect 94556 534080 94562 534132
rect 68922 533332 68928 533384
rect 68980 533372 68986 533384
rect 100018 533372 100024 533384
rect 68980 533344 100024 533372
rect 68980 533332 68986 533344
rect 100018 533332 100024 533344
rect 100076 533332 100082 533384
rect 82078 530612 82084 530664
rect 82136 530652 82142 530664
rect 91186 530652 91192 530664
rect 82136 530624 91192 530652
rect 82136 530612 82142 530624
rect 91186 530612 91192 530624
rect 91244 530612 91250 530664
rect 61930 530544 61936 530596
rect 61988 530584 61994 530596
rect 96798 530584 96804 530596
rect 61988 530556 96804 530584
rect 61988 530544 61994 530556
rect 96798 530544 96804 530556
rect 96856 530544 96862 530596
rect 88334 530136 88340 530188
rect 88392 530176 88398 530188
rect 88886 530176 88892 530188
rect 88392 530148 88892 530176
rect 88392 530136 88398 530148
rect 88886 530136 88892 530148
rect 88944 530136 88950 530188
rect 3510 527824 3516 527876
rect 3568 527864 3574 527876
rect 118694 527864 118700 527876
rect 3568 527836 118700 527864
rect 3568 527824 3574 527836
rect 118694 527824 118700 527836
rect 118752 527824 118758 527876
rect 83458 525036 83464 525088
rect 83516 525076 83522 525088
rect 100846 525076 100852 525088
rect 83516 525048 100852 525076
rect 83516 525036 83522 525048
rect 100846 525036 100852 525048
rect 100904 525036 100910 525088
rect 88242 522248 88248 522300
rect 88300 522288 88306 522300
rect 97994 522288 98000 522300
rect 88300 522260 98000 522288
rect 88300 522248 88306 522260
rect 97994 522248 98000 522260
rect 98052 522248 98058 522300
rect 76558 519528 76564 519580
rect 76616 519568 76622 519580
rect 102226 519568 102232 519580
rect 76616 519540 102232 519568
rect 76616 519528 76622 519540
rect 102226 519528 102232 519540
rect 102284 519528 102290 519580
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 11698 514808 11704 514820
rect 3568 514780 11704 514808
rect 3568 514768 3574 514780
rect 11698 514768 11704 514780
rect 11756 514768 11762 514820
rect 48222 511232 48228 511284
rect 48280 511272 48286 511284
rect 580166 511272 580172 511284
rect 48280 511244 580172 511272
rect 48280 511232 48286 511244
rect 580166 511232 580172 511244
rect 580224 511232 580230 511284
rect 82906 487772 82912 487824
rect 82964 487812 82970 487824
rect 111058 487812 111064 487824
rect 82964 487784 111064 487812
rect 82964 487772 82970 487784
rect 111058 487772 111064 487784
rect 111116 487772 111122 487824
rect 65978 485052 65984 485104
rect 66036 485092 66042 485104
rect 118786 485092 118792 485104
rect 66036 485064 118792 485092
rect 66036 485052 66042 485064
rect 118786 485052 118792 485064
rect 118844 485052 118850 485104
rect 82170 482264 82176 482316
rect 82228 482304 82234 482316
rect 109678 482304 109684 482316
rect 82228 482276 109684 482304
rect 82228 482264 82234 482276
rect 109678 482264 109684 482276
rect 109736 482264 109742 482316
rect 64690 479476 64696 479528
rect 64748 479516 64754 479528
rect 92566 479516 92572 479528
rect 64748 479488 92572 479516
rect 64748 479476 64754 479488
rect 92566 479476 92572 479488
rect 92624 479476 92630 479528
rect 86862 478116 86868 478168
rect 86920 478156 86926 478168
rect 95326 478156 95332 478168
rect 86920 478128 95332 478156
rect 86920 478116 86926 478128
rect 95326 478116 95332 478128
rect 95384 478116 95390 478168
rect 64690 476756 64696 476808
rect 64748 476796 64754 476808
rect 84194 476796 84200 476808
rect 64748 476768 84200 476796
rect 64748 476756 64754 476768
rect 84194 476756 84200 476768
rect 84252 476756 84258 476808
rect 2958 475668 2964 475720
rect 3016 475708 3022 475720
rect 4062 475708 4068 475720
rect 3016 475680 4068 475708
rect 3016 475668 3022 475680
rect 4062 475668 4068 475680
rect 4120 475708 4126 475720
rect 4798 475708 4804 475720
rect 4120 475680 4804 475708
rect 4120 475668 4126 475680
rect 4798 475668 4804 475680
rect 4856 475668 4862 475720
rect 66070 475328 66076 475380
rect 66128 475368 66134 475380
rect 98638 475368 98644 475380
rect 66128 475340 98644 475368
rect 66128 475328 66134 475340
rect 98638 475328 98644 475340
rect 98696 475328 98702 475380
rect 65978 474036 65984 474088
rect 66036 474076 66042 474088
rect 75914 474076 75920 474088
rect 66036 474048 75920 474076
rect 66036 474036 66042 474048
rect 75914 474036 75920 474048
rect 75972 474036 75978 474088
rect 67726 473968 67732 474020
rect 67784 474008 67790 474020
rect 120166 474008 120172 474020
rect 67784 473980 120172 474008
rect 67784 473968 67790 473980
rect 120166 473968 120172 473980
rect 120224 473968 120230 474020
rect 74442 471248 74448 471300
rect 74500 471288 74506 471300
rect 112714 471288 112720 471300
rect 74500 471260 112720 471288
rect 74500 471248 74506 471260
rect 112714 471248 112720 471260
rect 112772 471248 112778 471300
rect 67726 469820 67732 469872
rect 67784 469860 67790 469872
rect 96706 469860 96712 469872
rect 67784 469832 96712 469860
rect 67784 469820 67790 469832
rect 96706 469820 96712 469832
rect 96764 469820 96770 469872
rect 85574 468460 85580 468512
rect 85632 468500 85638 468512
rect 116118 468500 116124 468512
rect 85632 468472 116124 468500
rect 85632 468460 85638 468472
rect 116118 468460 116124 468472
rect 116176 468460 116182 468512
rect 77110 467100 77116 467152
rect 77168 467140 77174 467152
rect 89714 467140 89720 467152
rect 77168 467112 89720 467140
rect 77168 467100 77174 467112
rect 89714 467100 89720 467112
rect 89772 467100 89778 467152
rect 78674 465672 78680 465724
rect 78732 465712 78738 465724
rect 100110 465712 100116 465724
rect 78732 465684 100116 465712
rect 78732 465672 78738 465684
rect 100110 465672 100116 465684
rect 100168 465672 100174 465724
rect 67818 464312 67824 464364
rect 67876 464352 67882 464364
rect 118970 464352 118976 464364
rect 67876 464324 118976 464352
rect 67876 464312 67882 464324
rect 118970 464312 118976 464324
rect 119028 464312 119034 464364
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 29638 462380 29644 462392
rect 3292 462352 29644 462380
rect 3292 462340 3298 462352
rect 29638 462340 29644 462352
rect 29696 462340 29702 462392
rect 92474 461592 92480 461644
rect 92532 461632 92538 461644
rect 125870 461632 125876 461644
rect 92532 461604 125876 461632
rect 92532 461592 92538 461604
rect 125870 461592 125876 461604
rect 125928 461592 125934 461644
rect 77202 459688 77208 459740
rect 77260 459728 77266 459740
rect 77938 459728 77944 459740
rect 77260 459700 77944 459728
rect 77260 459688 77266 459700
rect 77938 459688 77944 459700
rect 77996 459688 78002 459740
rect 64782 458804 64788 458856
rect 64840 458844 64846 458856
rect 107010 458844 107016 458856
rect 64840 458816 107016 458844
rect 64840 458804 64846 458816
rect 107010 458804 107016 458816
rect 107068 458804 107074 458856
rect 79318 457444 79324 457496
rect 79376 457484 79382 457496
rect 121638 457484 121644 457496
rect 79376 457456 121644 457484
rect 79376 457444 79382 457456
rect 121638 457444 121644 457456
rect 121696 457444 121702 457496
rect 64782 456016 64788 456068
rect 64840 456056 64846 456068
rect 86954 456056 86960 456068
rect 64840 456028 86960 456056
rect 64840 456016 64846 456028
rect 86954 456016 86960 456028
rect 87012 456016 87018 456068
rect 99190 456016 99196 456068
rect 99248 456056 99254 456068
rect 117406 456056 117412 456068
rect 99248 456028 117412 456056
rect 99248 456016 99254 456028
rect 117406 456016 117412 456028
rect 117464 456016 117470 456068
rect 94498 452548 94504 452600
rect 94556 452588 94562 452600
rect 96706 452588 96712 452600
rect 94556 452560 96712 452588
rect 94556 452548 94562 452560
rect 96706 452548 96712 452560
rect 96764 452548 96770 452600
rect 68462 451868 68468 451920
rect 68520 451908 68526 451920
rect 90358 451908 90364 451920
rect 68520 451880 90364 451908
rect 68520 451868 68526 451880
rect 90358 451868 90364 451880
rect 90416 451868 90422 451920
rect 71866 450508 71872 450560
rect 71924 450548 71930 450560
rect 120350 450548 120356 450560
rect 71924 450520 120356 450548
rect 71924 450508 71930 450520
rect 120350 450508 120356 450520
rect 120408 450508 120414 450560
rect 53650 449148 53656 449200
rect 53708 449188 53714 449200
rect 85666 449188 85672 449200
rect 53708 449160 85672 449188
rect 53708 449148 53714 449160
rect 85666 449148 85672 449160
rect 85724 449148 85730 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 21358 448576 21364 448588
rect 3200 448548 21364 448576
rect 3200 448536 3206 448548
rect 21358 448536 21364 448548
rect 21416 448536 21422 448588
rect 11698 448468 11704 448520
rect 11756 448508 11762 448520
rect 103514 448508 103520 448520
rect 11756 448480 103520 448508
rect 11756 448468 11762 448480
rect 103514 448468 103520 448480
rect 103572 448508 103578 448520
rect 103698 448508 103704 448520
rect 103572 448480 103704 448508
rect 103572 448468 103578 448480
rect 103698 448468 103704 448480
rect 103756 448468 103762 448520
rect 66162 446360 66168 446412
rect 66220 446400 66226 446412
rect 80330 446400 80336 446412
rect 66220 446372 80336 446400
rect 66220 446360 66226 446372
rect 80330 446360 80336 446372
rect 80388 446360 80394 446412
rect 67634 445136 67640 445188
rect 67692 445176 67698 445188
rect 83090 445176 83096 445188
rect 67692 445148 83096 445176
rect 67692 445136 67698 445148
rect 83090 445136 83096 445148
rect 83148 445136 83154 445188
rect 82814 445000 82820 445052
rect 82872 445040 82878 445052
rect 109034 445040 109040 445052
rect 82872 445012 109040 445040
rect 82872 445000 82878 445012
rect 109034 445000 109040 445012
rect 109092 445000 109098 445052
rect 65886 444728 65892 444780
rect 65944 444768 65950 444780
rect 70486 444768 70492 444780
rect 65944 444740 70492 444768
rect 65944 444728 65950 444740
rect 70486 444728 70492 444740
rect 70544 444728 70550 444780
rect 81618 443640 81624 443692
rect 81676 443680 81682 443692
rect 100754 443680 100760 443692
rect 81676 443652 100760 443680
rect 81676 443640 81682 443652
rect 100754 443640 100760 443652
rect 100812 443640 100818 443692
rect 50982 442212 50988 442264
rect 51040 442252 51046 442264
rect 95234 442252 95240 442264
rect 51040 442224 95240 442252
rect 51040 442212 51046 442224
rect 95234 442212 95240 442224
rect 95292 442212 95298 442264
rect 102134 442008 102140 442060
rect 102192 442048 102198 442060
rect 102778 442048 102784 442060
rect 102192 442020 102784 442048
rect 102192 442008 102198 442020
rect 102778 442008 102784 442020
rect 102836 442008 102842 442060
rect 102778 441600 102784 441652
rect 102836 441640 102842 441652
rect 128446 441640 128452 441652
rect 102836 441612 128452 441640
rect 102836 441600 102842 441612
rect 128446 441600 128452 441612
rect 128504 441600 128510 441652
rect 52362 440852 52368 440904
rect 52420 440892 52426 440904
rect 88702 440892 88708 440904
rect 52420 440864 88708 440892
rect 52420 440852 52426 440864
rect 88702 440852 88708 440864
rect 88760 440852 88766 440904
rect 108114 440308 108120 440360
rect 108172 440348 108178 440360
rect 136726 440348 136732 440360
rect 108172 440320 136732 440348
rect 108172 440308 108178 440320
rect 136726 440308 136732 440320
rect 136784 440308 136790 440360
rect 46750 440240 46756 440292
rect 46808 440280 46814 440292
rect 52362 440280 52368 440292
rect 46808 440252 52368 440280
rect 46808 440240 46814 440252
rect 52362 440240 52368 440252
rect 52420 440240 52426 440292
rect 94130 440240 94136 440292
rect 94188 440280 94194 440292
rect 95142 440280 95148 440292
rect 94188 440252 95148 440280
rect 94188 440240 94194 440252
rect 95142 440240 95148 440252
rect 95200 440280 95206 440292
rect 125778 440280 125784 440292
rect 95200 440252 125784 440280
rect 95200 440240 95206 440252
rect 125778 440240 125784 440252
rect 125836 440240 125842 440292
rect 48222 439492 48228 439544
rect 48280 439532 48286 439544
rect 74718 439532 74724 439544
rect 48280 439504 74724 439532
rect 48280 439492 48286 439504
rect 74718 439492 74724 439504
rect 74776 439492 74782 439544
rect 105538 439492 105544 439544
rect 105596 439532 105602 439544
rect 116210 439532 116216 439544
rect 105596 439504 116216 439532
rect 105596 439492 105602 439504
rect 116210 439492 116216 439504
rect 116268 439492 116274 439544
rect 90082 438880 90088 438932
rect 90140 438920 90146 438932
rect 122926 438920 122932 438932
rect 90140 438892 122932 438920
rect 90140 438880 90146 438892
rect 122926 438880 122932 438892
rect 122984 438880 122990 438932
rect 55030 438132 55036 438184
rect 55088 438172 55094 438184
rect 83734 438172 83740 438184
rect 55088 438144 83740 438172
rect 55088 438132 55094 438144
rect 83734 438132 83740 438144
rect 83792 438132 83798 438184
rect 91002 438132 91008 438184
rect 91060 438172 91066 438184
rect 106090 438172 106096 438184
rect 91060 438144 106096 438172
rect 91060 438132 91066 438144
rect 106090 438132 106096 438144
rect 106148 438132 106154 438184
rect 106642 437520 106648 437572
rect 106700 437560 106706 437572
rect 118878 437560 118884 437572
rect 106700 437532 118884 437560
rect 106700 437520 106706 437532
rect 118878 437520 118884 437532
rect 118936 437520 118942 437572
rect 106090 437452 106096 437504
rect 106148 437492 106154 437504
rect 123018 437492 123024 437504
rect 106148 437464 123024 437492
rect 106148 437452 106154 437464
rect 123018 437452 123024 437464
rect 123076 437452 123082 437504
rect 71130 437384 71136 437436
rect 71188 437424 71194 437436
rect 75178 437424 75184 437436
rect 71188 437396 75184 437424
rect 71188 437384 71194 437396
rect 75178 437384 75184 437396
rect 75236 437384 75242 437436
rect 90450 437384 90456 437436
rect 90508 437424 90514 437436
rect 94222 437424 94228 437436
rect 90508 437396 94228 437424
rect 90508 437384 90514 437396
rect 94222 437384 94228 437396
rect 94280 437384 94286 437436
rect 100110 437384 100116 437436
rect 100168 437424 100174 437436
rect 104618 437424 104624 437436
rect 100168 437396 104624 437424
rect 100168 437384 100174 437396
rect 104618 437384 104624 437396
rect 104676 437384 104682 437436
rect 95234 437112 95240 437164
rect 95292 437152 95298 437164
rect 95878 437152 95884 437164
rect 95292 437124 95884 437152
rect 95292 437112 95298 437124
rect 95878 437112 95884 437124
rect 95936 437112 95942 437164
rect 67082 436704 67088 436756
rect 67140 436744 67146 436756
rect 74626 436744 74632 436756
rect 67140 436716 74632 436744
rect 67140 436704 67146 436716
rect 74626 436704 74632 436716
rect 74684 436704 74690 436756
rect 116026 436704 116032 436756
rect 116084 436744 116090 436756
rect 582374 436744 582380 436756
rect 116084 436716 582380 436744
rect 116084 436704 116090 436716
rect 582374 436704 582380 436716
rect 582432 436704 582438 436756
rect 85114 436568 85120 436620
rect 85172 436608 85178 436620
rect 87598 436608 87604 436620
rect 85172 436580 87604 436608
rect 85172 436568 85178 436580
rect 87598 436568 87604 436580
rect 87656 436568 87662 436620
rect 77386 436432 77392 436484
rect 77444 436472 77450 436484
rect 82078 436472 82084 436484
rect 77444 436444 82084 436472
rect 77444 436432 77450 436444
rect 82078 436432 82084 436444
rect 82136 436432 82142 436484
rect 103790 436160 103796 436212
rect 103848 436200 103854 436212
rect 104618 436200 104624 436212
rect 103848 436172 104624 436200
rect 103848 436160 103854 436172
rect 104618 436160 104624 436172
rect 104676 436200 104682 436212
rect 123478 436200 123484 436212
rect 104676 436172 123484 436200
rect 104676 436160 104682 436172
rect 123478 436160 123484 436172
rect 123536 436160 123542 436212
rect 18598 436092 18604 436144
rect 18656 436132 18662 436144
rect 71130 436132 71136 436144
rect 18656 436104 71136 436132
rect 18656 436092 18662 436104
rect 71130 436092 71136 436104
rect 71188 436092 71194 436144
rect 95878 436092 95884 436144
rect 95936 436132 95942 436144
rect 116026 436132 116032 436144
rect 95936 436104 116032 436132
rect 95936 436092 95942 436104
rect 116026 436092 116032 436104
rect 116084 436092 116090 436144
rect 69106 435208 69112 435260
rect 69164 435248 69170 435260
rect 69934 435248 69940 435260
rect 69164 435220 69940 435248
rect 69164 435208 69170 435220
rect 69934 435208 69940 435220
rect 69992 435208 69998 435260
rect 50982 434800 50988 434852
rect 51040 434840 51046 434852
rect 69106 434840 69112 434852
rect 51040 434812 69112 434840
rect 51040 434800 51046 434812
rect 69106 434800 69112 434812
rect 69164 434800 69170 434852
rect 111794 434840 111800 434852
rect 109006 434812 111800 434840
rect 4798 434732 4804 434784
rect 4856 434772 4862 434784
rect 109006 434772 109034 434812
rect 111794 434800 111800 434812
rect 111852 434840 111858 434852
rect 112622 434840 112628 434852
rect 111852 434812 112628 434840
rect 111852 434800 111858 434812
rect 112622 434800 112628 434812
rect 112680 434840 112686 434852
rect 112680 434812 118694 434840
rect 112680 434800 112686 434812
rect 4856 434744 109034 434772
rect 4856 434732 4862 434744
rect 109678 434732 109684 434784
rect 109736 434772 109742 434784
rect 114094 434772 114100 434784
rect 109736 434744 114100 434772
rect 109736 434732 109742 434744
rect 114094 434732 114100 434744
rect 114152 434732 114158 434784
rect 118666 434772 118694 434812
rect 134518 434772 134524 434784
rect 118666 434744 134524 434772
rect 134518 434732 134524 434744
rect 134576 434732 134582 434784
rect 71774 434528 71780 434580
rect 71832 434568 71838 434580
rect 73016 434568 73022 434580
rect 71832 434540 73022 434568
rect 71832 434528 71838 434540
rect 73016 434528 73022 434540
rect 73074 434528 73080 434580
rect 68646 434188 68652 434240
rect 68704 434228 68710 434240
rect 71774 434228 71780 434240
rect 68704 434200 71780 434228
rect 68704 434188 68710 434200
rect 71774 434188 71780 434200
rect 71832 434188 71838 434240
rect 53742 433984 53748 434036
rect 53800 434024 53806 434036
rect 63218 434024 63224 434036
rect 53800 433996 63224 434024
rect 53800 433984 53806 433996
rect 63218 433984 63224 433996
rect 63276 434024 63282 434036
rect 66346 434024 66352 434036
rect 63276 433996 66352 434024
rect 63276 433984 63282 433996
rect 66346 433984 66352 433996
rect 66404 433984 66410 434036
rect 72602 433780 72608 433832
rect 72660 433820 72666 433832
rect 72660 433792 74534 433820
rect 72660 433780 72666 433792
rect 73982 433712 73988 433764
rect 74040 433712 74046 433764
rect 68278 433644 68284 433696
rect 68336 433684 68342 433696
rect 69198 433684 69204 433696
rect 68336 433656 69204 433684
rect 68336 433644 68342 433656
rect 69198 433644 69204 433656
rect 69256 433644 69262 433696
rect 70854 433644 70860 433696
rect 70912 433644 70918 433696
rect 67450 433236 67456 433288
rect 67508 433276 67514 433288
rect 70872 433276 70900 433644
rect 67508 433248 70900 433276
rect 67508 433236 67514 433248
rect 39942 432556 39948 432608
rect 40000 432596 40006 432608
rect 74000 432596 74028 433712
rect 74506 433344 74534 433792
rect 111058 433780 111064 433832
rect 111116 433820 111122 433832
rect 113174 433820 113180 433832
rect 111116 433792 113180 433820
rect 111116 433780 111122 433792
rect 113174 433780 113180 433792
rect 113232 433780 113238 433832
rect 111610 433644 111616 433696
rect 111668 433684 111674 433696
rect 112806 433684 112812 433696
rect 111668 433656 112812 433684
rect 111668 433644 111674 433656
rect 112806 433644 112812 433656
rect 112864 433644 112870 433696
rect 106246 433384 115934 433412
rect 106246 433344 106274 433384
rect 74506 433316 106274 433344
rect 115906 433344 115934 433384
rect 132494 433344 132500 433356
rect 115906 433316 132500 433344
rect 132494 433304 132500 433316
rect 132552 433304 132558 433356
rect 112806 433236 112812 433288
rect 112864 433276 112870 433288
rect 120258 433276 120264 433288
rect 112864 433248 120264 433276
rect 112864 433236 112870 433248
rect 120258 433236 120264 433248
rect 120316 433236 120322 433288
rect 40000 432568 74028 432596
rect 40000 432556 40006 432568
rect 57514 431944 57520 431996
rect 57572 431984 57578 431996
rect 66806 431984 66812 431996
rect 57572 431956 66812 431984
rect 57572 431944 57578 431956
rect 66806 431944 66812 431956
rect 66864 431944 66870 431996
rect 114738 431944 114744 431996
rect 114796 431984 114802 431996
rect 124214 431984 124220 431996
rect 114796 431956 124220 431984
rect 114796 431944 114802 431956
rect 124214 431944 124220 431956
rect 124272 431944 124278 431996
rect 58894 430584 58900 430636
rect 58952 430624 58958 430636
rect 66806 430624 66812 430636
rect 58952 430596 66812 430624
rect 58952 430584 58958 430596
rect 66806 430584 66812 430596
rect 66864 430584 66870 430636
rect 114738 430584 114744 430636
rect 114796 430624 114802 430636
rect 135254 430624 135260 430636
rect 114796 430596 135260 430624
rect 114796 430584 114802 430596
rect 135254 430584 135260 430596
rect 135312 430584 135318 430636
rect 60550 429224 60556 429276
rect 60608 429264 60614 429276
rect 66254 429264 66260 429276
rect 60608 429236 66260 429264
rect 60608 429224 60614 429236
rect 66254 429224 66260 429236
rect 66312 429224 66318 429276
rect 53650 429156 53656 429208
rect 53708 429196 53714 429208
rect 66806 429196 66812 429208
rect 53708 429168 66812 429196
rect 53708 429156 53714 429168
rect 66806 429156 66812 429168
rect 66864 429156 66870 429208
rect 115382 427796 115388 427848
rect 115440 427836 115446 427848
rect 118786 427836 118792 427848
rect 115440 427808 118792 427836
rect 115440 427796 115446 427808
rect 118786 427796 118792 427808
rect 118844 427836 118850 427848
rect 121546 427836 121552 427848
rect 118844 427808 121552 427836
rect 118844 427796 118850 427808
rect 121546 427796 121552 427808
rect 121604 427796 121610 427848
rect 56410 426436 56416 426488
rect 56468 426476 56474 426488
rect 66806 426476 66812 426488
rect 56468 426448 66812 426476
rect 56468 426436 56474 426448
rect 66806 426436 66812 426448
rect 66864 426436 66870 426488
rect 114094 426436 114100 426488
rect 114152 426476 114158 426488
rect 141418 426476 141424 426488
rect 114152 426448 141424 426476
rect 114152 426436 114158 426448
rect 141418 426436 141424 426448
rect 141476 426436 141482 426488
rect 118786 426368 118792 426420
rect 118844 426408 118850 426420
rect 122834 426408 122840 426420
rect 118844 426380 122840 426408
rect 118844 426368 118850 426380
rect 122834 426368 122840 426380
rect 122892 426368 122898 426420
rect 45462 425688 45468 425740
rect 45520 425728 45526 425740
rect 65886 425728 65892 425740
rect 45520 425700 65892 425728
rect 45520 425688 45526 425700
rect 65886 425688 65892 425700
rect 65944 425728 65950 425740
rect 66530 425728 66536 425740
rect 65944 425700 66536 425728
rect 65944 425688 65950 425700
rect 66530 425688 66536 425700
rect 66588 425688 66594 425740
rect 115842 425076 115848 425128
rect 115900 425116 115906 425128
rect 118786 425116 118792 425128
rect 115900 425088 118792 425116
rect 115900 425076 115906 425088
rect 118786 425076 118792 425088
rect 118844 425076 118850 425128
rect 115842 424328 115848 424380
rect 115900 424368 115906 424380
rect 142154 424368 142160 424380
rect 115900 424340 142160 424368
rect 115900 424328 115906 424340
rect 142154 424328 142160 424340
rect 142212 424328 142218 424380
rect 52362 423648 52368 423700
rect 52420 423688 52426 423700
rect 66622 423688 66628 423700
rect 52420 423660 66628 423688
rect 52420 423648 52426 423660
rect 66622 423648 66628 423660
rect 66680 423648 66686 423700
rect 2774 423580 2780 423632
rect 2832 423620 2838 423632
rect 4798 423620 4804 423632
rect 2832 423592 4804 423620
rect 2832 423580 2838 423592
rect 4798 423580 4804 423592
rect 4856 423580 4862 423632
rect 60734 423444 60740 423496
rect 60792 423484 60798 423496
rect 61930 423484 61936 423496
rect 60792 423456 61936 423484
rect 60792 423444 60798 423456
rect 61930 423444 61936 423456
rect 61988 423484 61994 423496
rect 66806 423484 66812 423496
rect 61988 423456 66812 423484
rect 61988 423444 61994 423456
rect 66806 423444 66812 423456
rect 66864 423444 66870 423496
rect 37182 422900 37188 422952
rect 37240 422940 37246 422952
rect 60734 422940 60740 422952
rect 37240 422912 60740 422940
rect 37240 422900 37246 422912
rect 60734 422900 60740 422912
rect 60792 422900 60798 422952
rect 115842 422900 115848 422952
rect 115900 422940 115906 422952
rect 121638 422940 121644 422952
rect 115900 422912 121644 422940
rect 115900 422900 115906 422912
rect 121638 422900 121644 422912
rect 121696 422940 121702 422952
rect 144178 422940 144184 422952
rect 121696 422912 144184 422940
rect 121696 422900 121702 422912
rect 144178 422900 144184 422912
rect 144236 422900 144242 422952
rect 115842 421948 115848 422000
rect 115900 421988 115906 422000
rect 118970 421988 118976 422000
rect 115900 421960 118976 421988
rect 115900 421948 115906 421960
rect 118970 421948 118976 421960
rect 119028 421948 119034 422000
rect 118970 421540 118976 421592
rect 119028 421580 119034 421592
rect 151078 421580 151084 421592
rect 119028 421552 151084 421580
rect 119028 421540 119034 421552
rect 151078 421540 151084 421552
rect 151136 421540 151142 421592
rect 43990 420928 43996 420980
rect 44048 420968 44054 420980
rect 48222 420968 48228 420980
rect 44048 420940 48228 420968
rect 44048 420928 44054 420940
rect 48222 420928 48228 420940
rect 48280 420968 48286 420980
rect 66806 420968 66812 420980
rect 48280 420940 66812 420968
rect 48280 420928 48286 420940
rect 66806 420928 66812 420940
rect 66864 420928 66870 420980
rect 66990 419568 66996 419620
rect 67048 419568 67054 419620
rect 60458 419500 60464 419552
rect 60516 419540 60522 419552
rect 66806 419540 66812 419552
rect 60516 419512 66812 419540
rect 60516 419500 60522 419512
rect 66806 419500 66812 419512
rect 66864 419500 66870 419552
rect 66806 419364 66812 419416
rect 66864 419404 66870 419416
rect 67008 419404 67036 419568
rect 66864 419376 67036 419404
rect 66864 419364 66870 419376
rect 66806 418248 66812 418260
rect 45526 418220 66812 418248
rect 43898 418140 43904 418192
rect 43956 418180 43962 418192
rect 45526 418180 45554 418220
rect 66806 418208 66812 418220
rect 66864 418208 66870 418260
rect 43956 418152 45554 418180
rect 43956 418140 43962 418152
rect 64138 418140 64144 418192
rect 64196 418180 64202 418192
rect 66990 418180 66996 418192
rect 64196 418152 66996 418180
rect 64196 418140 64202 418152
rect 66990 418140 66996 418152
rect 67048 418140 67054 418192
rect 34238 416780 34244 416832
rect 34296 416820 34302 416832
rect 57238 416820 57244 416832
rect 34296 416792 57244 416820
rect 34296 416780 34302 416792
rect 57238 416780 57244 416792
rect 57296 416820 57302 416832
rect 57296 416792 57928 416820
rect 57296 416780 57302 416792
rect 57900 416752 57928 416792
rect 115842 416780 115848 416832
rect 115900 416820 115906 416832
rect 121638 416820 121644 416832
rect 115900 416792 121644 416820
rect 115900 416780 115906 416792
rect 121638 416780 121644 416792
rect 121696 416780 121702 416832
rect 66714 416752 66720 416764
rect 57900 416724 66720 416752
rect 66714 416712 66720 416724
rect 66772 416712 66778 416764
rect 115198 415692 115204 415744
rect 115256 415732 115262 415744
rect 116210 415732 116216 415744
rect 115256 415704 116216 415732
rect 115256 415692 115262 415704
rect 116210 415692 116216 415704
rect 116268 415692 116274 415744
rect 119338 415352 119344 415404
rect 119396 415392 119402 415404
rect 120166 415392 120172 415404
rect 119396 415364 120172 415392
rect 119396 415352 119402 415364
rect 120166 415352 120172 415364
rect 120224 415352 120230 415404
rect 115842 414876 115848 414928
rect 115900 414916 115906 414928
rect 119338 414916 119344 414928
rect 115900 414888 119344 414916
rect 115900 414876 115906 414888
rect 119338 414876 119344 414888
rect 119396 414876 119402 414928
rect 54846 414060 54852 414112
rect 54904 414100 54910 414112
rect 66714 414100 66720 414112
rect 54904 414072 66720 414100
rect 54904 414060 54910 414072
rect 66714 414060 66720 414072
rect 66772 414060 66778 414112
rect 49510 413992 49516 414044
rect 49568 414032 49574 414044
rect 67726 414032 67732 414044
rect 49568 414004 67732 414032
rect 49568 413992 49574 414004
rect 67726 413992 67732 414004
rect 67784 413992 67790 414044
rect 115198 413992 115204 414044
rect 115256 414032 115262 414044
rect 143534 414032 143540 414044
rect 115256 414004 143540 414032
rect 115256 413992 115262 414004
rect 143534 413992 143540 414004
rect 143592 413992 143598 414044
rect 115842 413924 115848 413976
rect 115900 413964 115906 413976
rect 128354 413964 128360 413976
rect 115900 413936 128360 413964
rect 115900 413924 115906 413936
rect 128354 413924 128360 413936
rect 128412 413924 128418 413976
rect 33042 413244 33048 413296
rect 33100 413284 33106 413296
rect 59262 413284 59268 413296
rect 33100 413256 59268 413284
rect 33100 413244 33106 413256
rect 59262 413244 59268 413256
rect 59320 413284 59326 413296
rect 66254 413284 66260 413296
rect 59320 413256 66260 413284
rect 59320 413244 59326 413256
rect 66254 413244 66260 413256
rect 66312 413244 66318 413296
rect 128354 413244 128360 413296
rect 128412 413284 128418 413296
rect 140774 413284 140780 413296
rect 128412 413256 140780 413284
rect 128412 413244 128418 413256
rect 140774 413244 140780 413256
rect 140832 413244 140838 413296
rect 115842 412020 115848 412072
rect 115900 412060 115906 412072
rect 120350 412060 120356 412072
rect 115900 412032 120356 412060
rect 115900 412020 115906 412032
rect 120350 412020 120356 412032
rect 120408 412060 120414 412072
rect 129734 412060 129740 412072
rect 120408 412032 129740 412060
rect 120408 412020 120414 412032
rect 129734 412020 129740 412032
rect 129792 412020 129798 412072
rect 115842 410524 115848 410576
rect 115900 410564 115906 410576
rect 117498 410564 117504 410576
rect 115900 410536 117504 410564
rect 115900 410524 115906 410536
rect 117498 410524 117504 410536
rect 117556 410564 117562 410576
rect 127066 410564 127072 410576
rect 117556 410536 127072 410564
rect 117556 410524 117562 410536
rect 127066 410524 127072 410536
rect 127124 410524 127130 410576
rect 2866 409844 2872 409896
rect 2924 409884 2930 409896
rect 7558 409884 7564 409896
rect 2924 409856 7564 409884
rect 2924 409844 2930 409856
rect 7558 409844 7564 409856
rect 7616 409844 7622 409896
rect 49602 409844 49608 409896
rect 49660 409884 49666 409896
rect 52270 409884 52276 409896
rect 49660 409856 52276 409884
rect 49660 409844 49666 409856
rect 52270 409844 52276 409856
rect 52328 409884 52334 409896
rect 66806 409884 66812 409896
rect 52328 409856 66812 409884
rect 52328 409844 52334 409856
rect 66806 409844 66812 409856
rect 66864 409844 66870 409896
rect 50798 408484 50804 408536
rect 50856 408524 50862 408536
rect 66622 408524 66628 408536
rect 50856 408496 66628 408524
rect 50856 408484 50862 408496
rect 66622 408484 66628 408496
rect 66680 408484 66686 408536
rect 115842 408484 115848 408536
rect 115900 408524 115906 408536
rect 147674 408524 147680 408536
rect 115900 408496 147680 408524
rect 115900 408484 115906 408496
rect 147674 408484 147680 408496
rect 147732 408484 147738 408536
rect 66806 407164 66812 407176
rect 41340 407136 66812 407164
rect 37090 407056 37096 407108
rect 37148 407096 37154 407108
rect 41230 407096 41236 407108
rect 37148 407068 41236 407096
rect 37148 407056 37154 407068
rect 41230 407056 41236 407068
rect 41288 407096 41294 407108
rect 41340 407096 41368 407136
rect 66806 407124 66812 407136
rect 66864 407124 66870 407176
rect 115842 407124 115848 407176
rect 115900 407164 115906 407176
rect 149054 407164 149060 407176
rect 115900 407136 149060 407164
rect 115900 407124 115906 407136
rect 149054 407124 149060 407136
rect 149112 407124 149118 407176
rect 41288 407068 41368 407096
rect 41288 407056 41294 407068
rect 115566 405628 115572 405680
rect 115624 405668 115630 405680
rect 132586 405668 132592 405680
rect 115624 405640 132592 405668
rect 115624 405628 115630 405640
rect 132586 405628 132592 405640
rect 132644 405668 132650 405680
rect 133782 405668 133788 405680
rect 132644 405640 133788 405668
rect 132644 405628 132650 405640
rect 133782 405628 133788 405640
rect 133840 405628 133846 405680
rect 39850 404948 39856 405000
rect 39908 404988 39914 405000
rect 59078 404988 59084 405000
rect 39908 404960 59084 404988
rect 39908 404948 39914 404960
rect 59078 404948 59084 404960
rect 59136 404948 59142 405000
rect 115842 404948 115848 405000
rect 115900 404988 115906 405000
rect 126974 404988 126980 405000
rect 115900 404960 126980 404988
rect 115900 404948 115906 404960
rect 126974 404948 126980 404960
rect 127032 404988 127038 405000
rect 127434 404988 127440 405000
rect 127032 404960 127440 404988
rect 127032 404948 127038 404960
rect 127434 404948 127440 404960
rect 127492 404948 127498 405000
rect 133782 404948 133788 405000
rect 133840 404988 133846 405000
rect 146294 404988 146300 405000
rect 133840 404960 146300 404988
rect 133840 404948 133846 404960
rect 146294 404948 146300 404960
rect 146352 404948 146358 405000
rect 64782 404336 64788 404388
rect 64840 404376 64846 404388
rect 66806 404376 66812 404388
rect 64840 404348 66812 404376
rect 64840 404336 64846 404348
rect 66806 404336 66812 404348
rect 66864 404336 66870 404388
rect 66346 404268 66352 404320
rect 66404 404308 66410 404320
rect 66898 404308 66904 404320
rect 66404 404280 66904 404308
rect 66404 404268 66410 404280
rect 66898 404268 66904 404280
rect 66956 404268 66962 404320
rect 127434 403588 127440 403640
rect 127492 403628 127498 403640
rect 144914 403628 144920 403640
rect 127492 403600 144920 403628
rect 127492 403588 127498 403600
rect 144914 403588 144920 403600
rect 144972 403588 144978 403640
rect 115842 403248 115848 403300
rect 115900 403288 115906 403300
rect 118602 403288 118608 403300
rect 115900 403260 118608 403288
rect 115900 403248 115906 403260
rect 118602 403248 118608 403260
rect 118660 403248 118666 403300
rect 66346 403084 66352 403096
rect 45526 403056 66352 403084
rect 39850 402976 39856 403028
rect 39908 403016 39914 403028
rect 45526 403016 45554 403056
rect 66346 403044 66352 403056
rect 66404 403044 66410 403096
rect 39908 402988 45554 403016
rect 39908 402976 39914 402988
rect 63310 402976 63316 403028
rect 63368 403016 63374 403028
rect 66806 403016 66812 403028
rect 63368 402988 66812 403016
rect 63368 402976 63374 402988
rect 66806 402976 66812 402988
rect 66864 402976 66870 403028
rect 118602 402228 118608 402280
rect 118660 402268 118666 402280
rect 142798 402268 142804 402280
rect 118660 402240 142804 402268
rect 118660 402228 118666 402240
rect 142798 402228 142804 402240
rect 142856 402228 142862 402280
rect 35618 400868 35624 400920
rect 35676 400908 35682 400920
rect 66438 400908 66444 400920
rect 35676 400880 66444 400908
rect 35676 400868 35682 400880
rect 66438 400868 66444 400880
rect 66496 400868 66502 400920
rect 115014 400392 115020 400444
rect 115072 400432 115078 400444
rect 117498 400432 117504 400444
rect 115072 400404 117504 400432
rect 115072 400392 115078 400404
rect 117498 400392 117504 400404
rect 117556 400392 117562 400444
rect 56502 400188 56508 400240
rect 56560 400228 56566 400240
rect 66806 400228 66812 400240
rect 56560 400200 66812 400228
rect 56560 400188 56566 400200
rect 66806 400188 66812 400200
rect 66864 400188 66870 400240
rect 115658 400188 115664 400240
rect 115716 400228 115722 400240
rect 151814 400228 151820 400240
rect 115716 400200 151820 400228
rect 115716 400188 115722 400200
rect 151814 400188 151820 400200
rect 151872 400188 151878 400240
rect 55030 398828 55036 398880
rect 55088 398868 55094 398880
rect 66806 398868 66812 398880
rect 55088 398840 66812 398868
rect 55088 398828 55094 398840
rect 66806 398828 66812 398840
rect 66864 398828 66870 398880
rect 114554 398080 114560 398132
rect 114612 398120 114618 398132
rect 114922 398120 114928 398132
rect 114612 398092 114928 398120
rect 114612 398080 114618 398092
rect 114922 398080 114928 398092
rect 114980 398080 114986 398132
rect 115842 398080 115848 398132
rect 115900 398120 115906 398132
rect 125686 398120 125692 398132
rect 115900 398092 125692 398120
rect 115900 398080 115906 398092
rect 125686 398080 125692 398092
rect 125744 398080 125750 398132
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 21450 397508 21456 397520
rect 3476 397480 21456 397508
rect 3476 397468 3482 397480
rect 21450 397468 21456 397480
rect 21508 397468 21514 397520
rect 42610 396720 42616 396772
rect 42668 396760 42674 396772
rect 60642 396760 60648 396772
rect 42668 396732 60648 396760
rect 42668 396720 42674 396732
rect 60642 396720 60648 396732
rect 60700 396760 60706 396772
rect 66806 396760 66812 396772
rect 60700 396732 66812 396760
rect 60700 396720 60706 396732
rect 66806 396720 66812 396732
rect 66864 396720 66870 396772
rect 115842 396720 115848 396772
rect 115900 396760 115906 396772
rect 124122 396760 124128 396772
rect 115900 396732 124128 396760
rect 115900 396720 115906 396732
rect 124122 396720 124128 396732
rect 124180 396720 124186 396772
rect 59078 396108 59084 396160
rect 59136 396148 59142 396160
rect 66806 396148 66812 396160
rect 59136 396120 66812 396148
rect 59136 396108 59142 396120
rect 66806 396108 66812 396120
rect 66864 396108 66870 396160
rect 115842 396040 115848 396092
rect 115900 396080 115906 396092
rect 131114 396080 131120 396092
rect 115900 396052 131120 396080
rect 115900 396040 115906 396052
rect 131114 396040 131120 396052
rect 131172 396040 131178 396092
rect 48038 395292 48044 395344
rect 48096 395332 48102 395344
rect 64690 395332 64696 395344
rect 48096 395304 64696 395332
rect 48096 395292 48102 395304
rect 64690 395292 64696 395304
rect 64748 395332 64754 395344
rect 66806 395332 66812 395344
rect 64748 395304 66812 395332
rect 64748 395292 64754 395304
rect 66806 395292 66812 395304
rect 66864 395292 66870 395344
rect 115842 394680 115848 394732
rect 115900 394720 115906 394732
rect 191098 394720 191104 394732
rect 115900 394692 191104 394720
rect 115900 394680 115906 394692
rect 191098 394680 191104 394692
rect 191156 394680 191162 394732
rect 64598 393320 64604 393372
rect 64656 393360 64662 393372
rect 66806 393360 66812 393372
rect 64656 393332 66812 393360
rect 64656 393320 64662 393332
rect 66806 393320 66812 393332
rect 66864 393320 66870 393372
rect 115566 393320 115572 393372
rect 115624 393360 115630 393372
rect 187694 393360 187700 393372
rect 115624 393332 187700 393360
rect 115624 393320 115630 393332
rect 187694 393320 187700 393332
rect 187752 393320 187758 393372
rect 115842 393116 115848 393168
rect 115900 393156 115906 393168
rect 118694 393156 118700 393168
rect 115900 393128 118700 393156
rect 115900 393116 115906 393128
rect 118694 393116 118700 393128
rect 118752 393116 118758 393168
rect 118694 392028 118700 392080
rect 118752 392068 118758 392080
rect 122834 392068 122840 392080
rect 118752 392040 122840 392068
rect 118752 392028 118758 392040
rect 122834 392028 122840 392040
rect 122892 392028 122898 392080
rect 57698 391960 57704 392012
rect 57756 392000 57762 392012
rect 66806 392000 66812 392012
rect 57756 391972 66812 392000
rect 57756 391960 57762 391972
rect 66806 391960 66812 391972
rect 66864 391960 66870 392012
rect 115842 391960 115848 392012
rect 115900 392000 115906 392012
rect 147766 392000 147772 392012
rect 115900 391972 147772 392000
rect 115900 391960 115906 391972
rect 147766 391960 147772 391972
rect 147824 391960 147830 392012
rect 63402 391280 63408 391332
rect 63460 391320 63466 391332
rect 63460 391292 85712 391320
rect 63460 391280 63466 391292
rect 48130 391212 48136 391264
rect 48188 391252 48194 391264
rect 48188 391224 80054 391252
rect 48188 391212 48194 391224
rect 80026 390912 80054 391224
rect 85684 391048 85712 391292
rect 117406 391252 117412 391264
rect 113146 391224 117412 391252
rect 87966 391048 87972 391060
rect 85684 391020 87972 391048
rect 87966 391008 87972 391020
rect 88024 391008 88030 391060
rect 99466 391048 99472 391060
rect 89686 391020 99472 391048
rect 89686 390912 89714 391020
rect 99466 391008 99472 391020
rect 99524 391008 99530 391060
rect 106642 391008 106648 391060
rect 106700 391048 106706 391060
rect 113146 391048 113174 391224
rect 117406 391212 117412 391224
rect 117464 391252 117470 391264
rect 128354 391252 128360 391264
rect 117464 391224 128360 391252
rect 117464 391212 117470 391224
rect 128354 391212 128360 391224
rect 128412 391212 128418 391264
rect 106700 391020 113174 391048
rect 106700 391008 106706 391020
rect 89898 390940 89904 390992
rect 89956 390980 89962 390992
rect 92934 390980 92940 390992
rect 89956 390952 92940 390980
rect 89956 390940 89962 390952
rect 92934 390940 92940 390952
rect 92992 390940 92998 390992
rect 80026 390884 89714 390912
rect 112162 390668 112168 390720
rect 112220 390708 112226 390720
rect 112714 390708 112720 390720
rect 112220 390680 112720 390708
rect 112220 390668 112226 390680
rect 112714 390668 112720 390680
rect 112772 390668 112778 390720
rect 88242 390260 88248 390312
rect 88300 390300 88306 390312
rect 88978 390300 88984 390312
rect 88300 390272 88984 390300
rect 88300 390260 88306 390272
rect 88978 390260 88984 390272
rect 89036 390260 89042 390312
rect 67634 390124 67640 390176
rect 67692 390164 67698 390176
rect 68784 390164 68790 390176
rect 67692 390136 68790 390164
rect 67692 390124 67698 390136
rect 68784 390124 68790 390136
rect 68842 390124 68848 390176
rect 41322 389852 41328 389904
rect 41380 389892 41386 389904
rect 53834 389892 53840 389904
rect 41380 389864 53840 389892
rect 41380 389852 41386 389864
rect 53834 389852 53840 389864
rect 53892 389852 53898 389904
rect 21358 389784 21364 389836
rect 21416 389824 21422 389836
rect 99190 389824 99196 389836
rect 21416 389796 99196 389824
rect 21416 389784 21422 389796
rect 99190 389784 99196 389796
rect 99248 389824 99254 389836
rect 100754 389824 100760 389836
rect 99248 389796 100760 389824
rect 99248 389784 99254 389796
rect 100754 389784 100760 389796
rect 100812 389784 100818 389836
rect 104802 389784 104808 389836
rect 104860 389824 104866 389836
rect 114922 389824 114928 389836
rect 104860 389796 114928 389824
rect 104860 389784 104866 389796
rect 114922 389784 114928 389796
rect 114980 389784 114986 389836
rect 53834 389172 53840 389224
rect 53892 389212 53898 389224
rect 54754 389212 54760 389224
rect 53892 389184 54760 389212
rect 53892 389172 53898 389184
rect 54754 389172 54760 389184
rect 54812 389212 54818 389224
rect 82998 389212 83004 389224
rect 54812 389184 83004 389212
rect 54812 389172 54818 389184
rect 82998 389172 83004 389184
rect 83056 389172 83062 389224
rect 65978 389104 65984 389156
rect 66036 389144 66042 389156
rect 72510 389144 72516 389156
rect 66036 389116 72516 389144
rect 66036 389104 66042 389116
rect 72510 389104 72516 389116
rect 72568 389104 72574 389156
rect 101674 389104 101680 389156
rect 101732 389144 101738 389156
rect 106642 389144 106648 389156
rect 101732 389116 106648 389144
rect 101732 389104 101738 389116
rect 106642 389104 106648 389116
rect 106700 389104 106706 389156
rect 110138 389104 110144 389156
rect 110196 389144 110202 389156
rect 121454 389144 121460 389156
rect 110196 389116 121460 389144
rect 110196 389104 110202 389116
rect 121454 389104 121460 389116
rect 121512 389104 121518 389156
rect 46658 388424 46664 388476
rect 46716 388464 46722 388476
rect 65978 388464 65984 388476
rect 46716 388436 65984 388464
rect 46716 388424 46722 388436
rect 65978 388424 65984 388436
rect 66036 388424 66042 388476
rect 91094 388424 91100 388476
rect 91152 388464 91158 388476
rect 100018 388464 100024 388476
rect 91152 388436 100024 388464
rect 91152 388424 91158 388436
rect 100018 388424 100024 388436
rect 100076 388424 100082 388476
rect 103698 388424 103704 388476
rect 103756 388464 103762 388476
rect 232498 388464 232504 388476
rect 103756 388436 232504 388464
rect 103756 388424 103762 388436
rect 232498 388424 232504 388436
rect 232556 388424 232562 388476
rect 93394 388288 93400 388340
rect 93452 388328 93458 388340
rect 95878 388328 95884 388340
rect 93452 388300 95884 388328
rect 93452 388288 93458 388300
rect 95878 388288 95884 388300
rect 95936 388288 95942 388340
rect 85390 387812 85396 387864
rect 85448 387852 85454 387864
rect 90358 387852 90364 387864
rect 85448 387824 90364 387852
rect 85448 387812 85454 387824
rect 90358 387812 90364 387824
rect 90416 387812 90422 387864
rect 44082 387744 44088 387796
rect 44140 387784 44146 387796
rect 55122 387784 55128 387796
rect 44140 387756 55128 387784
rect 44140 387744 44146 387756
rect 55122 387744 55128 387756
rect 55180 387784 55186 387796
rect 73982 387784 73988 387796
rect 55180 387756 73988 387784
rect 55180 387744 55186 387756
rect 73982 387744 73988 387756
rect 74040 387744 74046 387796
rect 74258 387744 74264 387796
rect 74316 387784 74322 387796
rect 75270 387784 75276 387796
rect 74316 387756 75276 387784
rect 74316 387744 74322 387756
rect 75270 387744 75276 387756
rect 75328 387744 75334 387796
rect 79870 387744 79876 387796
rect 79928 387784 79934 387796
rect 81526 387784 81532 387796
rect 79928 387756 81532 387784
rect 79928 387744 79934 387756
rect 81526 387744 81532 387756
rect 81584 387744 81590 387796
rect 120718 387744 120724 387796
rect 120776 387784 120782 387796
rect 121454 387784 121460 387796
rect 120776 387756 121460 387784
rect 120776 387744 120782 387756
rect 121454 387744 121460 387756
rect 121512 387744 121518 387796
rect 76558 387608 76564 387660
rect 76616 387648 76622 387660
rect 80054 387648 80060 387660
rect 76616 387620 80060 387648
rect 76616 387608 76622 387620
rect 80054 387608 80060 387620
rect 80112 387608 80118 387660
rect 86862 387064 86868 387116
rect 86920 387104 86926 387116
rect 120718 387104 120724 387116
rect 86920 387076 120724 387104
rect 86920 387064 86926 387076
rect 120718 387064 120724 387076
rect 120776 387064 120782 387116
rect 69014 386996 69020 387048
rect 69072 387036 69078 387048
rect 69750 387036 69756 387048
rect 69072 387008 69756 387036
rect 69072 386996 69078 387008
rect 69750 386996 69756 387008
rect 69808 386996 69814 387048
rect 77294 386996 77300 387048
rect 77352 387036 77358 387048
rect 78030 387036 78036 387048
rect 77352 387008 78036 387036
rect 77352 386996 77358 387008
rect 78030 386996 78036 387008
rect 78088 386996 78094 387048
rect 93854 386996 93860 387048
rect 93912 387036 93918 387048
rect 94774 387036 94780 387048
rect 93912 387008 94780 387036
rect 93912 386996 93918 387008
rect 94774 386996 94780 387008
rect 94832 386996 94838 387048
rect 111794 386996 111800 387048
rect 111852 387036 111858 387048
rect 112254 387036 112260 387048
rect 111852 387008 112260 387036
rect 111852 386996 111858 387008
rect 112254 386996 112260 387008
rect 112312 386996 112318 387048
rect 46842 386316 46848 386368
rect 46900 386356 46906 386368
rect 96614 386356 96620 386368
rect 46900 386328 96620 386356
rect 46900 386316 46906 386328
rect 96614 386316 96620 386328
rect 96672 386356 96678 386368
rect 97902 386356 97908 386368
rect 96672 386328 97908 386356
rect 96672 386316 96678 386328
rect 97902 386316 97908 386328
rect 97960 386316 97966 386368
rect 105170 386316 105176 386368
rect 105228 386356 105234 386368
rect 133874 386356 133880 386368
rect 105228 386328 133880 386356
rect 105228 386316 105234 386328
rect 133874 386316 133880 386328
rect 133932 386356 133938 386368
rect 136634 386356 136640 386368
rect 133932 386328 136640 386356
rect 133932 386316 133938 386328
rect 136634 386316 136640 386328
rect 136692 386316 136698 386368
rect 80882 386248 80888 386300
rect 80940 386288 80946 386300
rect 81342 386288 81348 386300
rect 80940 386260 81348 386288
rect 80940 386248 80946 386260
rect 81342 386248 81348 386260
rect 81400 386288 81406 386300
rect 115934 386288 115940 386300
rect 81400 386260 115940 386288
rect 81400 386248 81406 386260
rect 115934 386248 115940 386260
rect 115992 386248 115998 386300
rect 108666 384956 108672 385008
rect 108724 384996 108730 385008
rect 125870 384996 125876 385008
rect 108724 384968 125876 384996
rect 108724 384956 108730 384968
rect 125870 384956 125876 384968
rect 125928 384996 125934 385008
rect 126882 384996 126888 385008
rect 125928 384968 126888 384996
rect 125928 384956 125934 384968
rect 126882 384956 126888 384968
rect 126940 384956 126946 385008
rect 101398 384344 101404 384396
rect 101456 384384 101462 384396
rect 113174 384384 113180 384396
rect 101456 384356 113180 384384
rect 101456 384344 101462 384356
rect 113174 384344 113180 384356
rect 113232 384344 113238 384396
rect 57882 384276 57888 384328
rect 57940 384316 57946 384328
rect 104894 384316 104900 384328
rect 57940 384288 104900 384316
rect 57940 384276 57946 384288
rect 104894 384276 104900 384288
rect 104952 384276 104958 384328
rect 35802 383596 35808 383648
rect 35860 383636 35866 383648
rect 91830 383636 91836 383648
rect 35860 383608 91836 383636
rect 35860 383596 35866 383608
rect 91830 383596 91836 383608
rect 91888 383596 91894 383648
rect 77386 382984 77392 383036
rect 77444 383024 77450 383036
rect 106918 383024 106924 383036
rect 77444 382996 106924 383024
rect 77444 382984 77450 382996
rect 106918 382984 106924 382996
rect 106976 382984 106982 383036
rect 97902 382916 97908 382968
rect 97960 382956 97966 382968
rect 126974 382956 126980 382968
rect 97960 382928 126980 382956
rect 97960 382916 97966 382928
rect 126974 382916 126980 382928
rect 127032 382916 127038 382968
rect 91186 382440 91192 382492
rect 91244 382480 91250 382492
rect 91830 382480 91836 382492
rect 91244 382452 91836 382480
rect 91244 382440 91250 382452
rect 91830 382440 91836 382452
rect 91888 382440 91894 382492
rect 34422 382168 34428 382220
rect 34480 382208 34486 382220
rect 96706 382208 96712 382220
rect 34480 382180 96712 382208
rect 34480 382168 34486 382180
rect 96706 382168 96712 382180
rect 96764 382168 96770 382220
rect 96706 381556 96712 381608
rect 96764 381596 96770 381608
rect 117406 381596 117412 381608
rect 96764 381568 117412 381596
rect 96764 381556 96770 381568
rect 117406 381556 117412 381568
rect 117464 381556 117470 381608
rect 73062 381488 73068 381540
rect 73120 381528 73126 381540
rect 77478 381528 77484 381540
rect 73120 381500 77484 381528
rect 73120 381488 73126 381500
rect 77478 381488 77484 381500
rect 77536 381488 77542 381540
rect 107470 381488 107476 381540
rect 107528 381528 107534 381540
rect 139394 381528 139400 381540
rect 107528 381500 139400 381528
rect 107528 381488 107534 381500
rect 139394 381488 139400 381500
rect 139452 381488 139458 381540
rect 38562 380128 38568 380180
rect 38620 380168 38626 380180
rect 69106 380168 69112 380180
rect 38620 380140 69112 380168
rect 38620 380128 38626 380140
rect 69106 380128 69112 380140
rect 69164 380128 69170 380180
rect 93210 380128 93216 380180
rect 93268 380168 93274 380180
rect 115934 380168 115940 380180
rect 93268 380140 115940 380168
rect 93268 380128 93274 380140
rect 115934 380128 115940 380140
rect 115992 380128 115998 380180
rect 103514 378836 103520 378888
rect 103572 378876 103578 378888
rect 138014 378876 138020 378888
rect 103572 378848 138020 378876
rect 103572 378836 103578 378848
rect 138014 378836 138020 378848
rect 138072 378836 138078 378888
rect 21450 378768 21456 378820
rect 21508 378808 21514 378820
rect 114462 378808 114468 378820
rect 21508 378780 114468 378808
rect 21508 378768 21514 378780
rect 114462 378768 114468 378780
rect 114520 378808 114526 378820
rect 116210 378808 116216 378820
rect 114520 378780 116216 378808
rect 114520 378768 114526 378780
rect 116210 378768 116216 378780
rect 116268 378768 116274 378820
rect 95142 378224 95148 378276
rect 95200 378264 95206 378276
rect 102318 378264 102324 378276
rect 95200 378236 102324 378264
rect 95200 378224 95206 378236
rect 102318 378224 102324 378236
rect 102376 378224 102382 378276
rect 97902 377408 97908 377460
rect 97960 377448 97966 377460
rect 120258 377448 120264 377460
rect 97960 377420 120264 377448
rect 97960 377408 97966 377420
rect 120258 377408 120264 377420
rect 120316 377408 120322 377460
rect 92382 376048 92388 376100
rect 92440 376088 92446 376100
rect 97534 376088 97540 376100
rect 92440 376060 97540 376088
rect 92440 376048 92446 376060
rect 97534 376048 97540 376060
rect 97592 376048 97598 376100
rect 104250 376048 104256 376100
rect 104308 376088 104314 376100
rect 123018 376088 123024 376100
rect 104308 376060 123024 376088
rect 104308 376048 104314 376060
rect 123018 376048 123024 376060
rect 123076 376048 123082 376100
rect 48130 375980 48136 376032
rect 48188 376020 48194 376032
rect 76006 376020 76012 376032
rect 48188 375992 76012 376020
rect 48188 375980 48194 375992
rect 76006 375980 76012 375992
rect 76064 375980 76070 376032
rect 83458 375980 83464 376032
rect 83516 376020 83522 376032
rect 105538 376020 105544 376032
rect 83516 375992 105544 376020
rect 83516 375980 83522 375992
rect 105538 375980 105544 375992
rect 105596 375980 105602 376032
rect 101950 374620 101956 374672
rect 102008 374660 102014 374672
rect 113450 374660 113456 374672
rect 102008 374632 113456 374660
rect 102008 374620 102014 374632
rect 113450 374620 113456 374632
rect 113508 374620 113514 374672
rect 93946 373260 93952 373312
rect 94004 373300 94010 373312
rect 124306 373300 124312 373312
rect 94004 373272 124312 373300
rect 94004 373260 94010 373272
rect 124306 373260 124312 373272
rect 124364 373260 124370 373312
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 106090 371260 106096 371272
rect 3476 371232 106096 371260
rect 3476 371220 3482 371232
rect 106090 371220 106096 371232
rect 106148 371260 106154 371272
rect 106148 371232 106228 371260
rect 106148 371220 106154 371232
rect 106200 371192 106228 371232
rect 116118 371192 116124 371204
rect 106200 371164 116124 371192
rect 116118 371152 116124 371164
rect 116176 371152 116182 371204
rect 93854 370472 93860 370524
rect 93912 370512 93918 370524
rect 126238 370512 126244 370524
rect 93912 370484 126244 370512
rect 93912 370472 93918 370484
rect 126238 370472 126244 370484
rect 126296 370472 126302 370524
rect 86770 367752 86776 367804
rect 86828 367792 86834 367804
rect 117314 367792 117320 367804
rect 86828 367764 117320 367792
rect 86828 367752 86834 367764
rect 117314 367752 117320 367764
rect 117372 367752 117378 367804
rect 90358 366324 90364 366376
rect 90416 366364 90422 366376
rect 117958 366364 117964 366376
rect 90416 366336 117964 366364
rect 90416 366324 90422 366336
rect 117958 366324 117964 366336
rect 118016 366324 118022 366376
rect 88978 364964 88984 365016
rect 89036 365004 89042 365016
rect 121454 365004 121460 365016
rect 89036 364976 121460 365004
rect 89036 364964 89042 364976
rect 121454 364964 121460 364976
rect 121512 364964 121518 365016
rect 93118 363604 93124 363656
rect 93176 363644 93182 363656
rect 119062 363644 119068 363656
rect 93176 363616 119068 363644
rect 93176 363604 93182 363616
rect 119062 363604 119068 363616
rect 119120 363604 119126 363656
rect 95050 362176 95056 362228
rect 95108 362216 95114 362228
rect 118878 362216 118884 362228
rect 95108 362188 118884 362216
rect 95108 362176 95114 362188
rect 118878 362176 118884 362188
rect 118936 362176 118942 362228
rect 89438 359456 89444 359508
rect 89496 359496 89502 359508
rect 124398 359496 124404 359508
rect 89496 359468 124404 359496
rect 89496 359456 89502 359468
rect 124398 359456 124404 359468
rect 124456 359456 124462 359508
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 17218 358748 17224 358760
rect 3384 358720 17224 358748
rect 3384 358708 3390 358720
rect 17218 358708 17224 358720
rect 17276 358708 17282 358760
rect 84102 356668 84108 356720
rect 84160 356708 84166 356720
rect 112438 356708 112444 356720
rect 84160 356680 112444 356708
rect 84160 356668 84166 356680
rect 112438 356668 112444 356680
rect 112496 356668 112502 356720
rect 85574 353948 85580 354000
rect 85632 353988 85638 354000
rect 104158 353988 104164 354000
rect 85632 353960 104164 353988
rect 85632 353948 85638 353960
rect 104158 353948 104164 353960
rect 104216 353948 104222 354000
rect 113818 349120 113824 349172
rect 113876 349160 113882 349172
rect 260098 349160 260104 349172
rect 113876 349132 260104 349160
rect 113876 349120 113882 349132
rect 260098 349120 260104 349132
rect 260156 349120 260162 349172
rect 93118 346400 93124 346452
rect 93176 346440 93182 346452
rect 93670 346440 93676 346452
rect 93176 346412 93676 346440
rect 93176 346400 93182 346412
rect 93670 346400 93676 346412
rect 93728 346440 93734 346452
rect 272058 346440 272064 346452
rect 93728 346412 272064 346440
rect 93728 346400 93734 346412
rect 272058 346400 272064 346412
rect 272116 346400 272122 346452
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 11698 345080 11704 345092
rect 3384 345052 11704 345080
rect 3384 345040 3390 345052
rect 11698 345040 11704 345052
rect 11756 345040 11762 345092
rect 141418 345040 141424 345092
rect 141476 345080 141482 345092
rect 270586 345080 270592 345092
rect 141476 345052 270592 345080
rect 141476 345040 141482 345052
rect 270586 345040 270592 345052
rect 270644 345040 270650 345092
rect 123478 343680 123484 343732
rect 123536 343720 123542 343732
rect 269114 343720 269120 343732
rect 123536 343692 269120 343720
rect 123536 343680 123542 343692
rect 269114 343680 269120 343692
rect 269172 343680 269178 343732
rect 73798 343612 73804 343664
rect 73856 343652 73862 343664
rect 240134 343652 240140 343664
rect 73856 343624 240140 343652
rect 73856 343612 73862 343624
rect 240134 343612 240140 343624
rect 240192 343612 240198 343664
rect 66990 342252 66996 342304
rect 67048 342292 67054 342304
rect 67450 342292 67456 342304
rect 67048 342264 67456 342292
rect 67048 342252 67054 342264
rect 67450 342252 67456 342264
rect 67508 342292 67514 342304
rect 261478 342292 261484 342304
rect 67508 342264 261484 342292
rect 67508 342252 67514 342264
rect 261478 342252 261484 342264
rect 261536 342252 261542 342304
rect 151078 340960 151084 341012
rect 151136 341000 151142 341012
rect 271966 341000 271972 341012
rect 151136 340972 271972 341000
rect 151136 340960 151142 340972
rect 271966 340960 271972 340972
rect 272024 340960 272030 341012
rect 75270 340892 75276 340944
rect 75328 340932 75334 340944
rect 253290 340932 253296 340944
rect 75328 340904 253296 340932
rect 75328 340892 75334 340904
rect 253290 340892 253296 340904
rect 253348 340892 253354 340944
rect 142798 339532 142804 339584
rect 142856 339572 142862 339584
rect 240410 339572 240416 339584
rect 142856 339544 240416 339572
rect 142856 339532 142862 339544
rect 240410 339532 240416 339544
rect 240468 339532 240474 339584
rect 45278 339464 45284 339516
rect 45336 339504 45342 339516
rect 81434 339504 81440 339516
rect 45336 339476 81440 339504
rect 45336 339464 45342 339476
rect 81434 339464 81440 339476
rect 81492 339464 81498 339516
rect 83550 339464 83556 339516
rect 83608 339504 83614 339516
rect 266446 339504 266452 339516
rect 83608 339476 266452 339504
rect 83608 339464 83614 339476
rect 266446 339464 266452 339476
rect 266504 339464 266510 339516
rect 81434 338716 81440 338768
rect 81492 338756 81498 338768
rect 251174 338756 251180 338768
rect 81492 338728 251180 338756
rect 81492 338716 81498 338728
rect 251174 338716 251180 338728
rect 251232 338716 251238 338768
rect 97810 338104 97816 338156
rect 97868 338144 97874 338156
rect 242158 338144 242164 338156
rect 97868 338116 242164 338144
rect 97868 338104 97874 338116
rect 242158 338104 242164 338116
rect 242216 338104 242222 338156
rect 69658 336812 69664 336864
rect 69716 336852 69722 336864
rect 246390 336852 246396 336864
rect 69716 336824 246396 336852
rect 69716 336812 69722 336824
rect 246390 336812 246396 336824
rect 246448 336812 246454 336864
rect 53558 336744 53564 336796
rect 53616 336784 53622 336796
rect 249794 336784 249800 336796
rect 53616 336756 249800 336784
rect 53616 336744 53622 336756
rect 249794 336744 249800 336756
rect 249852 336744 249858 336796
rect 39666 335996 39672 336048
rect 39724 336036 39730 336048
rect 74626 336036 74632 336048
rect 39724 336008 74632 336036
rect 39724 335996 39730 336008
rect 74626 335996 74632 336008
rect 74684 336036 74690 336048
rect 238018 336036 238024 336048
rect 74684 336008 238024 336036
rect 74684 335996 74690 336008
rect 238018 335996 238024 336008
rect 238076 335996 238082 336048
rect 92382 335316 92388 335368
rect 92440 335356 92446 335368
rect 191190 335356 191196 335368
rect 92440 335328 191196 335356
rect 92440 335316 92446 335328
rect 191190 335316 191196 335328
rect 191248 335316 191254 335368
rect 95234 334568 95240 334620
rect 95292 334608 95298 334620
rect 122926 334608 122932 334620
rect 95292 334580 122932 334608
rect 95292 334568 95298 334580
rect 122926 334568 122932 334580
rect 122984 334608 122990 334620
rect 123846 334608 123852 334620
rect 122984 334580 123852 334608
rect 122984 334568 122990 334580
rect 123846 334568 123852 334580
rect 123904 334568 123910 334620
rect 123846 334024 123852 334076
rect 123904 334064 123910 334076
rect 233878 334064 233884 334076
rect 123904 334036 233884 334064
rect 123904 334024 123910 334036
rect 233878 334024 233884 334036
rect 233936 334024 233942 334076
rect 88242 333956 88248 334008
rect 88300 333996 88306 334008
rect 240778 333996 240784 334008
rect 88300 333968 240784 333996
rect 88300 333956 88306 333968
rect 240778 333956 240784 333968
rect 240836 333956 240842 334008
rect 89714 333208 89720 333260
rect 89772 333248 89778 333260
rect 120166 333248 120172 333260
rect 89772 333220 120172 333248
rect 89772 333208 89778 333220
rect 120166 333208 120172 333220
rect 120224 333208 120230 333260
rect 120166 332596 120172 332648
rect 120224 332636 120230 332648
rect 247678 332636 247684 332648
rect 120224 332608 247684 332636
rect 120224 332596 120230 332608
rect 247678 332596 247684 332608
rect 247736 332596 247742 332648
rect 80698 331304 80704 331356
rect 80756 331344 80762 331356
rect 81250 331344 81256 331356
rect 80756 331316 81256 331344
rect 80756 331304 80762 331316
rect 81250 331304 81256 331316
rect 81308 331344 81314 331356
rect 241514 331344 241520 331356
rect 81308 331316 241520 331344
rect 81308 331304 81314 331316
rect 241514 331304 241520 331316
rect 241572 331304 241578 331356
rect 101490 331236 101496 331288
rect 101548 331276 101554 331288
rect 101950 331276 101956 331288
rect 101548 331248 101956 331276
rect 101548 331236 101554 331248
rect 101950 331236 101956 331248
rect 102008 331276 102014 331288
rect 269206 331276 269212 331288
rect 102008 331248 269212 331276
rect 102008 331236 102014 331248
rect 269206 331236 269212 331248
rect 269264 331236 269270 331288
rect 42702 330488 42708 330540
rect 42760 330528 42766 330540
rect 66990 330528 66996 330540
rect 42760 330500 66996 330528
rect 42760 330488 42766 330500
rect 66990 330488 66996 330500
rect 67048 330488 67054 330540
rect 99282 329876 99288 329928
rect 99340 329916 99346 329928
rect 226978 329916 226984 329928
rect 99340 329888 226984 329916
rect 99340 329876 99346 329888
rect 226978 329876 226984 329888
rect 227036 329876 227042 329928
rect 53466 329808 53472 329860
rect 53524 329848 53530 329860
rect 53650 329848 53656 329860
rect 53524 329820 53656 329848
rect 53524 329808 53530 329820
rect 53650 329808 53656 329820
rect 53708 329848 53714 329860
rect 267826 329848 267832 329860
rect 53708 329820 267832 329848
rect 53708 329808 53714 329820
rect 267826 329808 267832 329820
rect 267884 329808 267890 329860
rect 89714 329060 89720 329112
rect 89772 329100 89778 329112
rect 123018 329100 123024 329112
rect 89772 329072 123024 329100
rect 89772 329060 89778 329072
rect 123018 329060 123024 329072
rect 123076 329100 123082 329112
rect 259638 329100 259644 329112
rect 123076 329072 259644 329100
rect 123076 329060 123082 329072
rect 259638 329060 259644 329072
rect 259696 329060 259702 329112
rect 100202 328448 100208 328500
rect 100260 328488 100266 328500
rect 100662 328488 100668 328500
rect 100260 328460 100668 328488
rect 100260 328448 100266 328460
rect 100662 328448 100668 328460
rect 100720 328488 100726 328500
rect 242894 328488 242900 328500
rect 100720 328460 242900 328488
rect 100720 328448 100726 328460
rect 242894 328448 242900 328460
rect 242952 328448 242958 328500
rect 63218 328380 63224 328432
rect 63276 328420 63282 328432
rect 63402 328420 63408 328432
rect 63276 328392 63408 328420
rect 63276 328380 63282 328392
rect 63402 328380 63408 328392
rect 63460 328380 63466 328432
rect 38470 328176 38476 328228
rect 38528 328216 38534 328228
rect 39850 328216 39856 328228
rect 38528 328188 39856 328216
rect 38528 328176 38534 328188
rect 39850 328176 39856 328188
rect 39908 328176 39914 328228
rect 39850 327700 39856 327752
rect 39908 327740 39914 327752
rect 67542 327740 67548 327752
rect 39908 327712 67548 327740
rect 39908 327700 39914 327712
rect 67542 327700 67548 327712
rect 67600 327700 67606 327752
rect 80238 327700 80244 327752
rect 80296 327740 80302 327752
rect 89714 327740 89720 327752
rect 80296 327712 89720 327740
rect 80296 327700 80302 327712
rect 89714 327700 89720 327712
rect 89772 327700 89778 327752
rect 115198 327156 115204 327208
rect 115256 327196 115262 327208
rect 246482 327196 246488 327208
rect 115256 327168 246488 327196
rect 115256 327156 115262 327168
rect 246482 327156 246488 327168
rect 246540 327156 246546 327208
rect 63402 327088 63408 327140
rect 63460 327128 63466 327140
rect 266538 327128 266544 327140
rect 63460 327100 266544 327128
rect 63460 327088 63466 327100
rect 266538 327088 266544 327100
rect 266596 327088 266602 327140
rect 108850 326340 108856 326392
rect 108908 326380 108914 326392
rect 116118 326380 116124 326392
rect 108908 326352 116124 326380
rect 108908 326340 108914 326352
rect 116118 326340 116124 326352
rect 116176 326340 116182 326392
rect 116118 325728 116124 325780
rect 116176 325768 116182 325780
rect 254026 325768 254032 325780
rect 116176 325740 254032 325768
rect 116176 325728 116182 325740
rect 254026 325728 254032 325740
rect 254084 325728 254090 325780
rect 78030 325660 78036 325712
rect 78088 325700 78094 325712
rect 84102 325700 84108 325712
rect 78088 325672 84108 325700
rect 78088 325660 78094 325672
rect 84102 325660 84108 325672
rect 84160 325700 84166 325712
rect 255406 325700 255412 325712
rect 84160 325672 255412 325700
rect 84160 325660 84166 325672
rect 255406 325660 255412 325672
rect 255464 325660 255470 325712
rect 128998 324912 129004 324964
rect 129056 324952 129062 324964
rect 151078 324952 151084 324964
rect 129056 324924 151084 324952
rect 129056 324912 129062 324924
rect 151078 324912 151084 324924
rect 151136 324912 151142 324964
rect 192478 324368 192484 324420
rect 192536 324408 192542 324420
rect 208670 324408 208676 324420
rect 192536 324380 208676 324408
rect 192536 324368 192542 324380
rect 208670 324368 208676 324380
rect 208728 324368 208734 324420
rect 49510 324300 49516 324352
rect 49568 324340 49574 324352
rect 258166 324340 258172 324352
rect 49568 324312 258172 324340
rect 49568 324300 49574 324312
rect 258166 324300 258172 324312
rect 258224 324300 258230 324352
rect 291838 324300 291844 324352
rect 291896 324340 291902 324352
rect 580166 324340 580172 324352
rect 291896 324312 580172 324340
rect 291896 324300 291902 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 96522 323552 96528 323604
rect 96580 323592 96586 323604
rect 136726 323592 136732 323604
rect 96580 323564 136732 323592
rect 96580 323552 96586 323564
rect 136726 323552 136732 323564
rect 136784 323592 136790 323604
rect 260926 323592 260932 323604
rect 136784 323564 260932 323592
rect 136784 323552 136790 323564
rect 260926 323552 260932 323564
rect 260984 323552 260990 323604
rect 75362 322940 75368 322992
rect 75420 322980 75426 322992
rect 75822 322980 75828 322992
rect 75420 322952 75828 322980
rect 75420 322940 75426 322952
rect 75822 322940 75828 322952
rect 75880 322980 75886 322992
rect 249058 322980 249064 322992
rect 75880 322952 249064 322980
rect 75880 322940 75886 322952
rect 249058 322940 249064 322952
rect 249116 322940 249122 322992
rect 119338 321920 119344 321972
rect 119396 321960 119402 321972
rect 123478 321960 123484 321972
rect 119396 321932 123484 321960
rect 119396 321920 119402 321932
rect 123478 321920 123484 321932
rect 123536 321920 123542 321972
rect 88150 321716 88156 321768
rect 88208 321756 88214 321768
rect 91186 321756 91192 321768
rect 88208 321728 91192 321756
rect 88208 321716 88214 321728
rect 91186 321716 91192 321728
rect 91244 321716 91250 321768
rect 125502 321648 125508 321700
rect 125560 321688 125566 321700
rect 259546 321688 259552 321700
rect 125560 321660 259552 321688
rect 125560 321648 125566 321660
rect 259546 321648 259552 321660
rect 259604 321648 259610 321700
rect 108850 321580 108856 321632
rect 108908 321620 108914 321632
rect 111886 321620 111892 321632
rect 108908 321592 111892 321620
rect 108908 321580 108914 321592
rect 111886 321580 111892 321592
rect 111944 321620 111950 321632
rect 265158 321620 265164 321632
rect 111944 321592 265164 321620
rect 111944 321580 111950 321592
rect 265158 321580 265164 321592
rect 265216 321580 265222 321632
rect 4798 320832 4804 320884
rect 4856 320872 4862 320884
rect 18598 320872 18604 320884
rect 4856 320844 18604 320872
rect 4856 320832 4862 320844
rect 18598 320832 18604 320844
rect 18656 320832 18662 320884
rect 113910 320628 113916 320680
rect 113968 320668 113974 320680
rect 114462 320668 114468 320680
rect 113968 320640 114468 320668
rect 113968 320628 113974 320640
rect 114462 320628 114468 320640
rect 114520 320628 114526 320680
rect 118878 320220 118884 320272
rect 118936 320260 118942 320272
rect 267734 320260 267740 320272
rect 118936 320232 267740 320260
rect 118936 320220 118942 320232
rect 267734 320220 267740 320232
rect 267792 320220 267798 320272
rect 56226 320152 56232 320204
rect 56284 320192 56290 320204
rect 88150 320192 88156 320204
rect 56284 320164 88156 320192
rect 56284 320152 56290 320164
rect 88150 320152 88156 320164
rect 88208 320152 88214 320204
rect 114462 320152 114468 320204
rect 114520 320192 114526 320204
rect 263594 320192 263600 320204
rect 114520 320164 263600 320192
rect 114520 320152 114526 320164
rect 263594 320152 263600 320164
rect 263652 320152 263658 320204
rect 3878 319200 3884 319252
rect 3936 319240 3942 319252
rect 4798 319240 4804 319252
rect 3936 319212 4804 319240
rect 3936 319200 3942 319212
rect 4798 319200 4804 319212
rect 4856 319200 4862 319252
rect 151078 318860 151084 318912
rect 151136 318900 151142 318912
rect 250438 318900 250444 318912
rect 151136 318872 250444 318900
rect 151136 318860 151142 318872
rect 250438 318860 250444 318872
rect 250496 318860 250502 318912
rect 41138 318792 41144 318844
rect 41196 318832 41202 318844
rect 63494 318832 63500 318844
rect 41196 318804 63500 318832
rect 41196 318792 41202 318804
rect 63494 318792 63500 318804
rect 63552 318832 63558 318844
rect 64138 318832 64144 318844
rect 63552 318804 64144 318832
rect 63552 318792 63558 318804
rect 64138 318792 64144 318804
rect 64196 318792 64202 318844
rect 72970 318792 72976 318844
rect 73028 318832 73034 318844
rect 251818 318832 251824 318844
rect 73028 318804 251824 318832
rect 73028 318792 73034 318804
rect 251818 318792 251824 318804
rect 251876 318792 251882 318844
rect 100110 318112 100116 318164
rect 100168 318152 100174 318164
rect 111886 318152 111892 318164
rect 100168 318124 111892 318152
rect 100168 318112 100174 318124
rect 111886 318112 111892 318124
rect 111944 318112 111950 318164
rect 63494 318044 63500 318096
rect 63552 318084 63558 318096
rect 250530 318084 250536 318096
rect 63552 318056 250536 318084
rect 63552 318044 63558 318056
rect 250530 318044 250536 318056
rect 250588 318044 250594 318096
rect 111886 317432 111892 317484
rect 111944 317472 111950 317484
rect 255498 317472 255504 317484
rect 111944 317444 255504 317472
rect 111944 317432 111950 317444
rect 255498 317432 255504 317444
rect 255556 317432 255562 317484
rect 63218 316684 63224 316736
rect 63276 316724 63282 316736
rect 72878 316724 72884 316736
rect 63276 316696 72884 316724
rect 63276 316684 63282 316696
rect 72878 316684 72884 316696
rect 72936 316724 72942 316736
rect 256694 316724 256700 316736
rect 72936 316696 256700 316724
rect 72936 316684 72942 316696
rect 256694 316684 256700 316696
rect 256752 316684 256758 316736
rect 84194 316004 84200 316056
rect 84252 316044 84258 316056
rect 85298 316044 85304 316056
rect 84252 316016 85304 316044
rect 84252 316004 84258 316016
rect 85298 316004 85304 316016
rect 85356 316044 85362 316056
rect 264974 316044 264980 316056
rect 85356 316016 264980 316044
rect 85356 316004 85362 316016
rect 264974 316004 264980 316016
rect 265032 316004 265038 316056
rect 106090 315256 106096 315308
rect 106148 315296 106154 315308
rect 137094 315296 137100 315308
rect 106148 315268 137100 315296
rect 106148 315256 106154 315268
rect 137094 315256 137100 315268
rect 137152 315256 137158 315308
rect 134610 314712 134616 314764
rect 134668 314752 134674 314764
rect 252738 314752 252744 314764
rect 134668 314724 252744 314752
rect 134668 314712 134674 314724
rect 252738 314712 252744 314724
rect 252796 314712 252802 314764
rect 136726 314644 136732 314696
rect 136784 314684 136790 314696
rect 137094 314684 137100 314696
rect 136784 314656 137100 314684
rect 136784 314644 136790 314656
rect 137094 314644 137100 314656
rect 137152 314684 137158 314696
rect 258350 314684 258356 314696
rect 137152 314656 258356 314684
rect 137152 314644 137158 314656
rect 258350 314644 258356 314656
rect 258408 314644 258414 314696
rect 117774 313896 117780 313948
rect 117832 313936 117838 313948
rect 125778 313936 125784 313948
rect 117832 313908 125784 313936
rect 117832 313896 117838 313908
rect 125778 313896 125784 313908
rect 125836 313936 125842 313948
rect 260834 313936 260840 313948
rect 125836 313908 260840 313936
rect 125836 313896 125842 313908
rect 260834 313896 260840 313908
rect 260892 313896 260898 313948
rect 71682 313284 71688 313336
rect 71740 313324 71746 313336
rect 75178 313324 75184 313336
rect 71740 313296 75184 313324
rect 71740 313284 71746 313296
rect 75178 313284 75184 313296
rect 75236 313324 75242 313336
rect 75822 313324 75828 313336
rect 75236 313296 75828 313324
rect 75236 313284 75242 313296
rect 75822 313284 75828 313296
rect 75880 313284 75886 313336
rect 82906 313284 82912 313336
rect 82964 313324 82970 313336
rect 117314 313324 117320 313336
rect 82964 313296 117320 313324
rect 82964 313284 82970 313296
rect 117314 313284 117320 313296
rect 117372 313324 117378 313336
rect 117774 313324 117780 313336
rect 117372 313296 117780 313324
rect 117372 313284 117378 313296
rect 117774 313284 117780 313296
rect 117832 313284 117838 313336
rect 186958 313284 186964 313336
rect 187016 313324 187022 313336
rect 266630 313324 266636 313336
rect 187016 313296 266636 313324
rect 187016 313284 187022 313296
rect 266630 313284 266636 313296
rect 266688 313284 266694 313336
rect 160738 311924 160744 311976
rect 160796 311964 160802 311976
rect 255314 311964 255320 311976
rect 160796 311936 255320 311964
rect 160796 311924 160802 311936
rect 255314 311924 255320 311936
rect 255372 311924 255378 311976
rect 144178 311856 144184 311908
rect 144236 311896 144242 311908
rect 258074 311896 258080 311908
rect 144236 311868 258080 311896
rect 144236 311856 144242 311868
rect 258074 311856 258080 311868
rect 258132 311856 258138 311908
rect 94590 311108 94596 311160
rect 94648 311148 94654 311160
rect 114462 311148 114468 311160
rect 94648 311120 114468 311148
rect 94648 311108 94654 311120
rect 114462 311108 114468 311120
rect 114520 311108 114526 311160
rect 160830 310564 160836 310616
rect 160888 310604 160894 310616
rect 261018 310604 261024 310616
rect 160888 310576 261024 310604
rect 160888 310564 160894 310576
rect 261018 310564 261024 310576
rect 261076 310564 261082 310616
rect 114462 310496 114468 310548
rect 114520 310536 114526 310548
rect 259730 310536 259736 310548
rect 114520 310508 259736 310536
rect 114520 310496 114526 310508
rect 259730 310496 259736 310508
rect 259788 310496 259794 310548
rect 78122 310428 78128 310480
rect 78180 310468 78186 310480
rect 78582 310468 78588 310480
rect 78180 310440 78588 310468
rect 78180 310428 78186 310440
rect 78582 310428 78588 310440
rect 78640 310428 78646 310480
rect 180058 309816 180064 309868
rect 180116 309856 180122 309868
rect 188338 309856 188344 309868
rect 180116 309828 188344 309856
rect 180116 309816 180122 309828
rect 188338 309816 188344 309828
rect 188396 309816 188402 309868
rect 78122 309748 78128 309800
rect 78180 309788 78186 309800
rect 266354 309788 266360 309800
rect 78180 309760 266360 309788
rect 78180 309748 78186 309760
rect 266354 309748 266360 309760
rect 266412 309748 266418 309800
rect 189718 309136 189724 309188
rect 189776 309176 189782 309188
rect 252830 309176 252836 309188
rect 189776 309148 252836 309176
rect 189776 309136 189782 309148
rect 252830 309136 252836 309148
rect 252888 309136 252894 309188
rect 79870 308388 79876 308440
rect 79928 308428 79934 308440
rect 109310 308428 109316 308440
rect 79928 308400 109316 308428
rect 79928 308388 79934 308400
rect 109310 308388 109316 308400
rect 109368 308388 109374 308440
rect 233878 308388 233884 308440
rect 233936 308428 233942 308440
rect 243906 308428 243912 308440
rect 233936 308400 243912 308428
rect 233936 308388 233942 308400
rect 243906 308388 243912 308400
rect 243964 308388 243970 308440
rect 245010 308388 245016 308440
rect 245068 308428 245074 308440
rect 256970 308428 256976 308440
rect 245068 308400 256976 308428
rect 245068 308388 245074 308400
rect 256970 308388 256976 308400
rect 257028 308388 257034 308440
rect 123478 307844 123484 307896
rect 123536 307884 123542 307896
rect 218238 307884 218244 307896
rect 123536 307856 218244 307884
rect 123536 307844 123542 307856
rect 218238 307844 218244 307856
rect 218296 307844 218302 307896
rect 109310 307776 109316 307828
rect 109368 307816 109374 307828
rect 262490 307816 262496 307828
rect 109368 307788 262496 307816
rect 109368 307776 109374 307788
rect 262490 307776 262496 307788
rect 262548 307776 262554 307828
rect 123110 307708 123116 307760
rect 123168 307748 123174 307760
rect 124214 307748 124220 307760
rect 123168 307720 124220 307748
rect 123168 307708 123174 307720
rect 124214 307708 124220 307720
rect 124272 307708 124278 307760
rect 240778 307708 240784 307760
rect 240836 307748 240842 307760
rect 244458 307748 244464 307760
rect 240836 307720 244464 307748
rect 240836 307708 240842 307720
rect 244458 307708 244464 307720
rect 244516 307708 244522 307760
rect 250438 307708 250444 307760
rect 250496 307748 250502 307760
rect 254118 307748 254124 307760
rect 250496 307720 254124 307748
rect 250496 307708 250502 307720
rect 254118 307708 254124 307720
rect 254176 307708 254182 307760
rect 250530 307640 250536 307692
rect 250588 307680 250594 307692
rect 255590 307680 255596 307692
rect 250588 307652 255596 307680
rect 250588 307640 250594 307652
rect 255590 307640 255596 307652
rect 255648 307640 255654 307692
rect 176010 306416 176016 306468
rect 176068 306456 176074 306468
rect 215938 306456 215944 306468
rect 176068 306428 215944 306456
rect 176068 306416 176074 306428
rect 215938 306416 215944 306428
rect 215996 306416 216002 306468
rect 100662 306348 100668 306400
rect 100720 306388 100726 306400
rect 123110 306388 123116 306400
rect 100720 306360 123116 306388
rect 100720 306348 100726 306360
rect 123110 306348 123116 306360
rect 123168 306348 123174 306400
rect 137278 306348 137284 306400
rect 137336 306388 137342 306400
rect 236362 306388 236368 306400
rect 137336 306360 236368 306388
rect 137336 306348 137342 306360
rect 236362 306348 236368 306360
rect 236420 306348 236426 306400
rect 246390 306348 246396 306400
rect 246448 306388 246454 306400
rect 250346 306388 250352 306400
rect 246448 306360 250352 306388
rect 246448 306348 246454 306360
rect 250346 306348 250352 306360
rect 250404 306348 250410 306400
rect 122834 306280 122840 306332
rect 122892 306320 122898 306332
rect 160738 306320 160744 306332
rect 122892 306292 160744 306320
rect 122892 306280 122898 306292
rect 160738 306280 160744 306292
rect 160796 306280 160802 306332
rect 249058 306008 249064 306060
rect 249116 306048 249122 306060
rect 254210 306048 254216 306060
rect 249116 306020 254216 306048
rect 249116 306008 249122 306020
rect 254210 306008 254216 306020
rect 254268 306008 254274 306060
rect 84102 305600 84108 305652
rect 84160 305640 84166 305652
rect 87046 305640 87052 305652
rect 84160 305612 87052 305640
rect 84160 305600 84166 305612
rect 87046 305600 87052 305612
rect 87104 305600 87110 305652
rect 111058 305600 111064 305652
rect 111116 305640 111122 305652
rect 122834 305640 122840 305652
rect 111116 305612 122840 305640
rect 111116 305600 111122 305612
rect 122834 305600 122840 305612
rect 122892 305600 122898 305652
rect 214558 305600 214564 305652
rect 214616 305640 214622 305652
rect 259454 305640 259460 305652
rect 214616 305612 259460 305640
rect 214616 305600 214622 305612
rect 259454 305600 259460 305612
rect 259512 305600 259518 305652
rect 126238 305396 126244 305448
rect 126296 305436 126302 305448
rect 128538 305436 128544 305448
rect 126296 305408 128544 305436
rect 126296 305396 126302 305408
rect 128538 305396 128544 305408
rect 128596 305396 128602 305448
rect 232498 305124 232504 305176
rect 232556 305164 232562 305176
rect 239858 305164 239864 305176
rect 232556 305136 239864 305164
rect 232556 305124 232562 305136
rect 239858 305124 239864 305136
rect 239916 305124 239922 305176
rect 182818 305056 182824 305108
rect 182876 305096 182882 305108
rect 197262 305096 197268 305108
rect 182876 305068 197268 305096
rect 182876 305056 182882 305068
rect 197262 305056 197268 305068
rect 197320 305056 197326 305108
rect 96430 304988 96436 305040
rect 96488 305028 96494 305040
rect 100202 305028 100208 305040
rect 96488 305000 100208 305028
rect 96488 304988 96494 305000
rect 100202 304988 100208 305000
rect 100260 304988 100266 305040
rect 155402 304988 155408 305040
rect 155460 305028 155466 305040
rect 214190 305028 214196 305040
rect 155460 305000 214196 305028
rect 155460 304988 155466 305000
rect 214190 304988 214196 305000
rect 214248 304988 214254 305040
rect 260098 304988 260104 305040
rect 260156 305028 260162 305040
rect 263870 305028 263876 305040
rect 260156 305000 263876 305028
rect 260156 304988 260162 305000
rect 263870 304988 263876 305000
rect 263928 304988 263934 305040
rect 62022 304920 62028 304972
rect 62080 304960 62086 304972
rect 66898 304960 66904 304972
rect 62080 304932 66904 304960
rect 62080 304920 62086 304932
rect 66898 304920 66904 304932
rect 66956 304960 66962 304972
rect 160830 304960 160836 304972
rect 66956 304932 160836 304960
rect 66956 304920 66962 304932
rect 160830 304920 160836 304932
rect 160888 304920 160894 304972
rect 246298 304444 246304 304496
rect 246356 304484 246362 304496
rect 249702 304484 249708 304496
rect 246356 304456 249708 304484
rect 246356 304444 246362 304456
rect 249702 304444 249708 304456
rect 249760 304444 249766 304496
rect 60366 304240 60372 304292
rect 60424 304280 60430 304292
rect 151078 304280 151084 304292
rect 60424 304252 151084 304280
rect 60424 304240 60430 304252
rect 151078 304240 151084 304252
rect 151136 304240 151142 304292
rect 200086 303844 209774 303872
rect 184198 303696 184204 303748
rect 184256 303736 184262 303748
rect 200086 303736 200114 303844
rect 205450 303736 205456 303748
rect 184256 303708 200114 303736
rect 200316 303708 205456 303736
rect 184256 303696 184262 303708
rect 160738 303628 160744 303680
rect 160796 303668 160802 303680
rect 200316 303668 200344 303708
rect 205450 303696 205456 303708
rect 205508 303696 205514 303748
rect 209746 303736 209774 303844
rect 211246 303736 211252 303748
rect 209746 303708 211252 303736
rect 211246 303696 211252 303708
rect 211304 303696 211310 303748
rect 245102 303696 245108 303748
rect 245160 303736 245166 303748
rect 289078 303736 289084 303748
rect 245160 303708 289084 303736
rect 245160 303696 245166 303708
rect 289078 303696 289084 303708
rect 289136 303696 289142 303748
rect 160796 303640 200344 303668
rect 160796 303628 160802 303640
rect 247402 303628 247408 303680
rect 247460 303668 247466 303680
rect 248322 303668 248328 303680
rect 247460 303640 248328 303668
rect 247460 303628 247466 303640
rect 248322 303628 248328 303640
rect 248380 303628 248386 303680
rect 252646 303628 252652 303680
rect 252704 303668 252710 303680
rect 335998 303668 336004 303680
rect 252704 303640 336004 303668
rect 252704 303628 252710 303640
rect 335998 303628 336004 303640
rect 336056 303628 336062 303680
rect 200298 303560 200304 303612
rect 200356 303600 200362 303612
rect 201126 303600 201132 303612
rect 200356 303572 201132 303600
rect 200356 303560 200362 303572
rect 201126 303560 201132 303572
rect 201184 303560 201190 303612
rect 242802 302880 242808 302932
rect 242860 302920 242866 302932
rect 273254 302920 273260 302932
rect 242860 302892 273260 302920
rect 242860 302880 242866 302892
rect 273254 302880 273260 302892
rect 273312 302880 273318 302932
rect 69750 302268 69756 302320
rect 69808 302308 69814 302320
rect 75822 302308 75828 302320
rect 69808 302280 75828 302308
rect 69808 302268 69814 302280
rect 75822 302268 75828 302280
rect 75880 302268 75886 302320
rect 184290 302268 184296 302320
rect 184348 302308 184354 302320
rect 200206 302308 200212 302320
rect 184348 302280 200212 302308
rect 184348 302268 184354 302280
rect 200206 302268 200212 302280
rect 200264 302268 200270 302320
rect 56502 302200 56508 302252
rect 56560 302240 56566 302252
rect 120902 302240 120908 302252
rect 56560 302212 120908 302240
rect 56560 302200 56566 302212
rect 120902 302200 120908 302212
rect 120960 302200 120966 302252
rect 173158 302200 173164 302252
rect 173216 302240 173222 302252
rect 249150 302240 249156 302252
rect 173216 302212 249156 302240
rect 173216 302200 173222 302212
rect 249150 302200 249156 302212
rect 249208 302200 249214 302252
rect 251818 302200 251824 302252
rect 251876 302240 251882 302252
rect 252922 302240 252928 302252
rect 251876 302212 252928 302240
rect 251876 302200 251882 302212
rect 252922 302200 252928 302212
rect 252980 302200 252986 302252
rect 240134 302132 240140 302184
rect 240192 302172 240198 302184
rect 240962 302172 240968 302184
rect 240192 302144 240968 302172
rect 240192 302132 240198 302144
rect 240962 302132 240968 302144
rect 241020 302132 241026 302184
rect 86862 301452 86868 301504
rect 86920 301492 86926 301504
rect 100110 301492 100116 301504
rect 86920 301464 100116 301492
rect 86920 301452 86926 301464
rect 100110 301452 100116 301464
rect 100168 301452 100174 301504
rect 118050 301452 118056 301504
rect 118108 301492 118114 301504
rect 142798 301492 142804 301504
rect 118108 301464 142804 301492
rect 118108 301452 118114 301464
rect 142798 301452 142804 301464
rect 142856 301452 142862 301504
rect 65978 301248 65984 301300
rect 66036 301288 66042 301300
rect 69014 301288 69020 301300
rect 66036 301260 69020 301288
rect 66036 301248 66042 301260
rect 69014 301248 69020 301260
rect 69072 301248 69078 301300
rect 241330 301112 241336 301164
rect 241388 301152 241394 301164
rect 262582 301152 262588 301164
rect 241388 301124 262588 301152
rect 241388 301112 241394 301124
rect 262582 301112 262588 301124
rect 262640 301112 262646 301164
rect 240778 301044 240784 301096
rect 240836 301084 240842 301096
rect 240836 301056 253244 301084
rect 240836 301044 240842 301056
rect 250622 301016 250628 301028
rect 245948 300988 250628 301016
rect 160830 300908 160836 300960
rect 160888 300948 160894 300960
rect 196342 300948 196348 300960
rect 160888 300920 196348 300948
rect 160888 300908 160894 300920
rect 196342 300908 196348 300920
rect 196400 300908 196406 300960
rect 66070 300840 66076 300892
rect 66128 300880 66134 300892
rect 141418 300880 141424 300892
rect 66128 300852 141424 300880
rect 66128 300840 66134 300852
rect 141418 300840 141424 300852
rect 141476 300840 141482 300892
rect 53742 300772 53748 300824
rect 53800 300812 53806 300824
rect 193490 300812 193496 300824
rect 53800 300784 193496 300812
rect 53800 300772 53806 300784
rect 193490 300772 193496 300784
rect 193548 300772 193554 300824
rect 245948 300812 245976 300988
rect 250622 300976 250628 300988
rect 250680 300976 250686 301028
rect 248046 300908 248052 300960
rect 248104 300908 248110 300960
rect 238726 300784 245976 300812
rect 193674 300092 193680 300144
rect 193732 300132 193738 300144
rect 238726 300132 238754 300784
rect 193732 300104 238754 300132
rect 193732 300092 193738 300104
rect 248064 299724 248092 300908
rect 253216 300880 253244 301056
rect 270494 300880 270500 300892
rect 253216 300852 270500 300880
rect 270494 300840 270500 300852
rect 270552 300840 270558 300892
rect 253198 299724 253204 299736
rect 248064 299696 253204 299724
rect 253198 299684 253204 299696
rect 253256 299684 253262 299736
rect 255682 299548 255688 299600
rect 255740 299588 255746 299600
rect 274634 299588 274640 299600
rect 255740 299560 274640 299588
rect 255740 299548 255746 299560
rect 274634 299548 274640 299560
rect 274692 299548 274698 299600
rect 134518 299480 134524 299532
rect 134576 299520 134582 299532
rect 193582 299520 193588 299532
rect 134576 299492 193588 299520
rect 134576 299480 134582 299492
rect 193582 299480 193588 299492
rect 193640 299480 193646 299532
rect 255866 299480 255872 299532
rect 255924 299520 255930 299532
rect 282178 299520 282184 299532
rect 255924 299492 282184 299520
rect 255924 299480 255930 299492
rect 282178 299480 282184 299492
rect 282236 299480 282242 299532
rect 255774 299412 255780 299464
rect 255832 299452 255838 299464
rect 263686 299452 263692 299464
rect 255832 299424 263692 299452
rect 255832 299412 255838 299424
rect 263686 299412 263692 299424
rect 263744 299412 263750 299464
rect 255682 299344 255688 299396
rect 255740 299384 255746 299396
rect 258258 299384 258264 299396
rect 255740 299356 258264 299384
rect 255740 299344 255746 299356
rect 258258 299344 258264 299356
rect 258316 299384 258322 299396
rect 259362 299384 259368 299396
rect 258316 299356 259368 299384
rect 258316 299344 258322 299356
rect 259362 299344 259368 299356
rect 259420 299344 259426 299396
rect 85758 299072 85764 299124
rect 85816 299112 85822 299124
rect 86770 299112 86776 299124
rect 85816 299084 86776 299112
rect 85816 299072 85822 299084
rect 86770 299072 86776 299084
rect 86828 299072 86834 299124
rect 100018 299004 100024 299056
rect 100076 299044 100082 299056
rect 105630 299044 105636 299056
rect 100076 299016 105636 299044
rect 100076 299004 100082 299016
rect 105630 299004 105636 299016
rect 105688 299004 105694 299056
rect 186314 298868 186320 298920
rect 186372 298908 186378 298920
rect 191742 298908 191748 298920
rect 186372 298880 191748 298908
rect 186372 298868 186378 298880
rect 191742 298868 191748 298880
rect 191800 298868 191806 298920
rect 259362 298732 259368 298784
rect 259420 298772 259426 298784
rect 280890 298772 280896 298784
rect 259420 298744 280896 298772
rect 259420 298732 259426 298744
rect 280890 298732 280896 298744
rect 280948 298732 280954 298784
rect 71038 298596 71044 298648
rect 71096 298636 71102 298648
rect 72602 298636 72608 298648
rect 71096 298608 72608 298636
rect 71096 298596 71102 298608
rect 72602 298596 72608 298608
rect 72660 298596 72666 298648
rect 86770 298120 86776 298172
rect 86828 298160 86834 298172
rect 139486 298160 139492 298172
rect 86828 298132 139492 298160
rect 86828 298120 86834 298132
rect 139486 298120 139492 298132
rect 139544 298120 139550 298172
rect 263686 298120 263692 298172
rect 263744 298160 263750 298172
rect 268470 298160 268476 298172
rect 263744 298132 268476 298160
rect 263744 298120 263750 298132
rect 268470 298120 268476 298132
rect 268528 298120 268534 298172
rect 298738 298120 298744 298172
rect 298796 298160 298802 298172
rect 580166 298160 580172 298172
rect 298796 298132 580172 298160
rect 298796 298120 298802 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 255774 298052 255780 298104
rect 255832 298092 255838 298104
rect 269206 298092 269212 298104
rect 255832 298064 269212 298092
rect 255832 298052 255838 298064
rect 269206 298052 269212 298064
rect 269264 298092 269270 298104
rect 270402 298092 270408 298104
rect 269264 298064 270408 298092
rect 269264 298052 269270 298064
rect 270402 298052 270408 298064
rect 270460 298052 270466 298104
rect 261478 297984 261484 298036
rect 261536 298024 261542 298036
rect 262214 298024 262220 298036
rect 261536 297996 262220 298024
rect 261536 297984 261542 297996
rect 262214 297984 262220 297996
rect 262272 297984 262278 298036
rect 255682 297372 255688 297424
rect 255740 297412 255746 297424
rect 262122 297412 262128 297424
rect 255740 297384 262128 297412
rect 255740 297372 255746 297384
rect 262122 297372 262128 297384
rect 262180 297372 262186 297424
rect 270402 297372 270408 297424
rect 270460 297412 270466 297424
rect 282086 297412 282092 297424
rect 270460 297384 282092 297412
rect 270460 297372 270466 297384
rect 282086 297372 282092 297384
rect 282144 297372 282150 297424
rect 282178 297372 282184 297424
rect 282236 297412 282242 297424
rect 317414 297412 317420 297424
rect 282236 297384 317420 297412
rect 282236 297372 282242 297384
rect 317414 297372 317420 297384
rect 317472 297372 317478 297424
rect 255682 296624 255688 296676
rect 255740 296664 255746 296676
rect 267826 296664 267832 296676
rect 255740 296636 267832 296664
rect 255740 296624 255746 296636
rect 267826 296624 267832 296636
rect 267884 296664 267890 296676
rect 269022 296664 269028 296676
rect 267884 296636 269028 296664
rect 267884 296624 267890 296636
rect 269022 296624 269028 296636
rect 269080 296624 269086 296676
rect 57606 295944 57612 295996
rect 57664 295984 57670 295996
rect 78582 295984 78588 295996
rect 57664 295956 78588 295984
rect 57664 295944 57670 295956
rect 78582 295944 78588 295956
rect 78640 295984 78646 295996
rect 191190 295984 191196 295996
rect 78640 295956 191196 295984
rect 78640 295944 78646 295956
rect 191190 295944 191196 295956
rect 191248 295944 191254 295996
rect 269022 295944 269028 295996
rect 269080 295984 269086 295996
rect 287054 295984 287060 295996
rect 269080 295956 287060 295984
rect 269080 295944 269086 295956
rect 287054 295944 287060 295956
rect 287112 295944 287118 295996
rect 255406 295808 255412 295860
rect 255464 295848 255470 295860
rect 255774 295848 255780 295860
rect 255464 295820 255780 295848
rect 255464 295808 255470 295820
rect 255774 295808 255780 295820
rect 255832 295808 255838 295860
rect 78674 295332 78680 295384
rect 78732 295372 78738 295384
rect 79962 295372 79968 295384
rect 78732 295344 79968 295372
rect 78732 295332 78738 295344
rect 79962 295332 79968 295344
rect 80020 295372 80026 295384
rect 110598 295372 110604 295384
rect 80020 295344 110604 295372
rect 80020 295332 80026 295344
rect 110598 295332 110604 295344
rect 110656 295332 110662 295384
rect 170398 295332 170404 295384
rect 170456 295372 170462 295384
rect 191742 295372 191748 295384
rect 170456 295344 191748 295372
rect 170456 295332 170462 295344
rect 191742 295332 191748 295344
rect 191800 295332 191806 295384
rect 255406 295332 255412 295384
rect 255464 295372 255470 295384
rect 259362 295372 259368 295384
rect 255464 295344 259368 295372
rect 255464 295332 255470 295344
rect 259362 295332 259368 295344
rect 259420 295372 259426 295384
rect 259638 295372 259644 295384
rect 259420 295344 259644 295372
rect 259420 295332 259426 295344
rect 259638 295332 259644 295344
rect 259696 295332 259702 295384
rect 120810 294584 120816 294636
rect 120868 294624 120874 294636
rect 191098 294624 191104 294636
rect 120868 294596 191104 294624
rect 120868 294584 120874 294596
rect 191098 294584 191104 294596
rect 191156 294584 191162 294636
rect 256786 294040 256792 294092
rect 256844 294080 256850 294092
rect 257338 294080 257344 294092
rect 256844 294052 257344 294080
rect 256844 294040 256850 294052
rect 257338 294040 257344 294052
rect 257396 294040 257402 294092
rect 39850 293972 39856 294024
rect 39908 294012 39914 294024
rect 75178 294012 75184 294024
rect 39908 293984 75184 294012
rect 39908 293972 39914 293984
rect 75178 293972 75184 293984
rect 75236 294012 75242 294024
rect 75362 294012 75368 294024
rect 75236 293984 75368 294012
rect 75236 293972 75242 293984
rect 75362 293972 75368 293984
rect 75420 293972 75426 294024
rect 93762 293972 93768 294024
rect 93820 294012 93826 294024
rect 124858 294012 124864 294024
rect 93820 293984 124864 294012
rect 93820 293972 93826 293984
rect 124858 293972 124864 293984
rect 124916 294012 124922 294024
rect 191650 294012 191656 294024
rect 124916 293984 191656 294012
rect 124916 293972 124922 293984
rect 191650 293972 191656 293984
rect 191708 293972 191714 294024
rect 255406 293972 255412 294024
rect 255464 294012 255470 294024
rect 263686 294012 263692 294024
rect 255464 293984 263692 294012
rect 255464 293972 255470 293984
rect 263686 293972 263692 293984
rect 263744 293972 263750 294024
rect 153102 293904 153108 293956
rect 153160 293944 153166 293956
rect 191742 293944 191748 293956
rect 153160 293916 191748 293944
rect 153160 293904 153166 293916
rect 191742 293904 191748 293916
rect 191800 293904 191806 293956
rect 255682 293904 255688 293956
rect 255740 293944 255746 293956
rect 263870 293944 263876 293956
rect 255740 293916 263876 293944
rect 255740 293904 255746 293916
rect 263870 293904 263876 293916
rect 263928 293904 263934 293956
rect 255406 293836 255412 293888
rect 255464 293876 255470 293888
rect 262214 293876 262220 293888
rect 255464 293848 262220 293876
rect 255464 293836 255470 293848
rect 262214 293836 262220 293848
rect 262272 293836 262278 293888
rect 95878 293224 95884 293276
rect 95936 293264 95942 293276
rect 104986 293264 104992 293276
rect 95936 293236 104992 293264
rect 95936 293224 95942 293236
rect 104986 293224 104992 293236
rect 105044 293224 105050 293276
rect 125502 293224 125508 293276
rect 125560 293264 125566 293276
rect 151814 293264 151820 293276
rect 125560 293236 151820 293264
rect 125560 293224 125566 293236
rect 151814 293224 151820 293236
rect 151872 293264 151878 293276
rect 153102 293264 153108 293276
rect 151872 293236 153108 293264
rect 151872 293224 151878 293236
rect 153102 293224 153108 293236
rect 153160 293224 153166 293276
rect 41322 292612 41328 292664
rect 41380 292652 41386 292664
rect 77846 292652 77852 292664
rect 41380 292624 77852 292652
rect 41380 292612 41386 292624
rect 77846 292612 77852 292624
rect 77904 292652 77910 292664
rect 78030 292652 78036 292664
rect 77904 292624 78036 292652
rect 77904 292612 77910 292624
rect 78030 292612 78036 292624
rect 78088 292612 78094 292664
rect 3510 292544 3516 292596
rect 3568 292584 3574 292596
rect 14458 292584 14464 292596
rect 3568 292556 14464 292584
rect 3568 292544 3574 292556
rect 14458 292544 14464 292556
rect 14516 292544 14522 292596
rect 60458 292544 60464 292596
rect 60516 292584 60522 292596
rect 60642 292584 60648 292596
rect 60516 292556 60648 292584
rect 60516 292544 60522 292556
rect 60642 292544 60648 292556
rect 60700 292584 60706 292596
rect 191466 292584 191472 292596
rect 60700 292556 191472 292584
rect 60700 292544 60706 292556
rect 191466 292544 191472 292556
rect 191524 292544 191530 292596
rect 255406 292068 255412 292120
rect 255464 292108 255470 292120
rect 256970 292108 256976 292120
rect 255464 292080 256976 292108
rect 255464 292068 255470 292080
rect 256970 292068 256976 292080
rect 257028 292068 257034 292120
rect 159358 291864 159364 291916
rect 159416 291904 159422 291916
rect 189810 291904 189816 291916
rect 159416 291876 189816 291904
rect 159416 291864 159422 291876
rect 189810 291864 189816 291876
rect 189868 291864 189874 291916
rect 77754 291796 77760 291848
rect 77812 291836 77818 291848
rect 78122 291836 78128 291848
rect 77812 291808 78128 291836
rect 77812 291796 77818 291808
rect 78122 291796 78128 291808
rect 78180 291796 78186 291848
rect 85574 291796 85580 291848
rect 85632 291836 85638 291848
rect 116026 291836 116032 291848
rect 85632 291808 116032 291836
rect 85632 291796 85638 291808
rect 116026 291796 116032 291808
rect 116084 291796 116090 291848
rect 120902 291796 120908 291848
rect 120960 291836 120966 291848
rect 191098 291836 191104 291848
rect 120960 291808 191104 291836
rect 120960 291796 120966 291808
rect 191098 291796 191104 291808
rect 191156 291796 191162 291848
rect 37090 291320 37096 291372
rect 37148 291360 37154 291372
rect 72418 291360 72424 291372
rect 37148 291332 72424 291360
rect 37148 291320 37154 291332
rect 72418 291320 72424 291332
rect 72476 291320 72482 291372
rect 41230 291252 41236 291304
rect 41288 291292 41294 291304
rect 77754 291292 77760 291304
rect 41288 291264 77760 291292
rect 41288 291252 41294 291264
rect 77754 291252 77760 291264
rect 77812 291252 77818 291304
rect 72050 291184 72056 291236
rect 72108 291224 72114 291236
rect 73062 291224 73068 291236
rect 72108 291196 73068 291224
rect 72108 291184 72114 291196
rect 73062 291184 73068 291196
rect 73120 291224 73126 291236
rect 131758 291224 131764 291236
rect 73120 291196 131764 291224
rect 73120 291184 73126 291196
rect 131758 291184 131764 291196
rect 131816 291184 131822 291236
rect 255682 291116 255688 291168
rect 255740 291156 255746 291168
rect 271966 291156 271972 291168
rect 255740 291128 271972 291156
rect 255740 291116 255746 291128
rect 271966 291116 271972 291128
rect 272024 291116 272030 291168
rect 255406 290844 255412 290896
rect 255464 290884 255470 290896
rect 258166 290884 258172 290896
rect 255464 290856 258172 290884
rect 255464 290844 255470 290856
rect 258166 290844 258172 290856
rect 258224 290844 258230 290896
rect 76190 290708 76196 290760
rect 76248 290748 76254 290760
rect 76742 290748 76748 290760
rect 76248 290720 76748 290748
rect 76248 290708 76254 290720
rect 76742 290708 76748 290720
rect 76800 290708 76806 290760
rect 162118 290436 162124 290488
rect 162176 290476 162182 290488
rect 192478 290476 192484 290488
rect 162176 290448 192484 290476
rect 162176 290436 162182 290448
rect 192478 290436 192484 290448
rect 192536 290436 192542 290488
rect 89530 289892 89536 289944
rect 89588 289932 89594 289944
rect 120902 289932 120908 289944
rect 89588 289904 120908 289932
rect 89588 289892 89594 289904
rect 120902 289892 120908 289904
rect 120960 289892 120966 289944
rect 39758 289824 39764 289876
rect 39816 289864 39822 289876
rect 76190 289864 76196 289876
rect 39816 289836 76196 289864
rect 39816 289824 39822 289836
rect 76190 289824 76196 289836
rect 76248 289824 76254 289876
rect 81986 289824 81992 289876
rect 82044 289864 82050 289876
rect 82722 289864 82728 289876
rect 82044 289836 82728 289864
rect 82044 289824 82050 289836
rect 82722 289824 82728 289836
rect 82780 289864 82786 289876
rect 112070 289864 112076 289876
rect 82780 289836 112076 289864
rect 82780 289824 82786 289836
rect 112070 289824 112076 289836
rect 112128 289864 112134 289876
rect 191742 289864 191748 289876
rect 112128 289836 191748 289864
rect 112128 289824 112134 289836
rect 191742 289824 191748 289836
rect 191800 289824 191806 289876
rect 46750 289756 46756 289808
rect 46808 289796 46814 289808
rect 52178 289796 52184 289808
rect 46808 289768 52184 289796
rect 46808 289756 46814 289768
rect 52178 289756 52184 289768
rect 52236 289756 52242 289808
rect 255682 289756 255688 289808
rect 255740 289796 255746 289808
rect 270586 289796 270592 289808
rect 255740 289768 270592 289796
rect 255740 289756 255746 289768
rect 270586 289756 270592 289768
rect 270644 289756 270650 289808
rect 255406 289688 255412 289740
rect 255464 289728 255470 289740
rect 260926 289728 260932 289740
rect 255464 289700 260932 289728
rect 255464 289688 255470 289700
rect 260926 289688 260932 289700
rect 260984 289688 260990 289740
rect 56318 288464 56324 288516
rect 56376 288504 56382 288516
rect 82998 288504 83004 288516
rect 56376 288476 83004 288504
rect 56376 288464 56382 288476
rect 82998 288464 83004 288476
rect 83056 288504 83062 288516
rect 83458 288504 83464 288516
rect 83056 288476 83464 288504
rect 83056 288464 83062 288476
rect 83458 288464 83464 288476
rect 83516 288464 83522 288516
rect 101582 288464 101588 288516
rect 101640 288504 101646 288516
rect 113818 288504 113824 288516
rect 101640 288476 113824 288504
rect 101640 288464 101646 288476
rect 113818 288464 113824 288476
rect 113876 288464 113882 288516
rect 52178 288396 52184 288448
rect 52236 288436 52242 288448
rect 79962 288436 79968 288448
rect 52236 288408 79968 288436
rect 52236 288396 52242 288408
rect 79962 288396 79968 288408
rect 80020 288396 80026 288448
rect 95234 288396 95240 288448
rect 95292 288436 95298 288448
rect 96522 288436 96528 288448
rect 95292 288408 96528 288436
rect 95292 288396 95298 288408
rect 96522 288396 96528 288408
rect 96580 288436 96586 288448
rect 109126 288436 109132 288448
rect 96580 288408 109132 288436
rect 96580 288396 96586 288408
rect 109126 288396 109132 288408
rect 109184 288396 109190 288448
rect 116578 288396 116584 288448
rect 116636 288436 116642 288448
rect 191742 288436 191748 288448
rect 116636 288408 191748 288436
rect 116636 288396 116642 288408
rect 191742 288396 191748 288408
rect 191800 288396 191806 288448
rect 88610 288328 88616 288380
rect 88668 288368 88674 288380
rect 89622 288368 89628 288380
rect 88668 288340 89628 288368
rect 88668 288328 88674 288340
rect 89622 288328 89628 288340
rect 89680 288328 89686 288380
rect 179414 288328 179420 288380
rect 179472 288368 179478 288380
rect 190822 288368 190828 288380
rect 179472 288340 190828 288368
rect 179472 288328 179478 288340
rect 190822 288328 190828 288340
rect 190880 288328 190886 288380
rect 255406 288328 255412 288380
rect 255464 288368 255470 288380
rect 269114 288368 269120 288380
rect 255464 288340 269120 288368
rect 255464 288328 255470 288340
rect 269114 288328 269120 288340
rect 269172 288328 269178 288380
rect 255682 288260 255688 288312
rect 255740 288300 255746 288312
rect 265158 288300 265164 288312
rect 255740 288272 265164 288300
rect 255740 288260 255746 288272
rect 265158 288260 265164 288272
rect 265216 288260 265222 288312
rect 78674 287716 78680 287768
rect 78732 287756 78738 287768
rect 79134 287756 79140 287768
rect 78732 287728 79140 287756
rect 78732 287716 78738 287728
rect 79134 287716 79140 287728
rect 79192 287716 79198 287768
rect 85666 287716 85672 287768
rect 85724 287756 85730 287768
rect 86310 287756 86316 287768
rect 85724 287728 86316 287756
rect 85724 287716 85730 287728
rect 86310 287716 86316 287728
rect 86368 287716 86374 287768
rect 11698 287648 11704 287700
rect 11756 287688 11762 287700
rect 34514 287688 34520 287700
rect 11756 287660 34520 287688
rect 11756 287648 11762 287660
rect 34514 287648 34520 287660
rect 34572 287648 34578 287700
rect 58986 287648 58992 287700
rect 59044 287688 59050 287700
rect 71682 287688 71688 287700
rect 59044 287660 71688 287688
rect 59044 287648 59050 287660
rect 71682 287648 71688 287660
rect 71740 287688 71746 287700
rect 74534 287688 74540 287700
rect 71740 287660 74540 287688
rect 71740 287648 71746 287660
rect 74534 287648 74540 287660
rect 74592 287648 74598 287700
rect 110506 287648 110512 287700
rect 110564 287688 110570 287700
rect 119338 287688 119344 287700
rect 110564 287660 119344 287688
rect 110564 287648 110570 287660
rect 119338 287648 119344 287660
rect 119396 287648 119402 287700
rect 169018 287648 169024 287700
rect 169076 287688 169082 287700
rect 187050 287688 187056 287700
rect 169076 287660 187056 287688
rect 169076 287648 169082 287660
rect 187050 287648 187056 287660
rect 187108 287648 187114 287700
rect 93670 287104 93676 287156
rect 93728 287144 93734 287156
rect 102226 287144 102232 287156
rect 93728 287116 102232 287144
rect 93728 287104 93734 287116
rect 102226 287104 102232 287116
rect 102284 287104 102290 287156
rect 34514 287036 34520 287088
rect 34572 287076 34578 287088
rect 35710 287076 35716 287088
rect 34572 287048 35716 287076
rect 34572 287036 34578 287048
rect 35710 287036 35716 287048
rect 35768 287076 35774 287088
rect 70946 287076 70952 287088
rect 35768 287048 70952 287076
rect 35768 287036 35774 287048
rect 70946 287036 70952 287048
rect 71004 287036 71010 287088
rect 91462 287036 91468 287088
rect 91520 287076 91526 287088
rect 110506 287076 110512 287088
rect 91520 287048 110512 287076
rect 91520 287036 91526 287048
rect 110506 287036 110512 287048
rect 110564 287036 110570 287088
rect 82906 286968 82912 287020
rect 82964 287008 82970 287020
rect 85482 287008 85488 287020
rect 82964 286980 85488 287008
rect 82964 286968 82970 286980
rect 85482 286968 85488 286980
rect 85540 286968 85546 287020
rect 255498 286968 255504 287020
rect 255556 287008 255562 287020
rect 265066 287008 265072 287020
rect 255556 286980 265072 287008
rect 255556 286968 255562 286980
rect 265066 286968 265072 286980
rect 265124 286968 265130 287020
rect 74074 286900 74080 286952
rect 74132 286940 74138 286952
rect 76558 286940 76564 286952
rect 74132 286912 76564 286940
rect 74132 286900 74138 286912
rect 76558 286900 76564 286912
rect 76616 286900 76622 286952
rect 77386 286356 77392 286408
rect 77444 286396 77450 286408
rect 77938 286396 77944 286408
rect 77444 286368 77944 286396
rect 77444 286356 77450 286368
rect 77938 286356 77944 286368
rect 77996 286356 78002 286408
rect 3418 286288 3424 286340
rect 3476 286328 3482 286340
rect 15838 286328 15844 286340
rect 3476 286300 15844 286328
rect 3476 286288 3482 286300
rect 15838 286288 15844 286300
rect 15896 286288 15902 286340
rect 93026 286288 93032 286340
rect 93084 286328 93090 286340
rect 93762 286328 93768 286340
rect 93084 286300 93768 286328
rect 93084 286288 93090 286300
rect 93762 286288 93768 286300
rect 93820 286288 93826 286340
rect 45370 285812 45376 285864
rect 45428 285852 45434 285864
rect 75270 285852 75276 285864
rect 45428 285824 75276 285852
rect 45428 285812 45434 285824
rect 75270 285812 75276 285824
rect 75328 285812 75334 285864
rect 72510 285784 72516 285796
rect 64156 285756 72516 285784
rect 64156 285660 64184 285756
rect 72510 285744 72516 285756
rect 72568 285744 72574 285796
rect 148318 285744 148324 285796
rect 148376 285784 148382 285796
rect 165522 285784 165528 285796
rect 148376 285756 165528 285784
rect 148376 285744 148382 285756
rect 165522 285744 165528 285756
rect 165580 285784 165586 285796
rect 191742 285784 191748 285796
rect 165580 285756 191748 285784
rect 165580 285744 165586 285756
rect 191742 285744 191748 285756
rect 191800 285744 191806 285796
rect 95602 285676 95608 285728
rect 95660 285716 95666 285728
rect 107562 285716 107568 285728
rect 95660 285688 107568 285716
rect 95660 285676 95666 285688
rect 107562 285676 107568 285688
rect 107620 285676 107626 285728
rect 115842 285676 115848 285728
rect 115900 285716 115906 285728
rect 190362 285716 190368 285728
rect 115900 285688 190368 285716
rect 115900 285676 115906 285688
rect 190362 285676 190368 285688
rect 190420 285676 190426 285728
rect 63218 285608 63224 285660
rect 63276 285648 63282 285660
rect 64138 285648 64144 285660
rect 63276 285620 64144 285648
rect 63276 285608 63282 285620
rect 64138 285608 64144 285620
rect 64196 285608 64202 285660
rect 43898 284928 43904 284980
rect 43956 284968 43962 284980
rect 60734 284968 60740 284980
rect 43956 284940 60740 284968
rect 43956 284928 43962 284940
rect 60734 284928 60740 284940
rect 60792 284928 60798 284980
rect 67542 284928 67548 284980
rect 67600 284968 67606 284980
rect 68646 284968 68652 284980
rect 67600 284940 68652 284968
rect 67600 284928 67606 284940
rect 68646 284928 68652 284940
rect 68704 284968 68710 284980
rect 98362 284968 98368 284980
rect 68704 284940 98368 284968
rect 68704 284928 68710 284940
rect 98362 284928 98368 284940
rect 98420 284928 98426 284980
rect 151170 284928 151176 284980
rect 151228 284968 151234 284980
rect 178770 284968 178776 284980
rect 151228 284940 178776 284968
rect 151228 284928 151234 284940
rect 178770 284928 178776 284940
rect 178828 284928 178834 284980
rect 255590 284928 255596 284980
rect 255648 284968 255654 284980
rect 267734 284968 267740 284980
rect 255648 284940 267740 284968
rect 255648 284928 255654 284940
rect 267734 284928 267740 284940
rect 267792 284928 267798 284980
rect 255406 284520 255412 284572
rect 255464 284560 255470 284572
rect 259546 284560 259552 284572
rect 255464 284532 259552 284560
rect 255464 284520 255470 284532
rect 259546 284520 259552 284532
rect 259604 284520 259610 284572
rect 52086 284316 52092 284368
rect 52144 284356 52150 284368
rect 76650 284356 76656 284368
rect 52144 284328 76656 284356
rect 52144 284316 52150 284328
rect 76650 284316 76656 284328
rect 76708 284316 76714 284368
rect 173250 284316 173256 284368
rect 173308 284356 173314 284368
rect 191742 284356 191748 284368
rect 173308 284328 191748 284356
rect 173308 284316 173314 284328
rect 191742 284316 191748 284328
rect 191800 284316 191806 284368
rect 255406 284248 255412 284300
rect 255464 284288 255470 284300
rect 261018 284288 261024 284300
rect 255464 284260 261024 284288
rect 255464 284248 255470 284260
rect 261018 284248 261024 284260
rect 261076 284248 261082 284300
rect 75040 283704 75046 283756
rect 75098 283744 75104 283756
rect 75270 283744 75276 283756
rect 75098 283716 75276 283744
rect 75098 283704 75104 283716
rect 75270 283704 75276 283716
rect 75328 283704 75334 283756
rect 39942 283568 39948 283620
rect 40000 283608 40006 283620
rect 52454 283608 52460 283620
rect 40000 283580 52460 283608
rect 40000 283568 40006 283580
rect 52454 283568 52460 283580
rect 52512 283568 52518 283620
rect 91370 283568 91376 283620
rect 91428 283608 91434 283620
rect 93118 283608 93124 283620
rect 91428 283580 93124 283608
rect 91428 283568 91434 283580
rect 93118 283568 93124 283580
rect 93176 283608 93182 283620
rect 99466 283608 99472 283620
rect 93176 283580 99472 283608
rect 93176 283568 93182 283580
rect 99466 283568 99472 283580
rect 99524 283568 99530 283620
rect 97902 283432 97908 283484
rect 97960 283472 97966 283484
rect 98454 283472 98460 283484
rect 97960 283444 98460 283472
rect 97960 283432 97966 283444
rect 98454 283432 98460 283444
rect 98512 283432 98518 283484
rect 69106 283132 69112 283144
rect 60706 283104 69112 283132
rect 47854 282956 47860 283008
rect 47912 282996 47918 283008
rect 60706 282996 60734 283104
rect 69106 283092 69112 283104
rect 69164 283132 69170 283144
rect 69842 283132 69848 283144
rect 69164 283104 69848 283132
rect 69164 283092 69170 283104
rect 69842 283092 69848 283104
rect 69900 283092 69906 283144
rect 68646 283024 68652 283076
rect 68704 283064 68710 283076
rect 80238 283064 80244 283076
rect 68704 283036 80244 283064
rect 68704 283024 68710 283036
rect 80238 283024 80244 283036
rect 80296 283024 80302 283076
rect 47912 282968 60734 282996
rect 47912 282956 47918 282968
rect 68370 282956 68376 283008
rect 68428 282996 68434 283008
rect 69198 282996 69204 283008
rect 68428 282968 69204 282996
rect 68428 282956 68434 282968
rect 69198 282956 69204 282968
rect 69256 282956 69262 283008
rect 69750 282956 69756 283008
rect 69808 282996 69814 283008
rect 69808 282968 69888 282996
rect 69808 282956 69814 282968
rect 64506 282208 64512 282260
rect 64564 282248 64570 282260
rect 69860 282248 69888 282968
rect 84746 282956 84752 283008
rect 84804 282996 84810 283008
rect 84804 282968 89714 282996
rect 84804 282956 84810 282968
rect 89686 282928 89714 282968
rect 106366 282928 106372 282940
rect 89686 282900 106372 282928
rect 106366 282888 106372 282900
rect 106424 282888 106430 282940
rect 126238 282888 126244 282940
rect 126296 282928 126302 282940
rect 191742 282928 191748 282940
rect 126296 282900 191748 282928
rect 126296 282888 126302 282900
rect 191742 282888 191748 282900
rect 191800 282888 191806 282940
rect 98914 282820 98920 282872
rect 98972 282860 98978 282872
rect 99374 282860 99380 282872
rect 98972 282832 99380 282860
rect 98972 282820 98978 282832
rect 99374 282820 99380 282832
rect 99432 282820 99438 282872
rect 255498 282820 255504 282872
rect 255556 282860 255562 282872
rect 266630 282860 266636 282872
rect 255556 282832 266636 282860
rect 255556 282820 255562 282832
rect 266630 282820 266636 282832
rect 266688 282820 266694 282872
rect 255406 282752 255412 282804
rect 255464 282792 255470 282804
rect 258350 282792 258356 282804
rect 255464 282764 258356 282792
rect 255464 282752 255470 282764
rect 258350 282752 258356 282764
rect 258408 282752 258414 282804
rect 64564 282220 69888 282248
rect 64564 282208 64570 282220
rect 52454 282140 52460 282192
rect 52512 282180 52518 282192
rect 53650 282180 53656 282192
rect 52512 282152 53656 282180
rect 52512 282140 52518 282152
rect 53650 282140 53656 282152
rect 53708 282180 53714 282192
rect 69014 282180 69020 282192
rect 53708 282152 69020 282180
rect 53708 282140 53714 282152
rect 69014 282140 69020 282152
rect 69072 282180 69078 282192
rect 187142 282180 187148 282192
rect 69072 282152 187148 282180
rect 69072 282140 69078 282152
rect 187142 282140 187148 282152
rect 187200 282140 187206 282192
rect 120902 281528 120908 281580
rect 120960 281568 120966 281580
rect 128446 281568 128452 281580
rect 120960 281540 128452 281568
rect 120960 281528 120966 281540
rect 128446 281528 128452 281540
rect 128504 281528 128510 281580
rect 48130 281460 48136 281512
rect 48188 281500 48194 281512
rect 53098 281500 53104 281512
rect 48188 281472 53104 281500
rect 48188 281460 48194 281472
rect 53098 281460 53104 281472
rect 53156 281460 53162 281512
rect 98362 281460 98368 281512
rect 98420 281500 98426 281512
rect 189718 281500 189724 281512
rect 98420 281472 189724 281500
rect 98420 281460 98426 281472
rect 189718 281460 189724 281472
rect 189776 281460 189782 281512
rect 255406 281460 255412 281512
rect 255464 281500 255470 281512
rect 262490 281500 262496 281512
rect 255464 281472 262496 281500
rect 255464 281460 255470 281472
rect 262490 281460 262496 281472
rect 262548 281460 262554 281512
rect 99374 280780 99380 280832
rect 99432 280820 99438 280832
rect 113358 280820 113364 280832
rect 99432 280792 113364 280820
rect 99432 280780 99438 280792
rect 113358 280780 113364 280792
rect 113416 280820 113422 280832
rect 134610 280820 134616 280832
rect 113416 280792 134616 280820
rect 113416 280780 113422 280792
rect 134610 280780 134616 280792
rect 134668 280780 134674 280832
rect 3418 280168 3424 280220
rect 3476 280208 3482 280220
rect 67542 280208 67548 280220
rect 3476 280180 67548 280208
rect 3476 280168 3482 280180
rect 67542 280168 67548 280180
rect 67600 280168 67606 280220
rect 169110 280168 169116 280220
rect 169168 280208 169174 280220
rect 191558 280208 191564 280220
rect 169168 280180 191564 280208
rect 169168 280168 169174 280180
rect 191558 280168 191564 280180
rect 191616 280168 191622 280220
rect 255498 280168 255504 280220
rect 255556 280208 255562 280220
rect 271874 280208 271880 280220
rect 255556 280180 271880 280208
rect 255556 280168 255562 280180
rect 271874 280168 271880 280180
rect 271932 280168 271938 280220
rect 108942 280100 108948 280152
rect 109000 280140 109006 280152
rect 186958 280140 186964 280152
rect 109000 280112 186964 280140
rect 109000 280100 109006 280112
rect 186958 280100 186964 280112
rect 187016 280100 187022 280152
rect 255314 280100 255320 280152
rect 255372 280140 255378 280152
rect 263778 280140 263784 280152
rect 255372 280112 263784 280140
rect 255372 280100 255378 280112
rect 263778 280100 263784 280112
rect 263836 280100 263842 280152
rect 255406 280032 255412 280084
rect 255464 280072 255470 280084
rect 259730 280072 259736 280084
rect 255464 280044 259736 280072
rect 255464 280032 255470 280044
rect 259730 280032 259736 280044
rect 259788 280032 259794 280084
rect 57882 279556 57888 279608
rect 57940 279596 57946 279608
rect 66070 279596 66076 279608
rect 57940 279568 66076 279596
rect 57940 279556 57946 279568
rect 66070 279556 66076 279568
rect 66128 279596 66134 279608
rect 66622 279596 66628 279608
rect 66128 279568 66628 279596
rect 66128 279556 66134 279568
rect 66622 279556 66628 279568
rect 66680 279556 66686 279608
rect 191742 279528 191748 279540
rect 190426 279500 191748 279528
rect 4798 279420 4804 279472
rect 4856 279460 4862 279472
rect 32858 279460 32864 279472
rect 4856 279432 32864 279460
rect 4856 279420 4862 279432
rect 32858 279420 32864 279432
rect 32916 279460 32922 279472
rect 60366 279460 60372 279472
rect 32916 279432 60372 279460
rect 32916 279420 32922 279432
rect 60366 279420 60372 279432
rect 60424 279460 60430 279472
rect 66806 279460 66812 279472
rect 60424 279432 66812 279460
rect 60424 279420 60430 279432
rect 66806 279420 66812 279432
rect 66864 279420 66870 279472
rect 99466 279420 99472 279472
rect 99524 279460 99530 279472
rect 107838 279460 107844 279472
rect 99524 279432 107844 279460
rect 99524 279420 99530 279432
rect 107838 279420 107844 279432
rect 107896 279420 107902 279472
rect 175182 279420 175188 279472
rect 175240 279460 175246 279472
rect 187694 279460 187700 279472
rect 175240 279432 187700 279460
rect 175240 279420 175246 279432
rect 187694 279420 187700 279432
rect 187752 279460 187758 279472
rect 190426 279460 190454 279500
rect 191742 279488 191748 279500
rect 191800 279488 191806 279540
rect 187752 279432 190454 279460
rect 187752 279420 187758 279432
rect 108298 279216 108304 279268
rect 108356 279256 108362 279268
rect 108942 279256 108948 279268
rect 108356 279228 108948 279256
rect 108356 279216 108362 279228
rect 108942 279216 108948 279228
rect 109000 279216 109006 279268
rect 142982 278740 142988 278792
rect 143040 278780 143046 278792
rect 175182 278780 175188 278792
rect 143040 278752 175188 278780
rect 143040 278740 143046 278752
rect 175182 278740 175188 278752
rect 175240 278740 175246 278792
rect 128446 278672 128452 278724
rect 128504 278712 128510 278724
rect 191742 278712 191748 278724
rect 128504 278684 191748 278712
rect 128504 278672 128510 278684
rect 191742 278672 191748 278684
rect 191800 278672 191806 278724
rect 259362 278672 259368 278724
rect 259420 278712 259426 278724
rect 259822 278712 259828 278724
rect 259420 278684 259828 278712
rect 259420 278672 259426 278684
rect 259822 278672 259828 278684
rect 259880 278672 259886 278724
rect 255406 278468 255412 278520
rect 255464 278508 255470 278520
rect 258074 278508 258080 278520
rect 255464 278480 258080 278508
rect 255464 278468 255470 278480
rect 258074 278468 258080 278480
rect 258132 278468 258138 278520
rect 50982 277992 50988 278044
rect 51040 278032 51046 278044
rect 59170 278032 59176 278044
rect 51040 278004 59176 278032
rect 51040 277992 51046 278004
rect 59170 277992 59176 278004
rect 59228 278032 59234 278044
rect 66806 278032 66812 278044
rect 59228 278004 66812 278032
rect 59228 277992 59234 278004
rect 66806 277992 66812 278004
rect 66864 277992 66870 278044
rect 102042 277992 102048 278044
rect 102100 278032 102106 278044
rect 131206 278032 131212 278044
rect 102100 278004 131212 278032
rect 102100 277992 102106 278004
rect 131206 277992 131212 278004
rect 131264 278032 131270 278044
rect 151078 278032 151084 278044
rect 131264 278004 151084 278032
rect 131264 277992 131270 278004
rect 151078 277992 151084 278004
rect 151136 277992 151142 278044
rect 255406 277448 255412 277500
rect 255464 277488 255470 277500
rect 258166 277488 258172 277500
rect 255464 277460 258172 277488
rect 255464 277448 255470 277460
rect 258166 277448 258172 277460
rect 258224 277448 258230 277500
rect 162210 277380 162216 277432
rect 162268 277420 162274 277432
rect 191650 277420 191656 277432
rect 162268 277392 191656 277420
rect 162268 277380 162274 277392
rect 191650 277380 191656 277392
rect 191708 277380 191714 277432
rect 66070 277312 66076 277364
rect 66128 277352 66134 277364
rect 68278 277352 68284 277364
rect 66128 277324 68284 277352
rect 66128 277312 66134 277324
rect 68278 277312 68284 277324
rect 68336 277312 68342 277364
rect 113818 276700 113824 276752
rect 113876 276740 113882 276752
rect 127158 276740 127164 276752
rect 113876 276712 127164 276740
rect 113876 276700 113882 276712
rect 127158 276700 127164 276712
rect 127216 276700 127222 276752
rect 100018 276632 100024 276684
rect 100076 276672 100082 276684
rect 118970 276672 118976 276684
rect 100076 276644 118976 276672
rect 100076 276632 100082 276644
rect 118970 276632 118976 276644
rect 119028 276632 119034 276684
rect 144822 276632 144828 276684
rect 144880 276672 144886 276684
rect 182818 276672 182824 276684
rect 144880 276644 182824 276672
rect 144880 276632 144886 276644
rect 182818 276632 182824 276644
rect 182876 276632 182882 276684
rect 102134 276292 102140 276344
rect 102192 276332 102198 276344
rect 102778 276332 102784 276344
rect 102192 276304 102784 276332
rect 102192 276292 102198 276304
rect 102778 276292 102784 276304
rect 102836 276292 102842 276344
rect 255498 276088 255504 276140
rect 255556 276128 255562 276140
rect 263594 276128 263600 276140
rect 255556 276100 263600 276128
rect 255556 276088 255562 276100
rect 263594 276088 263600 276100
rect 263652 276088 263658 276140
rect 43898 276020 43904 276072
rect 43956 276060 43962 276072
rect 52454 276060 52460 276072
rect 43956 276032 52460 276060
rect 43956 276020 43962 276032
rect 52454 276020 52460 276032
rect 52512 276060 52518 276072
rect 66806 276060 66812 276072
rect 52512 276032 66812 276060
rect 52512 276020 52518 276032
rect 66806 276020 66812 276032
rect 66864 276020 66870 276072
rect 136542 276020 136548 276072
rect 136600 276060 136606 276072
rect 144178 276060 144184 276072
rect 136600 276032 144184 276060
rect 136600 276020 136606 276032
rect 144178 276020 144184 276032
rect 144236 276020 144242 276072
rect 255314 276020 255320 276072
rect 255372 276060 255378 276072
rect 265250 276060 265256 276072
rect 255372 276032 265256 276060
rect 255372 276020 255378 276032
rect 265250 276020 265256 276032
rect 265308 276020 265314 276072
rect 63402 275952 63408 276004
rect 63460 275992 63466 276004
rect 66898 275992 66904 276004
rect 63460 275964 66904 275992
rect 63460 275952 63466 275964
rect 66898 275952 66904 275964
rect 66956 275952 66962 276004
rect 255406 275952 255412 276004
rect 255464 275992 255470 276004
rect 264974 275992 264980 276004
rect 255464 275964 264980 275992
rect 255464 275952 255470 275964
rect 264974 275952 264980 275964
rect 265032 275952 265038 276004
rect 261478 275340 261484 275392
rect 261536 275380 261542 275392
rect 269114 275380 269120 275392
rect 261536 275352 269120 275380
rect 261536 275340 261542 275352
rect 269114 275340 269120 275352
rect 269172 275340 269178 275392
rect 100754 275272 100760 275324
rect 100812 275312 100818 275324
rect 142154 275312 142160 275324
rect 100812 275284 142160 275312
rect 100812 275272 100818 275284
rect 142154 275272 142160 275284
rect 142212 275312 142218 275324
rect 142890 275312 142896 275324
rect 142212 275284 142896 275312
rect 142212 275272 142218 275284
rect 142890 275272 142896 275284
rect 142948 275272 142954 275324
rect 155218 275272 155224 275324
rect 155276 275312 155282 275324
rect 188338 275312 188344 275324
rect 155276 275284 188344 275312
rect 155276 275272 155282 275284
rect 188338 275272 188344 275284
rect 188396 275272 188402 275324
rect 188982 274728 188988 274780
rect 189040 274768 189046 274780
rect 191650 274768 191656 274780
rect 189040 274740 191656 274768
rect 189040 274728 189046 274740
rect 191650 274728 191656 274740
rect 191708 274728 191714 274780
rect 57790 274660 57796 274712
rect 57848 274700 57854 274712
rect 63402 274700 63408 274712
rect 57848 274672 63408 274700
rect 57848 274660 57854 274672
rect 63402 274660 63408 274672
rect 63460 274660 63466 274712
rect 130562 274660 130568 274712
rect 130620 274700 130626 274712
rect 168282 274700 168288 274712
rect 130620 274672 168288 274700
rect 130620 274660 130626 274672
rect 168282 274660 168288 274672
rect 168340 274700 168346 274712
rect 191742 274700 191748 274712
rect 168340 274672 191748 274700
rect 168340 274660 168346 274672
rect 191742 274660 191748 274672
rect 191800 274660 191806 274712
rect 58894 274592 58900 274644
rect 58952 274632 58958 274644
rect 65886 274632 65892 274644
rect 58952 274604 65892 274632
rect 58952 274592 58958 274604
rect 65886 274592 65892 274604
rect 65944 274632 65950 274644
rect 66530 274632 66536 274644
rect 65944 274604 66536 274632
rect 65944 274592 65950 274604
rect 66530 274592 66536 274604
rect 66588 274592 66594 274644
rect 141418 274592 141424 274644
rect 141476 274632 141482 274644
rect 193122 274632 193128 274644
rect 141476 274604 193128 274632
rect 141476 274592 141482 274604
rect 193122 274592 193128 274604
rect 193180 274592 193186 274644
rect 255406 274592 255412 274644
rect 255464 274632 255470 274644
rect 260834 274632 260840 274644
rect 255464 274604 260840 274632
rect 255464 274592 255470 274604
rect 260834 274592 260840 274604
rect 260892 274592 260898 274644
rect 58894 274116 58900 274168
rect 58952 274156 58958 274168
rect 59262 274156 59268 274168
rect 58952 274128 59268 274156
rect 58952 274116 58958 274128
rect 59262 274116 59268 274128
rect 59320 274116 59326 274168
rect 100754 273980 100760 274032
rect 100812 274020 100818 274032
rect 128446 274020 128452 274032
rect 100812 273992 128452 274020
rect 100812 273980 100818 273992
rect 128446 273980 128452 273992
rect 128504 273980 128510 274032
rect 100846 273912 100852 273964
rect 100904 273952 100910 273964
rect 135254 273952 135260 273964
rect 100904 273924 135260 273952
rect 100904 273912 100910 273924
rect 135254 273912 135260 273924
rect 135312 273952 135318 273964
rect 136542 273952 136548 273964
rect 135312 273924 136548 273952
rect 135312 273912 135318 273924
rect 136542 273912 136548 273924
rect 136600 273912 136606 273964
rect 255958 273912 255964 273964
rect 256016 273952 256022 273964
rect 582466 273952 582472 273964
rect 256016 273924 582472 273952
rect 256016 273912 256022 273924
rect 582466 273912 582472 273924
rect 582524 273912 582530 273964
rect 128446 273844 128452 273896
rect 128504 273884 128510 273896
rect 128998 273884 129004 273896
rect 128504 273856 129004 273884
rect 128504 273844 128510 273856
rect 128998 273844 129004 273856
rect 129056 273844 129062 273896
rect 104158 273164 104164 273216
rect 104216 273204 104222 273216
rect 116854 273204 116860 273216
rect 104216 273176 116860 273204
rect 104216 273164 104222 273176
rect 116854 273164 116860 273176
rect 116912 273164 116918 273216
rect 116854 272484 116860 272536
rect 116912 272524 116918 272536
rect 169110 272524 169116 272536
rect 116912 272496 169116 272524
rect 116912 272484 116918 272496
rect 169110 272484 169116 272496
rect 169168 272484 169174 272536
rect 62850 272076 62856 272128
rect 62908 272116 62914 272128
rect 63218 272116 63224 272128
rect 62908 272088 63224 272116
rect 62908 272076 62914 272088
rect 63218 272076 63224 272088
rect 63276 272116 63282 272128
rect 66806 272116 66812 272128
rect 63276 272088 66812 272116
rect 63276 272076 63282 272088
rect 66806 272076 66812 272088
rect 66864 272076 66870 272128
rect 171778 271940 171784 271992
rect 171836 271980 171842 271992
rect 191190 271980 191196 271992
rect 171836 271952 191196 271980
rect 171836 271940 171842 271952
rect 191190 271940 191196 271952
rect 191248 271940 191254 271992
rect 255498 271940 255504 271992
rect 255556 271980 255562 271992
rect 269206 271980 269212 271992
rect 255556 271952 269212 271980
rect 255556 271940 255562 271952
rect 269206 271940 269212 271952
rect 269264 271940 269270 271992
rect 109678 271872 109684 271924
rect 109736 271912 109742 271924
rect 112254 271912 112260 271924
rect 109736 271884 112260 271912
rect 109736 271872 109742 271884
rect 112254 271872 112260 271884
rect 112312 271912 112318 271924
rect 122834 271912 122840 271924
rect 112312 271884 122840 271912
rect 112312 271872 112318 271884
rect 122834 271872 122840 271884
rect 122892 271912 122898 271924
rect 160922 271912 160928 271924
rect 122892 271884 160928 271912
rect 122892 271872 122898 271884
rect 160922 271872 160928 271884
rect 160980 271872 160986 271924
rect 163590 271872 163596 271924
rect 163648 271912 163654 271924
rect 191742 271912 191748 271924
rect 163648 271884 191748 271912
rect 163648 271872 163654 271884
rect 191742 271872 191748 271884
rect 191800 271872 191806 271924
rect 255406 271872 255412 271924
rect 255464 271912 255470 271924
rect 265066 271912 265072 271924
rect 255464 271884 265072 271912
rect 255464 271872 255470 271884
rect 265066 271872 265072 271884
rect 265124 271872 265130 271924
rect 266998 271872 267004 271924
rect 267056 271912 267062 271924
rect 580166 271912 580172 271924
rect 267056 271884 580172 271912
rect 267056 271872 267062 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 54938 271804 54944 271856
rect 54996 271844 55002 271856
rect 56410 271844 56416 271856
rect 54996 271816 56416 271844
rect 54996 271804 55002 271816
rect 56410 271804 56416 271816
rect 56468 271844 56474 271856
rect 66806 271844 66812 271856
rect 56468 271816 66812 271844
rect 56468 271804 56474 271816
rect 66806 271804 66812 271816
rect 66864 271804 66870 271856
rect 255314 271804 255320 271856
rect 255372 271844 255378 271856
rect 266538 271844 266544 271856
rect 255372 271816 266544 271844
rect 255372 271804 255378 271816
rect 266538 271804 266544 271816
rect 266596 271804 266602 271856
rect 255498 271600 255504 271652
rect 255556 271640 255562 271652
rect 259454 271640 259460 271652
rect 255556 271612 259460 271640
rect 255556 271600 255562 271612
rect 259454 271600 259460 271612
rect 259512 271600 259518 271652
rect 101674 271124 101680 271176
rect 101732 271164 101738 271176
rect 103422 271164 103428 271176
rect 101732 271136 103428 271164
rect 101732 271124 101738 271136
rect 103422 271124 103428 271136
rect 103480 271164 103486 271176
rect 130378 271164 130384 271176
rect 103480 271136 130384 271164
rect 103480 271124 103486 271136
rect 130378 271124 130384 271136
rect 130436 271164 130442 271176
rect 173158 271164 173164 271176
rect 130436 271136 173164 271164
rect 130436 271124 130442 271136
rect 173158 271124 173164 271136
rect 173216 271124 173222 271176
rect 100754 269900 100760 269952
rect 100812 269940 100818 269952
rect 104434 269940 104440 269952
rect 100812 269912 104440 269940
rect 100812 269900 100818 269912
rect 104434 269900 104440 269912
rect 104492 269900 104498 269952
rect 135898 269764 135904 269816
rect 135956 269804 135962 269816
rect 188430 269804 188436 269816
rect 135956 269776 188436 269804
rect 135956 269764 135962 269776
rect 188430 269764 188436 269776
rect 188488 269764 188494 269816
rect 255590 269764 255596 269816
rect 255648 269804 255654 269816
rect 273346 269804 273352 269816
rect 255648 269776 273352 269804
rect 255648 269764 255654 269776
rect 273346 269764 273352 269776
rect 273404 269764 273410 269816
rect 103974 269084 103980 269136
rect 104032 269124 104038 269136
rect 106826 269124 106832 269136
rect 104032 269096 106832 269124
rect 104032 269084 104038 269096
rect 106826 269084 106832 269096
rect 106884 269124 106890 269136
rect 135898 269124 135904 269136
rect 106884 269096 135904 269124
rect 106884 269084 106890 269096
rect 135898 269084 135904 269096
rect 135956 269084 135962 269136
rect 181438 269084 181444 269136
rect 181496 269124 181502 269136
rect 191742 269124 191748 269136
rect 181496 269096 191748 269124
rect 181496 269084 181502 269096
rect 191742 269084 191748 269096
rect 191800 269084 191806 269136
rect 255406 269084 255412 269136
rect 255464 269124 255470 269136
rect 260926 269124 260932 269136
rect 255464 269096 260932 269124
rect 255464 269084 255470 269096
rect 260926 269084 260932 269096
rect 260984 269084 260990 269136
rect 104894 269016 104900 269068
rect 104952 269056 104958 269068
rect 109586 269056 109592 269068
rect 104952 269028 109592 269056
rect 104952 269016 104958 269028
rect 109586 269016 109592 269028
rect 109644 269016 109650 269068
rect 131758 269016 131764 269068
rect 131816 269056 131822 269068
rect 192478 269056 192484 269068
rect 131816 269028 192484 269056
rect 131816 269016 131822 269028
rect 192478 269016 192484 269028
rect 192536 269016 192542 269068
rect 116670 268880 116676 268932
rect 116728 268920 116734 268932
rect 118878 268920 118884 268932
rect 116728 268892 118884 268920
rect 116728 268880 116734 268892
rect 118878 268880 118884 268892
rect 118936 268880 118942 268932
rect 100754 268404 100760 268456
rect 100812 268444 100818 268456
rect 104894 268444 104900 268456
rect 100812 268416 104900 268444
rect 100812 268404 100818 268416
rect 104894 268404 104900 268416
rect 104952 268404 104958 268456
rect 52362 268336 52368 268388
rect 52420 268376 52426 268388
rect 66162 268376 66168 268388
rect 52420 268348 66168 268376
rect 52420 268336 52426 268348
rect 66162 268336 66168 268348
rect 66220 268336 66226 268388
rect 100846 268336 100852 268388
rect 100904 268376 100910 268388
rect 113266 268376 113272 268388
rect 100904 268348 113272 268376
rect 100904 268336 100910 268348
rect 113266 268336 113272 268348
rect 113324 268376 113330 268388
rect 113910 268376 113916 268388
rect 113324 268348 113916 268376
rect 113324 268336 113330 268348
rect 113910 268336 113916 268348
rect 113968 268336 113974 268388
rect 178770 267724 178776 267776
rect 178828 267764 178834 267776
rect 191650 267764 191656 267776
rect 178828 267736 191656 267764
rect 178828 267724 178834 267736
rect 191650 267724 191656 267736
rect 191708 267724 191714 267776
rect 255498 267724 255504 267776
rect 255556 267764 255562 267776
rect 261110 267764 261116 267776
rect 255556 267736 261116 267764
rect 255556 267724 255562 267736
rect 261110 267724 261116 267736
rect 261168 267724 261174 267776
rect 53742 267656 53748 267708
rect 53800 267696 53806 267708
rect 66254 267696 66260 267708
rect 53800 267668 66260 267696
rect 53800 267656 53806 267668
rect 66254 267656 66260 267668
rect 66312 267656 66318 267708
rect 255406 267656 255412 267708
rect 255464 267696 255470 267708
rect 285674 267696 285680 267708
rect 255464 267668 285680 267696
rect 255464 267656 255470 267668
rect 285674 267656 285680 267668
rect 285732 267656 285738 267708
rect 104434 266976 104440 267028
rect 104492 267016 104498 267028
rect 119430 267016 119436 267028
rect 104492 266988 119436 267016
rect 104492 266976 104498 266988
rect 119430 266976 119436 266988
rect 119488 266976 119494 267028
rect 141510 266976 141516 267028
rect 141568 267016 141574 267028
rect 180150 267016 180156 267028
rect 141568 266988 180156 267016
rect 141568 266976 141574 266988
rect 180150 266976 180156 266988
rect 180208 266976 180214 267028
rect 255406 266976 255412 267028
rect 255464 267016 255470 267028
rect 262214 267016 262220 267028
rect 255464 266988 262220 267016
rect 255464 266976 255470 266988
rect 262214 266976 262220 266988
rect 262272 266976 262278 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 11698 266404 11704 266416
rect 3108 266376 11704 266404
rect 3108 266364 3114 266376
rect 11698 266364 11704 266376
rect 11756 266364 11762 266416
rect 66806 266404 66812 266416
rect 50356 266376 66812 266404
rect 50356 266348 50384 266376
rect 66806 266364 66812 266376
rect 66864 266364 66870 266416
rect 115382 266364 115388 266416
rect 115440 266404 115446 266416
rect 120902 266404 120908 266416
rect 115440 266376 120908 266404
rect 115440 266364 115446 266376
rect 120902 266364 120908 266376
rect 120960 266364 120966 266416
rect 177390 266364 177396 266416
rect 177448 266404 177454 266416
rect 191466 266404 191472 266416
rect 177448 266376 191472 266404
rect 177448 266364 177454 266376
rect 191466 266364 191472 266376
rect 191524 266364 191530 266416
rect 37182 266296 37188 266348
rect 37240 266336 37246 266348
rect 50338 266336 50344 266348
rect 37240 266308 50344 266336
rect 37240 266296 37246 266308
rect 50338 266296 50344 266308
rect 50396 266296 50402 266348
rect 149054 266296 149060 266348
rect 149112 266336 149118 266348
rect 162210 266336 162216 266348
rect 149112 266308 162216 266336
rect 149112 266296 149118 266308
rect 162210 266296 162216 266308
rect 162268 266296 162274 266348
rect 255314 266296 255320 266348
rect 255372 266336 255378 266348
rect 276014 266336 276020 266348
rect 255372 266308 276020 266336
rect 255372 266296 255378 266308
rect 276014 266296 276020 266308
rect 276072 266296 276078 266348
rect 100110 265616 100116 265668
rect 100168 265656 100174 265668
rect 107654 265656 107660 265668
rect 100168 265628 107660 265656
rect 100168 265616 100174 265628
rect 107654 265616 107660 265628
rect 107712 265616 107718 265668
rect 133782 265616 133788 265668
rect 133840 265656 133846 265668
rect 149054 265656 149060 265668
rect 133840 265628 149060 265656
rect 133840 265616 133846 265628
rect 149054 265616 149060 265628
rect 149112 265616 149118 265668
rect 159450 265616 159456 265668
rect 159508 265656 159514 265668
rect 185578 265656 185584 265668
rect 159508 265628 185584 265656
rect 159508 265616 159514 265628
rect 185578 265616 185584 265628
rect 185636 265616 185642 265668
rect 255958 265616 255964 265668
rect 256016 265656 256022 265668
rect 583202 265656 583208 265668
rect 256016 265628 583208 265656
rect 256016 265616 256022 265628
rect 583202 265616 583208 265628
rect 583260 265616 583266 265668
rect 60642 265140 60648 265192
rect 60700 265180 60706 265192
rect 66806 265180 66812 265192
rect 60700 265152 66812 265180
rect 60700 265140 60706 265152
rect 66806 265140 66812 265152
rect 66864 265140 66870 265192
rect 100846 264936 100852 264988
rect 100904 264976 100910 264988
rect 133138 264976 133144 264988
rect 100904 264948 133144 264976
rect 100904 264936 100910 264948
rect 133138 264936 133144 264948
rect 133196 264976 133202 264988
rect 133782 264976 133788 264988
rect 133196 264948 133788 264976
rect 133196 264936 133202 264948
rect 133782 264936 133788 264948
rect 133840 264936 133846 264988
rect 182818 264936 182824 264988
rect 182876 264976 182882 264988
rect 191742 264976 191748 264988
rect 182876 264948 191748 264976
rect 182876 264936 182882 264948
rect 191742 264936 191748 264948
rect 191800 264936 191806 264988
rect 41138 264188 41144 264240
rect 41196 264228 41202 264240
rect 66622 264228 66628 264240
rect 41196 264200 66628 264228
rect 41196 264188 41202 264200
rect 66622 264188 66628 264200
rect 66680 264188 66686 264240
rect 100754 264188 100760 264240
rect 100812 264228 100818 264240
rect 127066 264228 127072 264240
rect 100812 264200 127072 264228
rect 100812 264188 100818 264200
rect 127066 264188 127072 264200
rect 127124 264188 127130 264240
rect 255406 263644 255412 263696
rect 255464 263684 255470 263696
rect 262214 263684 262220 263696
rect 255464 263656 262220 263684
rect 255464 263644 255470 263656
rect 262214 263644 262220 263656
rect 262272 263644 262278 263696
rect 36538 263576 36544 263628
rect 36596 263616 36602 263628
rect 41138 263616 41144 263628
rect 36596 263588 41144 263616
rect 36596 263576 36602 263588
rect 41138 263576 41144 263588
rect 41196 263576 41202 263628
rect 100754 263576 100760 263628
rect 100812 263616 100818 263628
rect 120074 263616 120080 263628
rect 100812 263588 120080 263616
rect 100812 263576 100818 263588
rect 120074 263576 120080 263588
rect 120132 263616 120138 263628
rect 147582 263616 147588 263628
rect 120132 263588 147588 263616
rect 120132 263576 120138 263588
rect 147582 263576 147588 263588
rect 147640 263576 147646 263628
rect 155310 263576 155316 263628
rect 155368 263616 155374 263628
rect 191006 263616 191012 263628
rect 155368 263588 191012 263616
rect 155368 263576 155374 263588
rect 191006 263576 191012 263588
rect 191064 263576 191070 263628
rect 115014 263508 115020 263560
rect 115072 263548 115078 263560
rect 118786 263548 118792 263560
rect 115072 263520 118792 263548
rect 115072 263508 115078 263520
rect 118786 263508 118792 263520
rect 118844 263548 118850 263560
rect 148318 263548 148324 263560
rect 118844 263520 148324 263548
rect 118844 263508 118850 263520
rect 148318 263508 148324 263520
rect 148376 263508 148382 263560
rect 255406 263508 255412 263560
rect 255464 263548 255470 263560
rect 262306 263548 262312 263560
rect 255464 263520 262312 263548
rect 255464 263508 255470 263520
rect 262306 263508 262312 263520
rect 262364 263508 262370 263560
rect 100754 262896 100760 262948
rect 100812 262936 100818 262948
rect 115014 262936 115020 262948
rect 100812 262908 115020 262936
rect 100812 262896 100818 262908
rect 115014 262896 115020 262908
rect 115072 262896 115078 262948
rect 33962 262828 33968 262880
rect 34020 262868 34026 262880
rect 60734 262868 60740 262880
rect 34020 262840 60740 262868
rect 34020 262828 34026 262840
rect 60734 262828 60740 262840
rect 60792 262868 60798 262880
rect 66898 262868 66904 262880
rect 60792 262840 66904 262868
rect 60792 262828 60798 262840
rect 66898 262828 66904 262840
rect 66956 262828 66962 262880
rect 104158 262828 104164 262880
rect 104216 262868 104222 262880
rect 124398 262868 124404 262880
rect 104216 262840 124404 262868
rect 104216 262828 104222 262840
rect 124398 262828 124404 262840
rect 124456 262828 124462 262880
rect 147582 262828 147588 262880
rect 147640 262868 147646 262880
rect 174538 262868 174544 262880
rect 147640 262840 174544 262868
rect 147640 262828 147646 262840
rect 174538 262828 174544 262840
rect 174596 262828 174602 262880
rect 268378 262828 268384 262880
rect 268436 262868 268442 262880
rect 580258 262868 580264 262880
rect 268436 262840 580264 262868
rect 268436 262828 268442 262840
rect 580258 262828 580264 262840
rect 580316 262828 580322 262880
rect 4798 262216 4804 262268
rect 4856 262256 4862 262268
rect 33962 262256 33968 262268
rect 4856 262228 33968 262256
rect 4856 262216 4862 262228
rect 33962 262216 33968 262228
rect 34020 262256 34026 262268
rect 34330 262256 34336 262268
rect 34020 262228 34336 262256
rect 34020 262216 34026 262228
rect 34330 262216 34336 262228
rect 34388 262216 34394 262268
rect 185578 262216 185584 262268
rect 185636 262256 185642 262268
rect 191006 262256 191012 262268
rect 185636 262228 191012 262256
rect 185636 262216 185642 262228
rect 191006 262216 191012 262228
rect 191064 262216 191070 262268
rect 63126 261536 63132 261588
rect 63184 261576 63190 261588
rect 68278 261576 68284 261588
rect 63184 261548 68284 261576
rect 63184 261536 63190 261548
rect 68278 261536 68284 261548
rect 68336 261536 68342 261588
rect 56410 261468 56416 261520
rect 56468 261508 56474 261520
rect 66714 261508 66720 261520
rect 56468 261480 66720 261508
rect 56468 261468 56474 261480
rect 66714 261468 66720 261480
rect 66772 261468 66778 261520
rect 100754 261468 100760 261520
rect 100812 261508 100818 261520
rect 104802 261508 104808 261520
rect 100812 261480 104808 261508
rect 100812 261468 100818 261480
rect 104802 261468 104808 261480
rect 104860 261508 104866 261520
rect 109218 261508 109224 261520
rect 104860 261480 109224 261508
rect 104860 261468 104866 261480
rect 109218 261468 109224 261480
rect 109276 261508 109282 261520
rect 134518 261508 134524 261520
rect 109276 261480 134524 261508
rect 109276 261468 109282 261480
rect 134518 261468 134524 261480
rect 134576 261468 134582 261520
rect 268470 261468 268476 261520
rect 268528 261508 268534 261520
rect 302234 261508 302240 261520
rect 268528 261480 302240 261508
rect 268528 261468 268534 261480
rect 302234 261468 302240 261480
rect 302292 261468 302298 261520
rect 104250 261060 104256 261112
rect 104308 261100 104314 261112
rect 108298 261100 108304 261112
rect 104308 261072 108304 261100
rect 104308 261060 104314 261072
rect 108298 261060 108304 261072
rect 108356 261060 108362 261112
rect 49510 260788 49516 260840
rect 49568 260828 49574 260840
rect 66438 260828 66444 260840
rect 49568 260800 66444 260828
rect 49568 260788 49574 260800
rect 66438 260788 66444 260800
rect 66496 260788 66502 260840
rect 113174 260720 113180 260772
rect 113232 260760 113238 260772
rect 115198 260760 115204 260772
rect 113232 260732 115204 260760
rect 113232 260720 113238 260732
rect 115198 260720 115204 260732
rect 115256 260720 115262 260772
rect 45462 260108 45468 260160
rect 45520 260148 45526 260160
rect 49510 260148 49516 260160
rect 45520 260120 49516 260148
rect 45520 260108 45526 260120
rect 49510 260108 49516 260120
rect 49568 260108 49574 260160
rect 135162 260108 135168 260160
rect 135220 260148 135226 260160
rect 144914 260148 144920 260160
rect 135220 260120 144920 260148
rect 135220 260108 135226 260120
rect 144914 260108 144920 260120
rect 144972 260148 144978 260160
rect 182910 260148 182916 260160
rect 144972 260120 182916 260148
rect 144972 260108 144978 260120
rect 182910 260108 182916 260120
rect 182968 260108 182974 260160
rect 271782 260108 271788 260160
rect 271840 260148 271846 260160
rect 582742 260148 582748 260160
rect 271840 260120 582748 260148
rect 271840 260108 271846 260120
rect 582742 260108 582748 260120
rect 582800 260108 582806 260160
rect 100846 259428 100852 259480
rect 100904 259468 100910 259480
rect 133966 259468 133972 259480
rect 100904 259440 133972 259468
rect 100904 259428 100910 259440
rect 133966 259428 133972 259440
rect 134024 259468 134030 259480
rect 135162 259468 135168 259480
rect 134024 259440 135168 259468
rect 134024 259428 134030 259440
rect 135162 259428 135168 259440
rect 135220 259428 135226 259480
rect 188246 259428 188252 259480
rect 188304 259468 188310 259480
rect 191742 259468 191748 259480
rect 188304 259440 191748 259468
rect 188304 259428 188310 259440
rect 191742 259428 191748 259440
rect 191800 259428 191806 259480
rect 255406 259428 255412 259480
rect 255464 259468 255470 259480
rect 260834 259468 260840 259480
rect 255464 259440 260840 259468
rect 255464 259428 255470 259440
rect 260834 259428 260840 259440
rect 260892 259428 260898 259480
rect 100754 258748 100760 258800
rect 100812 258788 100818 258800
rect 136726 258788 136732 258800
rect 100812 258760 136732 258788
rect 100812 258748 100818 258760
rect 136726 258748 136732 258760
rect 136784 258748 136790 258800
rect 266630 258748 266636 258800
rect 266688 258788 266694 258800
rect 307018 258788 307024 258800
rect 266688 258760 307024 258788
rect 266688 258748 266694 258760
rect 307018 258748 307024 258760
rect 307076 258748 307082 258800
rect 100846 258680 100852 258732
rect 100904 258720 100910 258732
rect 118050 258720 118056 258732
rect 100904 258692 118056 258720
rect 100904 258680 100910 258692
rect 118050 258680 118056 258692
rect 118108 258680 118114 258732
rect 133782 258680 133788 258732
rect 133840 258720 133846 258732
rect 173342 258720 173348 258732
rect 133840 258692 173348 258720
rect 133840 258680 133846 258692
rect 173342 258680 173348 258692
rect 173400 258680 173406 258732
rect 267918 258680 267924 258732
rect 267976 258720 267982 258732
rect 583294 258720 583300 258732
rect 267976 258692 583300 258720
rect 267976 258680 267982 258692
rect 583294 258680 583300 258692
rect 583352 258680 583358 258732
rect 45554 258136 45560 258188
rect 45612 258176 45618 258188
rect 46198 258176 46204 258188
rect 45612 258148 46204 258176
rect 45612 258136 45618 258148
rect 46198 258136 46204 258148
rect 46256 258176 46262 258188
rect 66254 258176 66260 258188
rect 46256 258148 66260 258176
rect 46256 258136 46262 258148
rect 66254 258136 66260 258148
rect 66312 258136 66318 258188
rect 100846 258176 100852 258188
rect 100772 258148 100852 258176
rect 100772 258120 100800 258148
rect 100846 258136 100852 258148
rect 100904 258136 100910 258188
rect 177298 258136 177304 258188
rect 177356 258176 177362 258188
rect 190638 258176 190644 258188
rect 177356 258148 190644 258176
rect 177356 258136 177362 258148
rect 190638 258136 190644 258148
rect 190696 258136 190702 258188
rect 42702 258068 42708 258120
rect 42760 258108 42766 258120
rect 66346 258108 66352 258120
rect 42760 258080 66352 258108
rect 42760 258068 42766 258080
rect 66346 258068 66352 258080
rect 66404 258068 66410 258120
rect 100754 258068 100760 258120
rect 100812 258068 100818 258120
rect 175918 258068 175924 258120
rect 175976 258108 175982 258120
rect 190546 258108 190552 258120
rect 175976 258080 190552 258108
rect 175976 258068 175982 258080
rect 190546 258068 190552 258080
rect 190604 258068 190610 258120
rect 255406 258068 255412 258120
rect 255464 258108 255470 258120
rect 266630 258108 266636 258120
rect 255464 258080 266636 258108
rect 255464 258068 255470 258080
rect 266630 258068 266636 258080
rect 266688 258068 266694 258120
rect 33042 258000 33048 258052
rect 33100 258040 33106 258052
rect 45554 258040 45560 258052
rect 33100 258012 45560 258040
rect 33100 258000 33106 258012
rect 45554 258000 45560 258012
rect 45612 258000 45618 258052
rect 66254 258000 66260 258052
rect 66312 258040 66318 258052
rect 68186 258040 68192 258052
rect 66312 258012 68192 258040
rect 66312 258000 66318 258012
rect 68186 258000 68192 258012
rect 68244 258000 68250 258052
rect 100846 258000 100852 258052
rect 100904 258040 100910 258052
rect 125502 258040 125508 258052
rect 100904 258012 125508 258040
rect 100904 258000 100910 258012
rect 125502 258000 125508 258012
rect 125560 258000 125566 258052
rect 190454 258000 190460 258052
rect 190512 258040 190518 258052
rect 193398 258040 193404 258052
rect 190512 258012 193404 258040
rect 190512 258000 190518 258012
rect 193398 258000 193404 258012
rect 193456 258000 193462 258052
rect 262674 258000 262680 258052
rect 262732 258040 262738 258052
rect 304258 258040 304264 258052
rect 262732 258012 304264 258040
rect 262732 258000 262738 258012
rect 304258 258000 304264 258012
rect 304316 258000 304322 258052
rect 255406 257388 255412 257440
rect 255464 257428 255470 257440
rect 262674 257428 262680 257440
rect 255464 257400 262680 257428
rect 255464 257388 255470 257400
rect 262674 257388 262680 257400
rect 262732 257388 262738 257440
rect 52270 257320 52276 257372
rect 52328 257360 52334 257372
rect 66622 257360 66628 257372
rect 52328 257332 66628 257360
rect 52328 257320 52334 257332
rect 66622 257320 66628 257332
rect 66680 257320 66686 257372
rect 110414 257320 110420 257372
rect 110472 257360 110478 257372
rect 130470 257360 130476 257372
rect 110472 257332 130476 257360
rect 110472 257320 110478 257332
rect 130470 257320 130476 257332
rect 130528 257320 130534 257372
rect 146938 257320 146944 257372
rect 146996 257360 147002 257372
rect 176010 257360 176016 257372
rect 146996 257332 176016 257360
rect 146996 257320 147002 257332
rect 176010 257320 176016 257332
rect 176068 257320 176074 257372
rect 255682 257320 255688 257372
rect 255740 257360 255746 257372
rect 583478 257360 583484 257372
rect 255740 257332 583484 257360
rect 255740 257320 255746 257332
rect 583478 257320 583484 257332
rect 583536 257320 583542 257372
rect 104342 256708 104348 256760
rect 104400 256748 104406 256760
rect 110414 256748 110420 256760
rect 104400 256720 110420 256748
rect 104400 256708 104406 256720
rect 110414 256708 110420 256720
rect 110472 256708 110478 256760
rect 125502 256708 125508 256760
rect 125560 256748 125566 256760
rect 127066 256748 127072 256760
rect 125560 256720 127072 256748
rect 125560 256708 125566 256720
rect 127066 256708 127072 256720
rect 127124 256708 127130 256760
rect 173158 256708 173164 256760
rect 173216 256748 173222 256760
rect 191742 256748 191748 256760
rect 173216 256720 191748 256748
rect 173216 256708 173222 256720
rect 191742 256708 191748 256720
rect 191800 256708 191806 256760
rect 50798 256640 50804 256692
rect 50856 256680 50862 256692
rect 66806 256680 66812 256692
rect 50856 256652 66812 256680
rect 50856 256640 50862 256652
rect 66806 256640 66812 256652
rect 66864 256640 66870 256692
rect 255498 256640 255504 256692
rect 255556 256680 255562 256692
rect 258350 256680 258356 256692
rect 255556 256652 258356 256680
rect 255556 256640 255562 256652
rect 258350 256640 258356 256652
rect 258408 256680 258414 256692
rect 582834 256680 582840 256692
rect 258408 256652 582840 256680
rect 258408 256640 258414 256652
rect 582834 256640 582840 256652
rect 582892 256640 582898 256692
rect 100846 255960 100852 256012
rect 100904 256000 100910 256012
rect 113174 256000 113180 256012
rect 100904 255972 113180 256000
rect 100904 255960 100910 255972
rect 113174 255960 113180 255972
rect 113232 255960 113238 256012
rect 142798 255960 142804 256012
rect 142856 256000 142862 256012
rect 155402 256000 155408 256012
rect 142856 255972 155408 256000
rect 142856 255960 142862 255972
rect 155402 255960 155408 255972
rect 155460 255960 155466 256012
rect 255406 255960 255412 256012
rect 255464 256000 255470 256012
rect 270770 256000 270776 256012
rect 255464 255972 270776 256000
rect 255464 255960 255470 255972
rect 270770 255960 270776 255972
rect 270828 255960 270834 256012
rect 270770 255484 270776 255536
rect 270828 255524 270834 255536
rect 271782 255524 271788 255536
rect 270828 255496 271788 255524
rect 270828 255484 270834 255496
rect 271782 255484 271788 255496
rect 271840 255484 271846 255536
rect 49418 255280 49424 255332
rect 49476 255320 49482 255332
rect 50798 255320 50804 255332
rect 49476 255292 50804 255320
rect 49476 255280 49482 255292
rect 50798 255280 50804 255292
rect 50856 255280 50862 255332
rect 100938 255280 100944 255332
rect 100996 255320 101002 255332
rect 106090 255320 106096 255332
rect 100996 255292 106096 255320
rect 100996 255280 101002 255292
rect 106090 255280 106096 255292
rect 106148 255320 106154 255332
rect 133230 255320 133236 255332
rect 106148 255292 133236 255320
rect 106148 255280 106154 255292
rect 133230 255280 133236 255292
rect 133288 255280 133294 255332
rect 148318 255280 148324 255332
rect 148376 255320 148382 255332
rect 191742 255320 191748 255332
rect 148376 255292 191748 255320
rect 148376 255280 148382 255292
rect 191742 255280 191748 255292
rect 191800 255280 191806 255332
rect 276014 254600 276020 254652
rect 276072 254640 276078 254652
rect 298738 254640 298744 254652
rect 276072 254612 298744 254640
rect 276072 254600 276078 254612
rect 298738 254600 298744 254612
rect 298796 254600 298802 254652
rect 102778 254532 102784 254584
rect 102836 254572 102842 254584
rect 123018 254572 123024 254584
rect 102836 254544 123024 254572
rect 102836 254532 102842 254544
rect 123018 254532 123024 254544
rect 123076 254532 123082 254584
rect 269022 254532 269028 254584
rect 269080 254572 269086 254584
rect 583110 254572 583116 254584
rect 269080 254544 583116 254572
rect 269080 254532 269086 254544
rect 583110 254532 583116 254544
rect 583168 254532 583174 254584
rect 151078 253988 151084 254040
rect 151136 254028 151142 254040
rect 191558 254028 191564 254040
rect 151136 254000 191564 254028
rect 151136 253988 151142 254000
rect 191558 253988 191564 254000
rect 191616 253988 191622 254040
rect 255406 253988 255412 254040
rect 255464 254028 255470 254040
rect 267734 254028 267740 254040
rect 255464 254000 267740 254028
rect 255464 253988 255470 254000
rect 267734 253988 267740 254000
rect 267792 254028 267798 254040
rect 269022 254028 269028 254040
rect 267792 254000 269028 254028
rect 267792 253988 267798 254000
rect 269022 253988 269028 254000
rect 269080 253988 269086 254040
rect 49510 253920 49516 253972
rect 49568 253960 49574 253972
rect 66806 253960 66812 253972
rect 49568 253932 66812 253960
rect 49568 253920 49574 253932
rect 66806 253920 66812 253932
rect 66864 253920 66870 253972
rect 106918 253920 106924 253972
rect 106976 253960 106982 253972
rect 180242 253960 180248 253972
rect 106976 253932 180248 253960
rect 106976 253920 106982 253932
rect 180242 253920 180248 253932
rect 180300 253920 180306 253972
rect 255314 253920 255320 253972
rect 255372 253960 255378 253972
rect 276014 253960 276020 253972
rect 255372 253932 276020 253960
rect 255372 253920 255378 253932
rect 276014 253920 276020 253932
rect 276072 253920 276078 253972
rect 15838 253852 15844 253904
rect 15896 253892 15902 253904
rect 35250 253892 35256 253904
rect 15896 253864 35256 253892
rect 15896 253852 15902 253864
rect 35250 253852 35256 253864
rect 35308 253892 35314 253904
rect 35618 253892 35624 253904
rect 35308 253864 35624 253892
rect 35308 253852 35314 253864
rect 35618 253852 35624 253864
rect 35676 253852 35682 253904
rect 266998 253852 267004 253904
rect 267056 253892 267062 253904
rect 268378 253892 268384 253904
rect 267056 253864 268384 253892
rect 267056 253852 267062 253864
rect 268378 253852 268384 253864
rect 268436 253852 268442 253904
rect 35250 253172 35256 253224
rect 35308 253212 35314 253224
rect 66990 253212 66996 253224
rect 35308 253184 66996 253212
rect 35308 253172 35314 253184
rect 66990 253172 66996 253184
rect 67048 253212 67054 253224
rect 67358 253212 67364 253224
rect 67048 253184 67364 253212
rect 67048 253172 67054 253184
rect 67358 253172 67364 253184
rect 67416 253172 67422 253224
rect 128998 253172 129004 253224
rect 129056 253212 129062 253224
rect 173250 253212 173256 253224
rect 129056 253184 173256 253212
rect 129056 253172 129062 253184
rect 173250 253172 173256 253184
rect 173308 253172 173314 253224
rect 271782 253172 271788 253224
rect 271840 253212 271846 253224
rect 583386 253212 583392 253224
rect 271840 253184 583392 253212
rect 271840 253172 271846 253184
rect 583386 253172 583392 253184
rect 583444 253172 583450 253224
rect 188338 252628 188344 252680
rect 188396 252668 188402 252680
rect 191006 252668 191012 252680
rect 188396 252640 191012 252668
rect 188396 252628 188402 252640
rect 191006 252628 191012 252640
rect 191064 252628 191070 252680
rect 255406 252628 255412 252680
rect 255464 252668 255470 252680
rect 266446 252668 266452 252680
rect 255464 252640 266452 252668
rect 255464 252628 255470 252640
rect 266446 252628 266452 252640
rect 266504 252668 266510 252680
rect 266998 252668 267004 252680
rect 266504 252640 267004 252668
rect 266504 252628 266510 252640
rect 266998 252628 267004 252640
rect 267056 252628 267062 252680
rect 107746 252560 107752 252612
rect 107804 252600 107810 252612
rect 111058 252600 111064 252612
rect 107804 252572 111064 252600
rect 107804 252560 107810 252572
rect 111058 252560 111064 252572
rect 111116 252560 111122 252612
rect 170490 252560 170496 252612
rect 170548 252600 170554 252612
rect 191742 252600 191748 252612
rect 170548 252572 191748 252600
rect 170548 252560 170554 252572
rect 191742 252560 191748 252572
rect 191800 252560 191806 252612
rect 255498 252560 255504 252612
rect 255556 252600 255562 252612
rect 270678 252600 270684 252612
rect 255556 252572 270684 252600
rect 255556 252560 255562 252572
rect 270678 252560 270684 252572
rect 270736 252600 270742 252612
rect 271782 252600 271788 252612
rect 270736 252572 271788 252600
rect 270736 252560 270742 252572
rect 271782 252560 271788 252572
rect 271840 252560 271846 252612
rect 100386 252492 100392 252544
rect 100444 252532 100450 252544
rect 120810 252532 120816 252544
rect 100444 252504 120816 252532
rect 100444 252492 100450 252504
rect 120810 252492 120816 252504
rect 120868 252492 120874 252544
rect 109034 252424 109040 252476
rect 109092 252464 109098 252476
rect 109678 252464 109684 252476
rect 109092 252436 109684 252464
rect 109092 252424 109098 252436
rect 109678 252424 109684 252436
rect 109736 252424 109742 252476
rect 263870 252288 263876 252340
rect 263928 252328 263934 252340
rect 266906 252328 266912 252340
rect 263928 252300 266912 252328
rect 263928 252288 263934 252300
rect 266906 252288 266912 252300
rect 266964 252288 266970 252340
rect 163498 251880 163504 251932
rect 163556 251920 163562 251932
rect 188246 251920 188252 251932
rect 163556 251892 188252 251920
rect 163556 251880 163562 251892
rect 188246 251880 188252 251892
rect 188304 251880 188310 251932
rect 38470 251812 38476 251864
rect 38528 251852 38534 251864
rect 45922 251852 45928 251864
rect 38528 251824 45928 251852
rect 38528 251812 38534 251824
rect 45922 251812 45928 251824
rect 45980 251812 45986 251864
rect 135162 251812 135168 251864
rect 135220 251852 135226 251864
rect 170398 251852 170404 251864
rect 135220 251824 170404 251852
rect 135220 251812 135226 251824
rect 170398 251812 170404 251824
rect 170456 251812 170462 251864
rect 259730 251852 259736 251864
rect 258046 251824 259736 251852
rect 255406 251540 255412 251592
rect 255464 251580 255470 251592
rect 258046 251580 258074 251824
rect 259730 251812 259736 251824
rect 259788 251852 259794 251864
rect 582374 251852 582380 251864
rect 259788 251824 582380 251852
rect 259788 251812 259794 251824
rect 582374 251812 582380 251824
rect 582432 251812 582438 251864
rect 255464 251552 258074 251580
rect 255464 251540 255470 251552
rect 45922 251200 45928 251252
rect 45980 251240 45986 251252
rect 46842 251240 46848 251252
rect 45980 251212 46848 251240
rect 45980 251200 45986 251212
rect 46842 251200 46848 251212
rect 46900 251240 46906 251252
rect 66806 251240 66812 251252
rect 46900 251212 66812 251240
rect 46900 251200 46906 251212
rect 66806 251200 66812 251212
rect 66864 251200 66870 251252
rect 109678 251200 109684 251252
rect 109736 251240 109742 251252
rect 134610 251240 134616 251252
rect 109736 251212 134616 251240
rect 109736 251200 109742 251212
rect 134610 251200 134616 251212
rect 134668 251240 134674 251252
rect 135162 251240 135168 251252
rect 134668 251212 135168 251240
rect 134668 251200 134674 251212
rect 135162 251200 135168 251212
rect 135220 251200 135226 251252
rect 186958 251200 186964 251252
rect 187016 251240 187022 251252
rect 191558 251240 191564 251252
rect 187016 251212 191564 251240
rect 187016 251200 187022 251212
rect 191558 251200 191564 251212
rect 191616 251200 191622 251252
rect 255498 251200 255504 251252
rect 255556 251240 255562 251252
rect 262490 251240 262496 251252
rect 255556 251212 262496 251240
rect 255556 251200 255562 251212
rect 262490 251200 262496 251212
rect 262548 251200 262554 251252
rect 61562 250452 61568 250504
rect 61620 250492 61626 250504
rect 66714 250492 66720 250504
rect 61620 250464 66720 250492
rect 61620 250452 61626 250464
rect 66714 250452 66720 250464
rect 66772 250452 66778 250504
rect 100846 250452 100852 250504
rect 100904 250492 100910 250504
rect 107746 250492 107752 250504
rect 100904 250464 107752 250492
rect 100904 250452 100910 250464
rect 107746 250452 107752 250464
rect 107804 250452 107810 250504
rect 112438 250452 112444 250504
rect 112496 250492 112502 250504
rect 114830 250492 114836 250504
rect 112496 250464 114836 250492
rect 112496 250452 112502 250464
rect 114830 250452 114836 250464
rect 114888 250492 114894 250504
rect 130562 250492 130568 250504
rect 114888 250464 130568 250492
rect 114888 250452 114894 250464
rect 130562 250452 130568 250464
rect 130620 250452 130626 250504
rect 133782 250452 133788 250504
rect 133840 250492 133846 250504
rect 147766 250492 147772 250504
rect 133840 250464 147772 250492
rect 133840 250452 133846 250464
rect 147766 250452 147772 250464
rect 147824 250492 147830 250504
rect 192570 250492 192576 250504
rect 147824 250464 192576 250492
rect 147824 250452 147830 250464
rect 192570 250452 192576 250464
rect 192628 250452 192634 250504
rect 265158 250452 265164 250504
rect 265216 250492 265222 250504
rect 582466 250492 582472 250504
rect 265216 250464 582472 250492
rect 265216 250452 265222 250464
rect 582466 250452 582472 250464
rect 582524 250452 582530 250504
rect 255314 249840 255320 249892
rect 255372 249880 255378 249892
rect 265158 249880 265164 249892
rect 255372 249852 265164 249880
rect 255372 249840 255378 249852
rect 265158 249840 265164 249852
rect 265216 249840 265222 249892
rect 56502 249772 56508 249824
rect 56560 249812 56566 249824
rect 56560 249784 61608 249812
rect 56560 249772 56566 249784
rect 61580 249756 61608 249784
rect 100846 249772 100852 249824
rect 100904 249812 100910 249824
rect 132586 249812 132592 249824
rect 100904 249784 132592 249812
rect 100904 249772 100910 249784
rect 132586 249772 132592 249784
rect 132644 249812 132650 249824
rect 133782 249812 133788 249824
rect 132644 249784 133788 249812
rect 132644 249772 132650 249784
rect 133782 249772 133788 249784
rect 133840 249772 133846 249824
rect 170398 249772 170404 249824
rect 170456 249812 170462 249824
rect 191742 249812 191748 249824
rect 170456 249784 191748 249812
rect 170456 249772 170462 249784
rect 191742 249772 191748 249784
rect 191800 249772 191806 249824
rect 255406 249772 255412 249824
rect 255464 249812 255470 249824
rect 266538 249812 266544 249824
rect 255464 249784 266544 249812
rect 255464 249772 255470 249784
rect 266538 249772 266544 249784
rect 266596 249812 266602 249824
rect 582374 249812 582380 249824
rect 266596 249784 582380 249812
rect 266596 249772 266602 249784
rect 582374 249772 582380 249784
rect 582432 249772 582438 249824
rect 61562 249704 61568 249756
rect 61620 249704 61626 249756
rect 100938 249704 100944 249756
rect 100996 249744 101002 249756
rect 111794 249744 111800 249756
rect 100996 249716 111800 249744
rect 100996 249704 101002 249716
rect 111794 249704 111800 249716
rect 111852 249744 111858 249756
rect 112346 249744 112352 249756
rect 111852 249716 112352 249744
rect 111852 249704 111858 249716
rect 112346 249704 112352 249716
rect 112404 249704 112410 249756
rect 112346 249092 112352 249144
rect 112404 249132 112410 249144
rect 131298 249132 131304 249144
rect 112404 249104 131304 249132
rect 112404 249092 112410 249104
rect 131298 249092 131304 249104
rect 131356 249092 131362 249144
rect 100846 249024 100852 249076
rect 100904 249064 100910 249076
rect 106642 249064 106648 249076
rect 100904 249036 106648 249064
rect 100904 249024 100910 249036
rect 106642 249024 106648 249036
rect 106700 249024 106706 249076
rect 122190 249024 122196 249076
rect 122248 249064 122254 249076
rect 124306 249064 124312 249076
rect 122248 249036 124312 249064
rect 122248 249024 122254 249036
rect 124306 249024 124312 249036
rect 124364 249064 124370 249076
rect 187234 249064 187240 249076
rect 124364 249036 187240 249064
rect 124364 249024 124370 249036
rect 187234 249024 187240 249036
rect 187292 249024 187298 249076
rect 255314 248480 255320 248532
rect 255372 248520 255378 248532
rect 268010 248520 268016 248532
rect 255372 248492 268016 248520
rect 255372 248480 255378 248492
rect 268010 248480 268016 248492
rect 268068 248480 268074 248532
rect 111610 248412 111616 248464
rect 111668 248452 111674 248464
rect 114646 248452 114652 248464
rect 111668 248424 114652 248452
rect 111668 248412 111674 248424
rect 114646 248412 114652 248424
rect 114704 248412 114710 248464
rect 180150 248412 180156 248464
rect 180208 248452 180214 248464
rect 190638 248452 190644 248464
rect 180208 248424 190644 248452
rect 180208 248412 180214 248424
rect 190638 248412 190644 248424
rect 190696 248412 190702 248464
rect 255682 248412 255688 248464
rect 255740 248452 255746 248464
rect 271966 248452 271972 248464
rect 255740 248424 271972 248452
rect 255740 248412 255746 248424
rect 271966 248412 271972 248424
rect 272024 248452 272030 248464
rect 582558 248452 582564 248464
rect 272024 248424 582564 248452
rect 272024 248412 272030 248424
rect 582558 248412 582564 248424
rect 582616 248412 582622 248464
rect 100846 248344 100852 248396
rect 100904 248384 100910 248396
rect 108942 248384 108948 248396
rect 100904 248356 108948 248384
rect 100904 248344 100910 248356
rect 108942 248344 108948 248356
rect 109000 248344 109006 248396
rect 42610 247664 42616 247716
rect 42668 247704 42674 247716
rect 52454 247704 52460 247716
rect 42668 247676 52460 247704
rect 42668 247664 42674 247676
rect 52454 247664 52460 247676
rect 52512 247664 52518 247716
rect 108942 247664 108948 247716
rect 109000 247704 109006 247716
rect 124214 247704 124220 247716
rect 109000 247676 124220 247704
rect 109000 247664 109006 247676
rect 124214 247664 124220 247676
rect 124272 247664 124278 247716
rect 254578 247664 254584 247716
rect 254636 247704 254642 247716
rect 582466 247704 582472 247716
rect 254636 247676 582472 247704
rect 254636 247664 254642 247676
rect 582466 247664 582472 247676
rect 582524 247664 582530 247716
rect 62022 247052 62028 247104
rect 62080 247092 62086 247104
rect 67450 247092 67456 247104
rect 62080 247064 67456 247092
rect 62080 247052 62086 247064
rect 67450 247052 67456 247064
rect 67508 247052 67514 247104
rect 188430 247052 188436 247104
rect 188488 247092 188494 247104
rect 191742 247092 191748 247104
rect 188488 247064 191748 247092
rect 188488 247052 188494 247064
rect 191742 247052 191748 247064
rect 191800 247052 191806 247104
rect 255406 247052 255412 247104
rect 255464 247092 255470 247104
rect 341518 247092 341524 247104
rect 255464 247064 341524 247092
rect 255464 247052 255470 247064
rect 341518 247052 341524 247064
rect 341576 247052 341582 247104
rect 100846 246916 100852 246968
rect 100904 246956 100910 246968
rect 104342 246956 104348 246968
rect 100904 246928 104348 246956
rect 100904 246916 100910 246928
rect 104342 246916 104348 246928
rect 104400 246916 104406 246968
rect 100846 246304 100852 246356
rect 100904 246344 100910 246356
rect 109034 246344 109040 246356
rect 100904 246316 109040 246344
rect 100904 246304 100910 246316
rect 109034 246304 109040 246316
rect 109092 246304 109098 246356
rect 120166 246304 120172 246356
rect 120224 246344 120230 246356
rect 178678 246344 178684 246356
rect 120224 246316 178684 246344
rect 120224 246304 120230 246316
rect 178678 246304 178684 246316
rect 178736 246304 178742 246356
rect 59078 246100 59084 246152
rect 59136 246140 59142 246152
rect 66990 246140 66996 246152
rect 59136 246112 66996 246140
rect 59136 246100 59142 246112
rect 66990 246100 66996 246112
rect 67048 246140 67054 246152
rect 67266 246140 67272 246152
rect 67048 246112 67272 246140
rect 67048 246100 67054 246112
rect 67266 246100 67272 246112
rect 67324 246100 67330 246152
rect 253198 245692 253204 245744
rect 253256 245732 253262 245744
rect 313918 245732 313924 245744
rect 253256 245704 313924 245732
rect 253256 245692 253262 245704
rect 313918 245692 313924 245704
rect 313976 245692 313982 245744
rect 184290 245624 184296 245676
rect 184348 245664 184354 245676
rect 191558 245664 191564 245676
rect 184348 245636 191564 245664
rect 184348 245624 184354 245636
rect 191558 245624 191564 245636
rect 191616 245624 191622 245676
rect 255406 245624 255412 245676
rect 255464 245664 255470 245676
rect 258258 245664 258264 245676
rect 255464 245636 258264 245664
rect 255464 245624 255470 245636
rect 258258 245624 258264 245636
rect 258316 245664 258322 245676
rect 583294 245664 583300 245676
rect 258316 245636 583300 245664
rect 258316 245624 258322 245636
rect 583294 245624 583300 245636
rect 583352 245624 583358 245676
rect 100938 245556 100944 245608
rect 100996 245596 101002 245608
rect 109678 245596 109684 245608
rect 100996 245568 109684 245596
rect 100996 245556 101002 245568
rect 109678 245556 109684 245568
rect 109736 245556 109742 245608
rect 254118 244944 254124 244996
rect 254176 244984 254182 244996
rect 255590 244984 255596 244996
rect 254176 244956 255596 244984
rect 254176 244944 254182 244956
rect 255590 244944 255596 244956
rect 255648 244944 255654 244996
rect 55122 244876 55128 244928
rect 55180 244916 55186 244928
rect 64598 244916 64604 244928
rect 55180 244888 64604 244916
rect 55180 244876 55186 244888
rect 64598 244876 64604 244888
rect 64656 244916 64662 244928
rect 66898 244916 66904 244928
rect 64656 244888 66904 244916
rect 64656 244876 64662 244888
rect 66898 244876 66904 244888
rect 66956 244876 66962 244928
rect 122098 244876 122104 244928
rect 122156 244916 122162 244928
rect 142154 244916 142160 244928
rect 122156 244888 142160 244916
rect 122156 244876 122162 244888
rect 142154 244876 142160 244888
rect 142212 244916 142218 244928
rect 143442 244916 143448 244928
rect 142212 244888 143448 244916
rect 142212 244876 142218 244888
rect 143442 244876 143448 244888
rect 143500 244876 143506 244928
rect 255682 244332 255688 244384
rect 255740 244372 255746 244384
rect 349798 244372 349804 244384
rect 255740 244344 349804 244372
rect 255740 244332 255746 244344
rect 349798 244332 349804 244344
rect 349856 244332 349862 244384
rect 100846 244264 100852 244316
rect 100904 244304 100910 244316
rect 124306 244304 124312 244316
rect 100904 244276 124312 244304
rect 100904 244264 100910 244276
rect 124306 244264 124312 244276
rect 124364 244264 124370 244316
rect 143442 244264 143448 244316
rect 143500 244304 143506 244316
rect 193030 244304 193036 244316
rect 143500 244276 193036 244304
rect 143500 244264 143506 244276
rect 193030 244264 193036 244276
rect 193088 244264 193094 244316
rect 260742 244264 260748 244316
rect 260800 244304 260806 244316
rect 583386 244304 583392 244316
rect 260800 244276 583392 244304
rect 260800 244264 260806 244276
rect 583386 244264 583392 244276
rect 583444 244264 583450 244316
rect 103422 243584 103428 243636
rect 103480 243624 103486 243636
rect 106274 243624 106280 243636
rect 103480 243596 106280 243624
rect 103480 243584 103486 243596
rect 106274 243584 106280 243596
rect 106332 243584 106338 243636
rect 105538 243516 105544 243568
rect 105596 243556 105602 243568
rect 111794 243556 111800 243568
rect 105596 243528 111800 243556
rect 105596 243516 105602 243528
rect 111794 243516 111800 243528
rect 111852 243556 111858 243568
rect 163590 243556 163596 243568
rect 111852 243528 163596 243556
rect 111852 243516 111858 243528
rect 163590 243516 163596 243528
rect 163648 243516 163654 243568
rect 255498 243516 255504 243568
rect 255556 243556 255562 243568
rect 262398 243556 262404 243568
rect 255556 243528 262404 243556
rect 255556 243516 255562 243528
rect 262398 243516 262404 243528
rect 262456 243516 262462 243568
rect 187050 242972 187056 243024
rect 187108 243012 187114 243024
rect 191742 243012 191748 243024
rect 187108 242984 191748 243012
rect 187108 242972 187114 242984
rect 191742 242972 191748 242984
rect 191800 242972 191806 243024
rect 261018 243012 261024 243024
rect 258046 242984 261024 243012
rect 49602 242904 49608 242956
rect 49660 242944 49666 242956
rect 55030 242944 55036 242956
rect 49660 242916 55036 242944
rect 49660 242904 49666 242916
rect 55030 242904 55036 242916
rect 55088 242944 55094 242956
rect 66806 242944 66812 242956
rect 55088 242916 66812 242944
rect 55088 242904 55094 242916
rect 66806 242904 66812 242916
rect 66864 242904 66870 242956
rect 98546 242904 98552 242956
rect 98604 242944 98610 242956
rect 99282 242944 99288 242956
rect 98604 242916 99288 242944
rect 98604 242904 98610 242916
rect 99282 242904 99288 242916
rect 99340 242944 99346 242956
rect 103422 242944 103428 242956
rect 99340 242916 103428 242944
rect 99340 242904 99346 242916
rect 103422 242904 103428 242916
rect 103480 242904 103486 242956
rect 117958 242904 117964 242956
rect 118016 242944 118022 242956
rect 193582 242944 193588 242956
rect 118016 242916 193588 242944
rect 118016 242904 118022 242916
rect 193582 242904 193588 242916
rect 193640 242904 193646 242956
rect 255406 242904 255412 242956
rect 255464 242944 255470 242956
rect 258046 242944 258074 242984
rect 261018 242972 261024 242984
rect 261076 243012 261082 243024
rect 304258 243012 304264 243024
rect 261076 242984 304264 243012
rect 261076 242972 261082 242984
rect 304258 242972 304264 242984
rect 304316 242972 304322 243024
rect 255464 242916 258074 242944
rect 255464 242904 255470 242916
rect 262398 242904 262404 242956
rect 262456 242944 262462 242956
rect 583110 242944 583116 242956
rect 262456 242916 583116 242944
rect 262456 242904 262462 242916
rect 583110 242904 583116 242916
rect 583168 242904 583174 242956
rect 253106 242836 253112 242888
rect 253164 242876 253170 242888
rect 255682 242876 255688 242888
rect 253164 242848 255688 242876
rect 253164 242836 253170 242848
rect 255682 242836 255688 242848
rect 255740 242836 255746 242888
rect 100846 242700 100852 242752
rect 100904 242740 100910 242752
rect 104250 242740 104256 242752
rect 100904 242712 104256 242740
rect 100904 242700 100910 242712
rect 104250 242700 104256 242712
rect 104308 242700 104314 242752
rect 54754 242156 54760 242208
rect 54812 242196 54818 242208
rect 69014 242196 69020 242208
rect 54812 242168 69020 242196
rect 54812 242156 54818 242168
rect 69014 242156 69020 242168
rect 69072 242156 69078 242208
rect 118970 242196 118976 242208
rect 94792 242168 118976 242196
rect 94792 241800 94820 242168
rect 118970 242156 118976 242168
rect 119028 242196 119034 242208
rect 180334 242196 180340 242208
rect 119028 242168 180340 242196
rect 119028 242156 119034 242168
rect 180334 242156 180340 242168
rect 180392 242156 180398 242208
rect 255406 242156 255412 242208
rect 255464 242196 255470 242208
rect 582742 242196 582748 242208
rect 255464 242168 582748 242196
rect 255464 242156 255470 242168
rect 582742 242156 582748 242168
rect 582800 242156 582806 242208
rect 251818 241884 251824 241936
rect 251876 241924 251882 241936
rect 254118 241924 254124 241936
rect 251876 241896 254124 241924
rect 251876 241884 251882 241896
rect 254118 241884 254124 241896
rect 254176 241884 254182 241936
rect 250438 241816 250444 241868
rect 250496 241856 250502 241868
rect 253106 241856 253112 241868
rect 250496 241828 253112 241856
rect 250496 241816 250502 241828
rect 253106 241816 253112 241828
rect 253164 241816 253170 241868
rect 69014 241748 69020 241800
rect 69072 241788 69078 241800
rect 69842 241788 69848 241800
rect 69072 241760 69848 241788
rect 69072 241748 69078 241760
rect 69842 241748 69848 241760
rect 69900 241748 69906 241800
rect 94774 241748 94780 241800
rect 94832 241748 94838 241800
rect 68554 241680 68560 241732
rect 68612 241720 68618 241732
rect 69290 241720 69296 241732
rect 68612 241692 69296 241720
rect 68612 241680 68618 241692
rect 69290 241680 69296 241692
rect 69348 241680 69354 241732
rect 111058 241544 111064 241596
rect 111116 241584 111122 241596
rect 193766 241584 193772 241596
rect 111116 241556 193772 241584
rect 111116 241544 111122 241556
rect 193766 241544 193772 241556
rect 193824 241544 193830 241596
rect 57606 241476 57612 241528
rect 57664 241516 57670 241528
rect 77432 241516 77438 241528
rect 57664 241488 77438 241516
rect 57664 241476 57670 241488
rect 77432 241476 77438 241488
rect 77490 241476 77496 241528
rect 193674 241476 193680 241528
rect 193732 241516 193738 241528
rect 213914 241516 213920 241528
rect 193732 241488 213920 241516
rect 193732 241476 193738 241488
rect 213914 241476 213920 241488
rect 213972 241516 213978 241528
rect 214742 241516 214748 241528
rect 213972 241488 214748 241516
rect 213972 241476 213978 241488
rect 214742 241476 214748 241488
rect 214800 241476 214806 241528
rect 255406 241476 255412 241528
rect 255464 241516 255470 241528
rect 263778 241516 263784 241528
rect 255464 241488 263784 241516
rect 255464 241476 255470 241488
rect 263778 241476 263784 241488
rect 263836 241516 263842 241528
rect 291930 241516 291936 241528
rect 263836 241488 291936 241516
rect 263836 241476 263842 241488
rect 291930 241476 291936 241488
rect 291988 241476 291994 241528
rect 46658 241408 46664 241460
rect 46716 241448 46722 241460
rect 71912 241448 71918 241460
rect 46716 241420 71918 241448
rect 46716 241408 46722 241420
rect 71912 241408 71918 241420
rect 71970 241408 71976 241460
rect 117222 241408 117228 241460
rect 117280 241448 117286 241460
rect 255314 241448 255320 241460
rect 117280 241420 255320 241448
rect 117280 241408 117286 241420
rect 255314 241408 255320 241420
rect 255372 241408 255378 241460
rect 193030 241340 193036 241392
rect 193088 241380 193094 241392
rect 199746 241380 199752 241392
rect 193088 241352 199752 241380
rect 193088 241340 193094 241352
rect 199746 241340 199752 241352
rect 199804 241340 199810 241392
rect 249242 241340 249248 241392
rect 249300 241380 249306 241392
rect 253198 241380 253204 241392
rect 249300 241352 253204 241380
rect 249300 241340 249306 241352
rect 253198 241340 253204 241352
rect 253256 241340 253262 241392
rect 2774 241204 2780 241256
rect 2832 241244 2838 241256
rect 4798 241244 4804 241256
rect 2832 241216 4804 241244
rect 2832 241204 2838 241216
rect 4798 241204 4804 241216
rect 4856 241204 4862 241256
rect 84654 240796 84660 240848
rect 84712 240836 84718 240848
rect 112162 240836 112168 240848
rect 84712 240808 112168 240836
rect 84712 240796 84718 240808
rect 112162 240796 112168 240808
rect 112220 240836 112226 240848
rect 115934 240836 115940 240848
rect 112220 240808 115940 240836
rect 112220 240796 112226 240808
rect 115934 240796 115940 240808
rect 115992 240836 115998 240848
rect 117222 240836 117228 240848
rect 115992 240808 117228 240836
rect 115992 240796 115998 240808
rect 117222 240796 117228 240808
rect 117280 240796 117286 240848
rect 14458 240728 14464 240780
rect 14516 240768 14522 240780
rect 88150 240768 88156 240780
rect 14516 240740 88156 240768
rect 14516 240728 14522 240740
rect 88150 240728 88156 240740
rect 88208 240728 88214 240780
rect 255314 240728 255320 240780
rect 255372 240768 255378 240780
rect 580258 240768 580264 240780
rect 255372 240740 580264 240768
rect 255372 240728 255378 240740
rect 580258 240728 580264 240740
rect 580316 240728 580322 240780
rect 74534 240116 74540 240168
rect 74592 240156 74598 240168
rect 74902 240156 74908 240168
rect 74592 240128 74908 240156
rect 74592 240116 74598 240128
rect 74902 240116 74908 240128
rect 74960 240116 74966 240168
rect 77294 240116 77300 240168
rect 77352 240156 77358 240168
rect 78214 240156 78220 240168
rect 77352 240128 78220 240156
rect 77352 240116 77358 240128
rect 78214 240116 78220 240128
rect 78272 240116 78278 240168
rect 83090 240116 83096 240168
rect 83148 240156 83154 240168
rect 83734 240156 83740 240168
rect 83148 240128 83740 240156
rect 83148 240116 83154 240128
rect 83734 240116 83740 240128
rect 83792 240116 83798 240168
rect 85574 240116 85580 240168
rect 85632 240156 85638 240168
rect 85942 240156 85948 240168
rect 85632 240128 85948 240156
rect 85632 240116 85638 240128
rect 85942 240116 85948 240128
rect 86000 240116 86006 240168
rect 88334 240116 88340 240168
rect 88392 240156 88398 240168
rect 88702 240156 88708 240168
rect 88392 240128 88708 240156
rect 88392 240116 88398 240128
rect 88702 240116 88708 240128
rect 88760 240116 88766 240168
rect 91094 240116 91100 240168
rect 91152 240156 91158 240168
rect 92290 240156 92296 240168
rect 91152 240128 92296 240156
rect 91152 240116 91158 240128
rect 92290 240116 92296 240128
rect 92348 240116 92354 240168
rect 96614 240116 96620 240168
rect 96672 240156 96678 240168
rect 96982 240156 96988 240168
rect 96672 240128 96988 240156
rect 96672 240116 96678 240128
rect 96982 240116 96988 240128
rect 97040 240116 97046 240168
rect 55950 240048 55956 240100
rect 56008 240088 56014 240100
rect 56226 240088 56232 240100
rect 56008 240060 56232 240088
rect 56008 240048 56014 240060
rect 56226 240048 56232 240060
rect 56284 240088 56290 240100
rect 87046 240088 87052 240100
rect 56284 240060 87052 240088
rect 56284 240048 56290 240060
rect 87046 240048 87052 240060
rect 87104 240048 87110 240100
rect 93854 240048 93860 240100
rect 93912 240088 93918 240100
rect 94222 240088 94228 240100
rect 93912 240060 94228 240088
rect 93912 240048 93918 240060
rect 94222 240048 94228 240060
rect 94280 240048 94286 240100
rect 103422 240048 103428 240100
rect 103480 240088 103486 240100
rect 194778 240088 194784 240100
rect 103480 240060 194784 240088
rect 103480 240048 103486 240060
rect 194778 240048 194784 240060
rect 194836 240048 194842 240100
rect 250622 240048 250628 240100
rect 250680 240088 250686 240100
rect 253014 240088 253020 240100
rect 250680 240060 253020 240088
rect 250680 240048 250686 240060
rect 253014 240048 253020 240060
rect 253072 240048 253078 240100
rect 64506 239980 64512 240032
rect 64564 240020 64570 240032
rect 74626 240020 74632 240032
rect 64564 239992 74632 240020
rect 64564 239980 64570 239992
rect 74626 239980 74632 239992
rect 74684 239980 74690 240032
rect 82998 239980 83004 240032
rect 83056 240020 83062 240032
rect 84010 240020 84016 240032
rect 83056 239992 84016 240020
rect 83056 239980 83062 239992
rect 84010 239980 84016 239992
rect 84068 239980 84074 240032
rect 128538 239980 128544 240032
rect 128596 240020 128602 240032
rect 212258 240020 212264 240032
rect 128596 239992 212264 240020
rect 128596 239980 128602 239992
rect 212258 239980 212264 239992
rect 212316 239980 212322 240032
rect 80054 239436 80060 239488
rect 80112 239476 80118 239488
rect 80422 239476 80428 239488
rect 80112 239448 80428 239476
rect 80112 239436 80118 239448
rect 80422 239436 80428 239448
rect 80480 239436 80486 239488
rect 252646 239436 252652 239488
rect 252704 239476 252710 239488
rect 261110 239476 261116 239488
rect 252704 239448 261116 239476
rect 252704 239436 252710 239448
rect 261110 239436 261116 239448
rect 261168 239436 261174 239488
rect 11698 239368 11704 239420
rect 11756 239408 11762 239420
rect 52362 239408 52368 239420
rect 11756 239380 52368 239408
rect 11756 239368 11762 239380
rect 52362 239368 52368 239380
rect 52420 239408 52426 239420
rect 55950 239408 55956 239420
rect 52420 239380 55956 239408
rect 52420 239368 52426 239380
rect 55950 239368 55956 239380
rect 56008 239368 56014 239420
rect 89622 239368 89628 239420
rect 89680 239408 89686 239420
rect 106458 239408 106464 239420
rect 89680 239380 106464 239408
rect 89680 239368 89686 239380
rect 106458 239368 106464 239380
rect 106516 239408 106522 239420
rect 128538 239408 128544 239420
rect 106516 239380 128544 239408
rect 106516 239368 106522 239380
rect 128538 239368 128544 239380
rect 128596 239368 128602 239420
rect 243630 239368 243636 239420
rect 243688 239408 243694 239420
rect 254578 239408 254584 239420
rect 243688 239380 254584 239408
rect 243688 239368 243694 239380
rect 254578 239368 254584 239380
rect 254636 239368 254642 239420
rect 249150 238796 249156 238808
rect 231826 238768 249156 238796
rect 38562 238688 38568 238740
rect 38620 238728 38626 238740
rect 69106 238728 69112 238740
rect 38620 238700 69112 238728
rect 38620 238688 38626 238700
rect 69106 238688 69112 238700
rect 69164 238688 69170 238740
rect 69842 238688 69848 238740
rect 69900 238728 69906 238740
rect 80146 238728 80152 238740
rect 69900 238700 80152 238728
rect 69900 238688 69906 238700
rect 80146 238688 80152 238700
rect 80204 238688 80210 238740
rect 83182 238688 83188 238740
rect 83240 238728 83246 238740
rect 103514 238728 103520 238740
rect 83240 238700 103520 238728
rect 83240 238688 83246 238700
rect 103514 238688 103520 238700
rect 103572 238688 103578 238740
rect 192570 238688 192576 238740
rect 192628 238728 192634 238740
rect 231826 238728 231854 238768
rect 249150 238756 249156 238768
rect 249208 238756 249214 238808
rect 258350 238756 258356 238808
rect 258408 238796 258414 238808
rect 580350 238796 580356 238808
rect 258408 238768 580356 238796
rect 258408 238756 258414 238768
rect 580350 238756 580356 238768
rect 580408 238756 580414 238808
rect 192628 238700 231854 238728
rect 192628 238688 192634 238700
rect 53098 238620 53104 238672
rect 53156 238660 53162 238672
rect 74534 238660 74540 238672
rect 53156 238632 74540 238660
rect 53156 238620 53162 238632
rect 74534 238620 74540 238632
rect 74592 238620 74598 238672
rect 88058 238620 88064 238672
rect 88116 238660 88122 238672
rect 104986 238660 104992 238672
rect 88116 238632 104992 238660
rect 88116 238620 88122 238632
rect 104986 238620 104992 238632
rect 105044 238620 105050 238672
rect 180242 238620 180248 238672
rect 180300 238660 180306 238672
rect 197262 238660 197268 238672
rect 180300 238632 197268 238660
rect 180300 238620 180306 238632
rect 197262 238620 197268 238632
rect 197320 238620 197326 238672
rect 87046 238076 87052 238128
rect 87104 238116 87110 238128
rect 88058 238116 88064 238128
rect 87104 238088 88064 238116
rect 87104 238076 87110 238088
rect 88058 238076 88064 238088
rect 88116 238076 88122 238128
rect 104250 238008 104256 238060
rect 104308 238048 104314 238060
rect 114738 238048 114744 238060
rect 104308 238020 114744 238048
rect 104308 238008 104314 238020
rect 114738 238008 114744 238020
rect 114796 238008 114802 238060
rect 119338 238008 119344 238060
rect 119396 238048 119402 238060
rect 191282 238048 191288 238060
rect 119396 238020 191288 238048
rect 119396 238008 119402 238020
rect 191282 238008 191288 238020
rect 191340 238008 191346 238060
rect 232222 238008 232228 238060
rect 232280 238048 232286 238060
rect 241514 238048 241520 238060
rect 232280 238020 241520 238048
rect 232280 238008 232286 238020
rect 241514 238008 241520 238020
rect 241572 238008 241578 238060
rect 243538 238008 243544 238060
rect 243596 238048 243602 238060
rect 258166 238048 258172 238060
rect 243596 238020 258172 238048
rect 243596 238008 243602 238020
rect 258166 238008 258172 238020
rect 258224 238008 258230 238060
rect 69106 237396 69112 237448
rect 69164 237436 69170 237448
rect 69658 237436 69664 237448
rect 69164 237408 69664 237436
rect 69164 237396 69170 237408
rect 69658 237396 69664 237408
rect 69716 237396 69722 237448
rect 80146 237396 80152 237448
rect 80204 237436 80210 237448
rect 80698 237436 80704 237448
rect 80204 237408 80704 237436
rect 80204 237396 80210 237408
rect 80698 237396 80704 237408
rect 80756 237396 80762 237448
rect 82722 237396 82728 237448
rect 82780 237436 82786 237448
rect 83182 237436 83188 237448
rect 82780 237408 83188 237436
rect 82780 237396 82786 237408
rect 83182 237396 83188 237408
rect 83240 237396 83246 237448
rect 39666 237328 39672 237380
rect 39724 237368 39730 237380
rect 73246 237368 73252 237380
rect 39724 237340 73252 237368
rect 39724 237328 39730 237340
rect 73246 237328 73252 237340
rect 73304 237328 73310 237380
rect 88150 237328 88156 237380
rect 88208 237368 88214 237380
rect 92566 237368 92572 237380
rect 88208 237340 92572 237368
rect 88208 237328 88214 237340
rect 92566 237328 92572 237340
rect 92624 237368 92630 237380
rect 92624 237340 93854 237368
rect 92624 237328 92630 237340
rect 93826 237300 93854 237340
rect 102226 237328 102232 237380
rect 102284 237368 102290 237380
rect 252830 237368 252836 237380
rect 102284 237340 252836 237368
rect 102284 237328 102290 237340
rect 252830 237328 252836 237340
rect 252888 237328 252894 237380
rect 111886 237300 111892 237312
rect 93826 237272 111892 237300
rect 111886 237260 111892 237272
rect 111944 237260 111950 237312
rect 187234 237260 187240 237312
rect 187292 237300 187298 237312
rect 224770 237300 224776 237312
rect 187292 237272 224776 237300
rect 187292 237260 187298 237272
rect 224770 237260 224776 237272
rect 224828 237260 224834 237312
rect 74718 236716 74724 236768
rect 74776 236756 74782 236768
rect 89162 236756 89168 236768
rect 74776 236728 89168 236756
rect 74776 236716 74782 236728
rect 89162 236716 89168 236728
rect 89220 236716 89226 236768
rect 60458 236648 60464 236700
rect 60516 236688 60522 236700
rect 76098 236688 76104 236700
rect 60516 236660 76104 236688
rect 60516 236648 60522 236660
rect 76098 236648 76104 236660
rect 76156 236648 76162 236700
rect 93118 236648 93124 236700
rect 93176 236688 93182 236700
rect 102226 236688 102232 236700
rect 93176 236660 102232 236688
rect 93176 236648 93182 236660
rect 102226 236648 102232 236660
rect 102284 236648 102290 236700
rect 253198 236648 253204 236700
rect 253256 236688 253262 236700
rect 263686 236688 263692 236700
rect 253256 236660 263692 236688
rect 253256 236648 253262 236660
rect 263686 236648 263692 236660
rect 263744 236648 263750 236700
rect 90818 235968 90824 236020
rect 90876 236008 90882 236020
rect 91094 236008 91100 236020
rect 90876 235980 91100 236008
rect 90876 235968 90882 235980
rect 91094 235968 91100 235980
rect 91152 235968 91158 236020
rect 67358 235900 67364 235952
rect 67416 235940 67422 235952
rect 111058 235940 111064 235952
rect 67416 235912 111064 235940
rect 67416 235900 67422 235912
rect 111058 235900 111064 235912
rect 111116 235900 111122 235952
rect 180334 235900 180340 235952
rect 180392 235940 180398 235952
rect 202230 235940 202236 235952
rect 180392 235912 202236 235940
rect 180392 235900 180398 235912
rect 202230 235900 202236 235912
rect 202288 235940 202294 235952
rect 202782 235940 202788 235952
rect 202288 235912 202788 235940
rect 202288 235900 202294 235912
rect 202782 235900 202788 235912
rect 202840 235900 202846 235952
rect 50982 235832 50988 235884
rect 51040 235872 51046 235884
rect 77294 235872 77300 235884
rect 51040 235844 77300 235872
rect 51040 235832 51046 235844
rect 77294 235832 77300 235844
rect 77352 235832 77358 235884
rect 94038 235492 94044 235544
rect 94096 235532 94102 235544
rect 94498 235532 94504 235544
rect 94096 235504 94504 235532
rect 94096 235492 94102 235504
rect 94498 235492 94504 235504
rect 94556 235532 94562 235544
rect 102318 235532 102324 235544
rect 94556 235504 102324 235532
rect 94556 235492 94562 235504
rect 102318 235492 102324 235504
rect 102376 235492 102382 235544
rect 84102 235220 84108 235272
rect 84160 235260 84166 235272
rect 89714 235260 89720 235272
rect 84160 235232 89720 235260
rect 84160 235220 84166 235232
rect 89714 235220 89720 235232
rect 89772 235220 89778 235272
rect 102778 235220 102784 235272
rect 102836 235260 102842 235272
rect 107010 235260 107016 235272
rect 102836 235232 107016 235260
rect 102836 235220 102842 235232
rect 107010 235220 107016 235232
rect 107068 235220 107074 235272
rect 134702 235220 134708 235272
rect 134760 235260 134766 235272
rect 142890 235260 142896 235272
rect 134760 235232 142896 235260
rect 134760 235220 134766 235232
rect 142890 235220 142896 235232
rect 142948 235220 142954 235272
rect 202782 235220 202788 235272
rect 202840 235260 202846 235272
rect 246298 235260 246304 235272
rect 202840 235232 246304 235260
rect 202840 235220 202846 235232
rect 246298 235220 246304 235232
rect 246356 235220 246362 235272
rect 217318 234608 217324 234660
rect 217376 234648 217382 234660
rect 266998 234648 267004 234660
rect 217376 234620 267004 234648
rect 217376 234608 217382 234620
rect 266998 234608 267004 234620
rect 267056 234608 267062 234660
rect 80054 234540 80060 234592
rect 80112 234580 80118 234592
rect 111794 234580 111800 234592
rect 80112 234552 111800 234580
rect 80112 234540 80118 234552
rect 111794 234540 111800 234552
rect 111852 234540 111858 234592
rect 117682 234540 117688 234592
rect 117740 234580 117746 234592
rect 117958 234580 117964 234592
rect 117740 234552 117964 234580
rect 117740 234540 117746 234552
rect 117958 234540 117964 234552
rect 118016 234580 118022 234592
rect 122190 234580 122196 234592
rect 118016 234552 122196 234580
rect 118016 234540 118022 234552
rect 122190 234540 122196 234552
rect 122248 234540 122254 234592
rect 182910 234540 182916 234592
rect 182968 234580 182974 234592
rect 254026 234580 254032 234592
rect 182968 234552 254032 234580
rect 182968 234540 182974 234552
rect 254026 234540 254032 234552
rect 254084 234540 254090 234592
rect 193674 234472 193680 234524
rect 193732 234512 193738 234524
rect 219710 234512 219716 234524
rect 193732 234484 219716 234512
rect 193732 234472 193738 234484
rect 219710 234472 219716 234484
rect 219768 234472 219774 234524
rect 68278 233928 68284 233980
rect 68336 233968 68342 233980
rect 80422 233968 80428 233980
rect 68336 233940 80428 233968
rect 68336 233928 68342 233940
rect 80422 233928 80428 233940
rect 80480 233928 80486 233980
rect 4798 233860 4804 233912
rect 4856 233900 4862 233912
rect 97810 233900 97816 233912
rect 4856 233872 97816 233900
rect 4856 233860 4862 233872
rect 97810 233860 97816 233872
rect 97868 233860 97874 233912
rect 114462 233860 114468 233912
rect 114520 233900 114526 233912
rect 115934 233900 115940 233912
rect 114520 233872 115940 233900
rect 114520 233860 114526 233872
rect 115934 233860 115940 233872
rect 115992 233860 115998 233912
rect 122098 233860 122104 233912
rect 122156 233900 122162 233912
rect 191098 233900 191104 233912
rect 122156 233872 191104 233900
rect 122156 233860 122162 233872
rect 191098 233860 191104 233872
rect 191156 233860 191162 233912
rect 100662 233248 100668 233300
rect 100720 233288 100726 233300
rect 100846 233288 100852 233300
rect 100720 233260 100852 233288
rect 100720 233248 100726 233260
rect 100846 233248 100852 233260
rect 100904 233248 100910 233300
rect 103514 233248 103520 233300
rect 103572 233288 103578 233300
rect 114646 233288 114652 233300
rect 103572 233260 114652 233288
rect 103572 233248 103578 233260
rect 114646 233248 114652 233260
rect 114704 233288 114710 233300
rect 138658 233288 138664 233300
rect 114704 233260 138664 233288
rect 114704 233248 114710 233260
rect 138658 233248 138664 233260
rect 138716 233248 138722 233300
rect 236638 233248 236644 233300
rect 236696 233288 236702 233300
rect 237190 233288 237196 233300
rect 236696 233260 237196 233288
rect 236696 233248 236702 233260
rect 237190 233248 237196 233260
rect 237248 233288 237254 233300
rect 298094 233288 298100 233300
rect 237248 233260 298100 233288
rect 237248 233248 237254 233260
rect 298094 233248 298100 233260
rect 298152 233248 298158 233300
rect 76650 233180 76656 233232
rect 76708 233220 76714 233232
rect 78674 233220 78680 233232
rect 76708 233192 78680 233220
rect 76708 233180 76714 233192
rect 78674 233180 78680 233192
rect 78732 233220 78738 233232
rect 80974 233220 80980 233232
rect 78732 233192 80980 233220
rect 78732 233180 78738 233192
rect 80974 233180 80980 233192
rect 81032 233180 81038 233232
rect 106918 233220 106924 233232
rect 86926 233192 106924 233220
rect 72786 233112 72792 233164
rect 72844 233152 72850 233164
rect 75914 233152 75920 233164
rect 72844 233124 75920 233152
rect 72844 233112 72850 233124
rect 75914 233112 75920 233124
rect 75972 233112 75978 233164
rect 86926 233152 86954 233192
rect 106918 233180 106924 233192
rect 106976 233180 106982 233232
rect 193766 233180 193772 233232
rect 193824 233220 193830 233232
rect 259546 233220 259552 233232
rect 193824 233192 259552 233220
rect 193824 233180 193830 233192
rect 259546 233180 259552 233192
rect 259604 233180 259610 233232
rect 109310 233152 109316 233164
rect 77266 233124 86954 233152
rect 89686 233124 109316 233152
rect 74810 233044 74816 233096
rect 74868 233084 74874 233096
rect 77266 233084 77294 233124
rect 74868 233056 77294 233084
rect 74868 233044 74874 233056
rect 80974 232976 80980 233028
rect 81032 233016 81038 233028
rect 89686 233016 89714 233124
rect 109310 233112 109316 233124
rect 109368 233112 109374 233164
rect 81032 232988 89714 233016
rect 81032 232976 81038 232988
rect 43806 232500 43812 232552
rect 43864 232540 43870 232552
rect 71958 232540 71964 232552
rect 43864 232512 71964 232540
rect 43864 232500 43870 232512
rect 71958 232500 71964 232512
rect 72016 232540 72022 232552
rect 72786 232540 72792 232552
rect 72016 232512 72792 232540
rect 72016 232500 72022 232512
rect 72786 232500 72792 232512
rect 72844 232500 72850 232552
rect 199746 232500 199752 232552
rect 199804 232540 199810 232552
rect 250438 232540 250444 232552
rect 199804 232512 250444 232540
rect 199804 232500 199810 232512
rect 250438 232500 250444 232512
rect 250496 232500 250502 232552
rect 255958 231820 255964 231872
rect 256016 231860 256022 231872
rect 582558 231860 582564 231872
rect 256016 231832 582564 231860
rect 256016 231820 256022 231832
rect 582558 231820 582564 231832
rect 582616 231820 582622 231872
rect 174538 231752 174544 231804
rect 174596 231792 174602 231804
rect 256786 231792 256792 231804
rect 174596 231764 256792 231792
rect 174596 231752 174602 231764
rect 256786 231752 256792 231764
rect 256844 231752 256850 231804
rect 207198 231684 207204 231736
rect 207256 231724 207262 231736
rect 207658 231724 207664 231736
rect 207256 231696 207664 231724
rect 207256 231684 207262 231696
rect 207658 231684 207664 231696
rect 207716 231684 207722 231736
rect 39942 231072 39948 231124
rect 40000 231112 40006 231124
rect 189810 231112 189816 231124
rect 40000 231084 189816 231112
rect 40000 231072 40006 231084
rect 189810 231072 189816 231084
rect 189868 231072 189874 231124
rect 207658 230460 207664 230512
rect 207716 230500 207722 230512
rect 270586 230500 270592 230512
rect 207716 230472 270592 230500
rect 207716 230460 207722 230472
rect 270586 230460 270592 230472
rect 270644 230460 270650 230512
rect 133230 230392 133236 230444
rect 133288 230432 133294 230444
rect 263870 230432 263876 230444
rect 133288 230404 263876 230432
rect 133288 230392 133294 230404
rect 263870 230392 263876 230404
rect 263928 230392 263934 230444
rect 80330 229780 80336 229832
rect 80388 229820 80394 229832
rect 92382 229820 92388 229832
rect 80388 229792 92388 229820
rect 80388 229780 80394 229792
rect 92382 229780 92388 229792
rect 92440 229820 92446 229832
rect 114830 229820 114836 229832
rect 92440 229792 114836 229820
rect 92440 229780 92446 229792
rect 114830 229780 114836 229792
rect 114888 229780 114894 229832
rect 12342 229712 12348 229764
rect 12400 229752 12406 229764
rect 191834 229752 191840 229764
rect 12400 229724 191840 229752
rect 12400 229712 12406 229724
rect 191834 229712 191840 229724
rect 191892 229712 191898 229764
rect 193214 229712 193220 229764
rect 193272 229752 193278 229764
rect 251266 229752 251272 229764
rect 193272 229724 251272 229752
rect 193272 229712 193278 229724
rect 251266 229712 251272 229724
rect 251324 229712 251330 229764
rect 122742 229100 122748 229152
rect 122800 229140 122806 229152
rect 123110 229140 123116 229152
rect 122800 229112 123116 229140
rect 122800 229100 122806 229112
rect 123110 229100 123116 229112
rect 123168 229100 123174 229152
rect 119430 228556 119436 228608
rect 119488 228596 119494 228608
rect 120258 228596 120264 228608
rect 119488 228568 120264 228596
rect 119488 228556 119494 228568
rect 120258 228556 120264 228568
rect 120316 228556 120322 228608
rect 57698 228352 57704 228404
rect 57756 228392 57762 228404
rect 70394 228392 70400 228404
rect 57756 228364 70400 228392
rect 57756 228352 57762 228364
rect 70394 228352 70400 228364
rect 70452 228352 70458 228404
rect 252922 228392 252928 228404
rect 122806 228364 252928 228392
rect 120258 228284 120264 228336
rect 120316 228324 120322 228336
rect 122806 228324 122834 228364
rect 252922 228352 252928 228364
rect 252980 228352 252986 228404
rect 255498 228352 255504 228404
rect 255556 228392 255562 228404
rect 583202 228392 583208 228404
rect 255556 228364 583208 228392
rect 255556 228352 255562 228364
rect 583202 228352 583208 228364
rect 583260 228352 583266 228404
rect 120316 228296 122834 228324
rect 120316 228284 120322 228296
rect 81434 227944 81440 227996
rect 81492 227984 81498 227996
rect 85574 227984 85580 227996
rect 81492 227956 85580 227984
rect 81492 227944 81498 227956
rect 85574 227944 85580 227956
rect 85632 227944 85638 227996
rect 92198 227808 92204 227860
rect 92256 227848 92262 227860
rect 92256 227820 93854 227848
rect 92256 227808 92262 227820
rect 88334 227740 88340 227792
rect 88392 227780 88398 227792
rect 93118 227780 93124 227792
rect 88392 227752 93124 227780
rect 88392 227740 88398 227752
rect 93118 227740 93124 227752
rect 93176 227740 93182 227792
rect 93826 227780 93854 227820
rect 94498 227780 94504 227792
rect 93826 227752 94504 227780
rect 94498 227740 94504 227752
rect 94556 227740 94562 227792
rect 95970 227740 95976 227792
rect 96028 227780 96034 227792
rect 100754 227780 100760 227792
rect 96028 227752 100760 227780
rect 96028 227740 96034 227752
rect 100754 227740 100760 227752
rect 100812 227740 100818 227792
rect 209774 227740 209780 227792
rect 209832 227780 209838 227792
rect 256050 227780 256056 227792
rect 209832 227752 256056 227780
rect 209832 227740 209838 227752
rect 256050 227740 256056 227752
rect 256108 227740 256114 227792
rect 95142 227672 95148 227724
rect 95200 227712 95206 227724
rect 128998 227712 129004 227724
rect 95200 227684 129004 227712
rect 95200 227672 95206 227684
rect 128998 227672 129004 227684
rect 129056 227672 129062 227724
rect 181530 227672 181536 227724
rect 181588 227712 181594 227724
rect 244734 227712 244740 227724
rect 181588 227684 244740 227712
rect 181588 227672 181594 227684
rect 244734 227672 244740 227684
rect 244792 227672 244798 227724
rect 82078 227604 82084 227656
rect 82136 227644 82142 227656
rect 103514 227644 103520 227656
rect 82136 227616 103520 227644
rect 82136 227604 82142 227616
rect 103514 227604 103520 227616
rect 103572 227604 103578 227656
rect 108298 226992 108304 227044
rect 108356 227032 108362 227044
rect 191190 227032 191196 227044
rect 108356 227004 191196 227032
rect 108356 226992 108362 227004
rect 191190 226992 191196 227004
rect 191248 226992 191254 227044
rect 234614 226992 234620 227044
rect 234672 227032 234678 227044
rect 291838 227032 291844 227044
rect 234672 227004 291844 227032
rect 234672 226992 234678 227004
rect 291838 226992 291844 227004
rect 291896 226992 291902 227044
rect 291930 226992 291936 227044
rect 291988 227032 291994 227044
rect 582374 227032 582380 227044
rect 291988 227004 582380 227032
rect 291988 226992 291994 227004
rect 582374 226992 582380 227004
rect 582432 226992 582438 227044
rect 68922 226312 68928 226364
rect 68980 226352 68986 226364
rect 71774 226352 71780 226364
rect 68980 226324 71780 226352
rect 68980 226312 68986 226324
rect 71774 226312 71780 226324
rect 71832 226312 71838 226364
rect 128538 226312 128544 226364
rect 128596 226352 128602 226364
rect 128998 226352 129004 226364
rect 128596 226324 129004 226352
rect 128596 226312 128602 226324
rect 128998 226312 129004 226324
rect 129056 226312 129062 226364
rect 52178 226244 52184 226296
rect 52236 226284 52242 226296
rect 77386 226284 77392 226296
rect 52236 226256 77392 226284
rect 52236 226244 52242 226256
rect 77386 226244 77392 226256
rect 77444 226284 77450 226296
rect 78582 226284 78588 226296
rect 77444 226256 78588 226284
rect 77444 226244 77450 226256
rect 78582 226244 78588 226256
rect 78640 226244 78646 226296
rect 125686 226244 125692 226296
rect 125744 226284 125750 226296
rect 265066 226284 265072 226296
rect 125744 226256 265072 226284
rect 125744 226244 125750 226256
rect 265066 226244 265072 226256
rect 265124 226244 265130 226296
rect 88242 225632 88248 225684
rect 88300 225672 88306 225684
rect 102134 225672 102140 225684
rect 88300 225644 102140 225672
rect 88300 225632 88306 225644
rect 102134 225632 102140 225644
rect 102192 225632 102198 225684
rect 101490 225564 101496 225616
rect 101548 225604 101554 225616
rect 111978 225604 111984 225616
rect 101548 225576 111984 225604
rect 101548 225564 101554 225576
rect 111978 225564 111984 225576
rect 112036 225604 112042 225616
rect 125686 225604 125692 225616
rect 112036 225576 125692 225604
rect 112036 225564 112042 225576
rect 125686 225564 125692 225576
rect 125744 225564 125750 225616
rect 251910 224952 251916 225004
rect 251968 224992 251974 225004
rect 351914 224992 351920 225004
rect 251968 224964 351920 224992
rect 251968 224952 251974 224964
rect 351914 224952 351920 224964
rect 351972 224952 351978 225004
rect 88426 224884 88432 224936
rect 88484 224924 88490 224936
rect 115934 224924 115940 224936
rect 88484 224896 115940 224924
rect 88484 224884 88490 224896
rect 115934 224884 115940 224896
rect 115992 224884 115998 224936
rect 136542 224884 136548 224936
rect 136600 224924 136606 224936
rect 255958 224924 255964 224936
rect 136600 224896 255964 224924
rect 136600 224884 136606 224896
rect 255958 224884 255964 224896
rect 256016 224884 256022 224936
rect 52270 224204 52276 224256
rect 52328 224244 52334 224256
rect 76742 224244 76748 224256
rect 52328 224216 76748 224244
rect 52328 224204 52334 224216
rect 76742 224204 76748 224216
rect 76800 224204 76806 224256
rect 131758 224204 131764 224256
rect 131816 224244 131822 224256
rect 135438 224244 135444 224256
rect 131816 224216 135444 224244
rect 131816 224204 131822 224216
rect 135438 224204 135444 224216
rect 135496 224244 135502 224256
rect 136542 224244 136548 224256
rect 135496 224216 136548 224244
rect 135496 224204 135502 224216
rect 136542 224204 136548 224216
rect 136600 224204 136606 224256
rect 89714 224136 89720 224188
rect 89772 224176 89778 224188
rect 94774 224176 94780 224188
rect 89772 224148 94780 224176
rect 89772 224136 89778 224148
rect 94774 224136 94780 224148
rect 94832 224136 94838 224188
rect 229738 223592 229744 223644
rect 229796 223632 229802 223644
rect 288434 223632 288440 223644
rect 229796 223604 288440 223632
rect 229796 223592 229802 223604
rect 288434 223592 288440 223604
rect 288492 223592 288498 223644
rect 130470 223524 130476 223576
rect 130528 223564 130534 223576
rect 131022 223564 131028 223576
rect 130528 223536 131028 223564
rect 130528 223524 130534 223536
rect 131022 223524 131028 223536
rect 131080 223564 131086 223576
rect 222194 223564 222200 223576
rect 131080 223536 222200 223564
rect 131080 223524 131086 223536
rect 222194 223524 222200 223536
rect 222252 223524 222258 223576
rect 184382 223456 184388 223508
rect 184440 223496 184446 223508
rect 265158 223496 265164 223508
rect 184440 223468 265164 223496
rect 184440 223456 184446 223468
rect 265158 223456 265164 223468
rect 265216 223456 265222 223508
rect 86862 222844 86868 222896
rect 86920 222884 86926 222896
rect 112070 222884 112076 222896
rect 86920 222856 112076 222884
rect 86920 222844 86926 222856
rect 112070 222844 112076 222856
rect 112128 222844 112134 222896
rect 242250 222164 242256 222216
rect 242308 222204 242314 222216
rect 306374 222204 306380 222216
rect 242308 222176 306380 222204
rect 242308 222164 242314 222176
rect 306374 222164 306380 222176
rect 306432 222164 306438 222216
rect 50338 222096 50344 222148
rect 50396 222136 50402 222148
rect 50890 222136 50896 222148
rect 50396 222108 50896 222136
rect 50396 222096 50402 222108
rect 50890 222096 50896 222108
rect 50948 222136 50954 222148
rect 266538 222136 266544 222148
rect 50948 222108 266544 222136
rect 50948 222096 50954 222108
rect 266538 222096 266544 222108
rect 266596 222096 266602 222148
rect 126238 221416 126244 221468
rect 126296 221456 126302 221468
rect 234706 221456 234712 221468
rect 126296 221428 234712 221456
rect 126296 221416 126302 221428
rect 234706 221416 234712 221428
rect 234764 221416 234770 221468
rect 244734 221416 244740 221468
rect 244792 221456 244798 221468
rect 309778 221456 309784 221468
rect 244792 221428 309784 221456
rect 244792 221416 244798 221428
rect 309778 221416 309784 221428
rect 309836 221416 309842 221468
rect 98638 220804 98644 220856
rect 98696 220844 98702 220856
rect 126882 220844 126888 220856
rect 98696 220816 126888 220844
rect 98696 220804 98702 220816
rect 126882 220804 126888 220816
rect 126940 220804 126946 220856
rect 69658 220736 69664 220788
rect 69716 220776 69722 220788
rect 209774 220776 209780 220788
rect 69716 220748 209780 220776
rect 69716 220736 69722 220748
rect 209774 220736 209780 220748
rect 209832 220736 209838 220788
rect 247218 220736 247224 220788
rect 247276 220776 247282 220788
rect 247678 220776 247684 220788
rect 247276 220748 247684 220776
rect 247276 220736 247282 220748
rect 247678 220736 247684 220748
rect 247736 220736 247742 220788
rect 58986 220056 58992 220108
rect 59044 220096 59050 220108
rect 71774 220096 71780 220108
rect 59044 220068 71780 220096
rect 59044 220056 59050 220068
rect 71774 220056 71780 220068
rect 71832 220056 71838 220108
rect 247678 219444 247684 219496
rect 247736 219484 247742 219496
rect 331214 219484 331220 219496
rect 247736 219456 331220 219484
rect 247736 219444 247742 219456
rect 331214 219444 331220 219456
rect 331272 219444 331278 219496
rect 41138 219376 41144 219428
rect 41196 219416 41202 219428
rect 243630 219416 243636 219428
rect 41196 219388 243636 219416
rect 41196 219376 41202 219388
rect 243630 219376 243636 219388
rect 243688 219376 243694 219428
rect 268378 219376 268384 219428
rect 268436 219416 268442 219428
rect 580166 219416 580172 219428
rect 268436 219388 580172 219416
rect 268436 219376 268442 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 107562 218696 107568 218748
rect 107620 218736 107626 218748
rect 177390 218736 177396 218748
rect 107620 218708 177396 218736
rect 107620 218696 107626 218708
rect 177390 218696 177396 218708
rect 177448 218696 177454 218748
rect 213914 218696 213920 218748
rect 213972 218736 213978 218748
rect 267918 218736 267924 218748
rect 213972 218708 267924 218736
rect 213972 218696 213978 218708
rect 267918 218696 267924 218708
rect 267976 218696 267982 218748
rect 53466 217948 53472 218000
rect 53524 217988 53530 218000
rect 273438 217988 273444 218000
rect 53524 217960 273444 217988
rect 53524 217948 53530 217960
rect 273438 217948 273444 217960
rect 273496 217948 273502 218000
rect 104158 217404 104164 217456
rect 104216 217444 104222 217456
rect 110414 217444 110420 217456
rect 104216 217416 110420 217444
rect 104216 217404 104222 217416
rect 110414 217404 110420 217416
rect 110472 217404 110478 217456
rect 125502 217268 125508 217320
rect 125560 217308 125566 217320
rect 171778 217308 171784 217320
rect 125560 217280 171784 217308
rect 125560 217268 125566 217280
rect 171778 217268 171784 217280
rect 171836 217268 171842 217320
rect 280890 217268 280896 217320
rect 280948 217308 280954 217320
rect 303614 217308 303620 217320
rect 280948 217280 303620 217308
rect 280948 217268 280954 217280
rect 303614 217268 303620 217280
rect 303672 217268 303678 217320
rect 73798 216588 73804 216640
rect 73856 216628 73862 216640
rect 74442 216628 74448 216640
rect 73856 216600 74448 216628
rect 73856 216588 73862 216600
rect 74442 216588 74448 216600
rect 74500 216628 74506 216640
rect 267734 216628 267740 216640
rect 74500 216600 267740 216628
rect 74500 216588 74506 216600
rect 267734 216588 267740 216600
rect 267792 216588 267798 216640
rect 110598 216520 110604 216572
rect 110656 216560 110662 216572
rect 242158 216560 242164 216572
rect 110656 216532 242164 216560
rect 110656 216520 110662 216532
rect 242158 216520 242164 216532
rect 242216 216520 242222 216572
rect 75914 215908 75920 215960
rect 75972 215948 75978 215960
rect 110598 215948 110604 215960
rect 75972 215920 110604 215948
rect 75972 215908 75978 215920
rect 110598 215908 110604 215920
rect 110656 215908 110662 215960
rect 249150 215908 249156 215960
rect 249208 215948 249214 215960
rect 338114 215948 338120 215960
rect 249208 215920 338120 215948
rect 249208 215908 249214 215920
rect 338114 215908 338120 215920
rect 338172 215908 338178 215960
rect 115750 215228 115756 215280
rect 115808 215268 115814 215280
rect 261018 215268 261024 215280
rect 115808 215240 261024 215268
rect 115808 215228 115814 215240
rect 261018 215228 261024 215240
rect 261076 215228 261082 215280
rect 117222 215160 117228 215212
rect 117280 215200 117286 215212
rect 241514 215200 241520 215212
rect 117280 215172 241520 215200
rect 117280 215160 117286 215172
rect 241514 215160 241520 215172
rect 241572 215200 241578 215212
rect 242158 215200 242164 215212
rect 241572 215172 242164 215200
rect 241572 215160 241578 215172
rect 242158 215160 242164 215172
rect 242216 215160 242222 215212
rect 88978 214616 88984 214668
rect 89036 214656 89042 214668
rect 114554 214656 114560 214668
rect 89036 214628 114560 214656
rect 89036 214616 89042 214628
rect 114554 214616 114560 214628
rect 114612 214656 114618 214668
rect 115750 214656 115756 214668
rect 114612 214628 115756 214656
rect 114612 214616 114618 214628
rect 115750 214616 115756 214628
rect 115808 214616 115814 214668
rect 84838 214548 84844 214600
rect 84896 214588 84902 214600
rect 116026 214588 116032 214600
rect 84896 214560 116032 214588
rect 84896 214548 84902 214560
rect 116026 214548 116032 214560
rect 116084 214588 116090 214600
rect 117222 214588 117228 214600
rect 116084 214560 117228 214588
rect 116084 214548 116090 214560
rect 117222 214548 117228 214560
rect 117280 214548 117286 214600
rect 3142 213936 3148 213988
rect 3200 213976 3206 213988
rect 3200 213948 6914 213976
rect 3200 213936 3206 213948
rect 6886 213908 6914 213948
rect 8202 213908 8208 213920
rect 6886 213880 8208 213908
rect 8202 213868 8208 213880
rect 8260 213908 8266 213920
rect 36538 213908 36544 213920
rect 8260 213880 36544 213908
rect 8260 213868 8266 213880
rect 36538 213868 36544 213880
rect 36596 213868 36602 213920
rect 243538 213908 243544 213920
rect 74506 213880 243544 213908
rect 66806 213800 66812 213852
rect 66864 213840 66870 213852
rect 67266 213840 67272 213852
rect 66864 213812 67272 213840
rect 66864 213800 66870 213812
rect 67266 213800 67272 213812
rect 67324 213840 67330 213852
rect 74506 213840 74534 213880
rect 243538 213868 243544 213880
rect 243596 213868 243602 213920
rect 67324 213812 74534 213840
rect 67324 213800 67330 213812
rect 139394 213800 139400 213852
rect 139452 213840 139458 213852
rect 200758 213840 200764 213852
rect 139452 213812 200764 213840
rect 139452 213800 139458 213812
rect 200758 213800 200764 213812
rect 200816 213800 200822 213852
rect 100662 213188 100668 213240
rect 100720 213228 100726 213240
rect 127250 213228 127256 213240
rect 100720 213200 127256 213228
rect 100720 213188 100726 213200
rect 127250 213188 127256 213200
rect 127308 213228 127314 213240
rect 139394 213228 139400 213240
rect 127308 213200 139400 213228
rect 127308 213188 127314 213200
rect 139394 213188 139400 213200
rect 139452 213188 139458 213240
rect 55122 212440 55128 212492
rect 55180 212480 55186 212492
rect 247678 212480 247684 212492
rect 55180 212452 247684 212480
rect 55180 212440 55186 212452
rect 247678 212440 247684 212452
rect 247736 212440 247742 212492
rect 128630 212372 128636 212424
rect 128688 212412 128694 212424
rect 250622 212412 250628 212424
rect 128688 212384 250628 212412
rect 128688 212372 128694 212384
rect 250622 212372 250628 212384
rect 250680 212372 250686 212424
rect 48038 211760 48044 211812
rect 48096 211800 48102 211812
rect 76650 211800 76656 211812
rect 48096 211772 76656 211800
rect 48096 211760 48102 211772
rect 76650 211760 76656 211772
rect 76708 211760 76714 211812
rect 88058 211760 88064 211812
rect 88116 211800 88122 211812
rect 116762 211800 116768 211812
rect 88116 211772 116768 211800
rect 88116 211760 88122 211772
rect 116762 211760 116768 211772
rect 116820 211760 116826 211812
rect 68462 211080 68468 211132
rect 68520 211120 68526 211132
rect 68922 211120 68928 211132
rect 68520 211092 68928 211120
rect 68520 211080 68526 211092
rect 68922 211080 68928 211092
rect 68980 211120 68986 211132
rect 253934 211120 253940 211132
rect 68980 211092 253940 211120
rect 68980 211080 68986 211092
rect 253934 211080 253940 211092
rect 253992 211080 253998 211132
rect 54938 211012 54944 211064
rect 54996 211052 55002 211064
rect 217318 211052 217324 211064
rect 54996 211024 217324 211052
rect 54996 211012 55002 211024
rect 217318 211012 217324 211024
rect 217376 211012 217382 211064
rect 92198 209108 92204 209160
rect 92256 209148 92262 209160
rect 118694 209148 118700 209160
rect 92256 209120 118700 209148
rect 92256 209108 92262 209120
rect 118694 209108 118700 209120
rect 118752 209148 118758 209160
rect 271874 209148 271880 209160
rect 118752 209120 271880 209148
rect 118752 209108 118758 209120
rect 271874 209108 271880 209120
rect 271932 209108 271938 209160
rect 80698 209040 80704 209092
rect 80756 209080 80762 209092
rect 103606 209080 103612 209092
rect 80756 209052 103612 209080
rect 80756 209040 80762 209052
rect 103606 209040 103612 209052
rect 103664 209080 103670 209092
rect 266446 209080 266452 209092
rect 103664 209052 266452 209080
rect 103664 209040 103670 209052
rect 266446 209040 266452 209052
rect 266504 209040 266510 209092
rect 61654 208292 61660 208344
rect 61712 208332 61718 208344
rect 236638 208332 236644 208344
rect 61712 208304 236644 208332
rect 61712 208292 61718 208304
rect 236638 208292 236644 208304
rect 236696 208292 236702 208344
rect 136634 208224 136640 208276
rect 136692 208264 136698 208276
rect 265250 208264 265256 208276
rect 136692 208236 265256 208264
rect 136692 208224 136698 208236
rect 265250 208224 265256 208236
rect 265308 208224 265314 208276
rect 96614 207612 96620 207664
rect 96672 207652 96678 207664
rect 128354 207652 128360 207664
rect 96672 207624 128360 207652
rect 96672 207612 96678 207624
rect 128354 207612 128360 207624
rect 128412 207652 128418 207664
rect 136634 207652 136640 207664
rect 128412 207624 136640 207652
rect 128412 207612 128418 207624
rect 136634 207612 136640 207624
rect 136692 207612 136698 207664
rect 56410 206932 56416 206984
rect 56468 206972 56474 206984
rect 207658 206972 207664 206984
rect 56468 206944 207664 206972
rect 56468 206932 56474 206944
rect 207658 206932 207664 206944
rect 207716 206932 207722 206984
rect 99190 206252 99196 206304
rect 99248 206292 99254 206304
rect 99248 206264 219434 206292
rect 99248 206252 99254 206264
rect 219406 206224 219434 206264
rect 240134 206224 240140 206236
rect 219406 206196 240140 206224
rect 240134 206184 240140 206196
rect 240192 206224 240198 206236
rect 240778 206224 240784 206236
rect 240192 206196 240784 206224
rect 240192 206184 240198 206196
rect 240778 206184 240784 206196
rect 240836 206184 240842 206236
rect 98730 205640 98736 205692
rect 98788 205680 98794 205692
rect 99190 205680 99196 205692
rect 98788 205652 99196 205680
rect 98788 205640 98794 205652
rect 99190 205640 99196 205652
rect 99248 205640 99254 205692
rect 61930 205572 61936 205624
rect 61988 205612 61994 205624
rect 229738 205612 229744 205624
rect 61988 205584 229744 205612
rect 61988 205572 61994 205584
rect 229738 205572 229744 205584
rect 229796 205572 229802 205624
rect 126974 205504 126980 205556
rect 127032 205544 127038 205556
rect 263594 205544 263600 205556
rect 127032 205516 263600 205544
rect 127032 205504 127038 205516
rect 263594 205504 263600 205516
rect 263652 205504 263658 205556
rect 91002 204892 91008 204944
rect 91060 204932 91066 204944
rect 106274 204932 106280 204944
rect 91060 204904 106280 204932
rect 91060 204892 91066 204904
rect 106274 204892 106280 204904
rect 106332 204932 106338 204944
rect 126974 204932 126980 204944
rect 106332 204904 126980 204932
rect 106332 204892 106338 204904
rect 126974 204892 126980 204904
rect 127032 204892 127038 204944
rect 102962 204212 102968 204264
rect 103020 204252 103026 204264
rect 103422 204252 103428 204264
rect 103020 204224 103428 204252
rect 103020 204212 103026 204224
rect 103422 204212 103428 204224
rect 103480 204252 103486 204264
rect 262398 204252 262404 204264
rect 103480 204224 262404 204252
rect 103480 204212 103486 204224
rect 262398 204212 262404 204224
rect 262456 204212 262462 204264
rect 82906 203532 82912 203584
rect 82964 203572 82970 203584
rect 105078 203572 105084 203584
rect 82964 203544 105084 203572
rect 82964 203532 82970 203544
rect 105078 203532 105084 203544
rect 105136 203532 105142 203584
rect 138658 202784 138664 202836
rect 138716 202824 138722 202836
rect 263778 202824 263784 202836
rect 138716 202796 263784 202824
rect 138716 202784 138722 202796
rect 263778 202784 263784 202796
rect 263836 202784 263842 202836
rect 3234 202104 3240 202156
rect 3292 202144 3298 202156
rect 124214 202144 124220 202156
rect 3292 202116 124220 202144
rect 3292 202104 3298 202116
rect 124214 202104 124220 202116
rect 124272 202104 124278 202156
rect 105630 202036 105636 202088
rect 105688 202076 105694 202088
rect 112162 202076 112168 202088
rect 105688 202048 112168 202076
rect 105688 202036 105694 202048
rect 112162 202036 112168 202048
rect 112220 202036 112226 202088
rect 128998 201492 129004 201544
rect 129056 201532 129062 201544
rect 132586 201532 132592 201544
rect 129056 201504 132592 201532
rect 129056 201492 129062 201504
rect 132586 201492 132592 201504
rect 132644 201492 132650 201544
rect 122190 201424 122196 201476
rect 122248 201464 122254 201476
rect 122742 201464 122748 201476
rect 122248 201436 122748 201464
rect 122248 201424 122254 201436
rect 122742 201424 122748 201436
rect 122800 201464 122806 201476
rect 271966 201464 271972 201476
rect 122800 201436 271972 201464
rect 122800 201424 122806 201436
rect 271966 201424 271972 201436
rect 272024 201424 272030 201476
rect 147030 200744 147036 200796
rect 147088 200784 147094 200796
rect 163498 200784 163504 200796
rect 147088 200756 163504 200784
rect 147088 200744 147094 200756
rect 163498 200744 163504 200756
rect 163556 200744 163562 200796
rect 82722 199520 82728 199572
rect 82780 199560 82786 199572
rect 90358 199560 90364 199572
rect 82780 199532 90364 199560
rect 82780 199520 82786 199532
rect 90358 199520 90364 199532
rect 90416 199520 90422 199572
rect 89806 199452 89812 199504
rect 89864 199492 89870 199504
rect 102962 199492 102968 199504
rect 89864 199464 102968 199492
rect 89864 199452 89870 199464
rect 102962 199452 102968 199464
rect 103020 199452 103026 199504
rect 56318 199384 56324 199436
rect 56376 199424 56382 199436
rect 80054 199424 80060 199436
rect 56376 199396 80060 199424
rect 56376 199384 56382 199396
rect 80054 199384 80060 199396
rect 80112 199384 80118 199436
rect 88150 199384 88156 199436
rect 88208 199424 88214 199436
rect 102134 199424 102140 199436
rect 88208 199396 102140 199424
rect 88208 199384 88214 199396
rect 102134 199384 102140 199396
rect 102192 199384 102198 199436
rect 50982 198636 50988 198688
rect 51040 198676 51046 198688
rect 249058 198676 249064 198688
rect 51040 198648 249064 198676
rect 51040 198636 51046 198648
rect 249058 198636 249064 198648
rect 249116 198636 249122 198688
rect 88150 197956 88156 198008
rect 88208 197996 88214 198008
rect 115382 197996 115388 198008
rect 88208 197968 115388 197996
rect 88208 197956 88214 197968
rect 115382 197956 115388 197968
rect 115440 197956 115446 198008
rect 46750 197276 46756 197328
rect 46808 197316 46814 197328
rect 276014 197316 276020 197328
rect 46808 197288 276020 197316
rect 46808 197276 46814 197288
rect 276014 197276 276020 197288
rect 276072 197276 276078 197328
rect 46198 196936 46204 196988
rect 46256 196976 46262 196988
rect 46750 196976 46756 196988
rect 46256 196948 46756 196976
rect 46256 196936 46262 196948
rect 46750 196936 46756 196948
rect 46808 196936 46814 196988
rect 59170 196596 59176 196648
rect 59228 196636 59234 196648
rect 77478 196636 77484 196648
rect 59228 196608 77484 196636
rect 59228 196596 59234 196608
rect 77478 196596 77484 196608
rect 77536 196596 77542 196648
rect 88058 196596 88064 196648
rect 88116 196636 88122 196648
rect 107838 196636 107844 196648
rect 88116 196608 107844 196636
rect 88116 196596 88122 196608
rect 107838 196596 107844 196608
rect 107896 196596 107902 196648
rect 116762 195916 116768 195968
rect 116820 195956 116826 195968
rect 269206 195956 269212 195968
rect 116820 195928 269212 195956
rect 116820 195916 116826 195928
rect 269206 195916 269212 195928
rect 269264 195916 269270 195968
rect 55030 194488 55036 194540
rect 55088 194528 55094 194540
rect 267826 194528 267832 194540
rect 55088 194500 267832 194528
rect 55088 194488 55094 194500
rect 267826 194488 267832 194500
rect 267884 194488 267890 194540
rect 37090 193808 37096 193860
rect 37148 193848 37154 193860
rect 68278 193848 68284 193860
rect 37148 193820 68284 193848
rect 37148 193808 37154 193820
rect 68278 193808 68284 193820
rect 68336 193808 68342 193860
rect 86770 193808 86776 193860
rect 86828 193848 86834 193860
rect 114646 193848 114652 193860
rect 86828 193820 114652 193848
rect 86828 193808 86834 193820
rect 114646 193808 114652 193820
rect 114704 193808 114710 193860
rect 313918 193128 313924 193180
rect 313976 193168 313982 193180
rect 580166 193168 580172 193180
rect 313976 193140 580172 193168
rect 313976 193128 313982 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 85574 191156 85580 191208
rect 85632 191196 85638 191208
rect 142154 191196 142160 191208
rect 85632 191168 142160 191196
rect 85632 191156 85638 191168
rect 142154 191156 142160 191168
rect 142212 191156 142218 191208
rect 1302 191088 1308 191140
rect 1360 191128 1366 191140
rect 157978 191128 157984 191140
rect 1360 191100 157984 191128
rect 1360 191088 1366 191100
rect 157978 191088 157984 191100
rect 158036 191088 158042 191140
rect 118602 189728 118608 189780
rect 118660 189768 118666 189780
rect 181438 189768 181444 189780
rect 118660 189740 181444 189768
rect 118660 189728 118666 189740
rect 181438 189728 181444 189740
rect 181496 189728 181502 189780
rect 2774 188844 2780 188896
rect 2832 188884 2838 188896
rect 4798 188884 4804 188896
rect 2832 188856 4804 188884
rect 2832 188844 2838 188856
rect 4798 188844 4804 188856
rect 4856 188844 4862 188896
rect 204898 185580 204904 185632
rect 204956 185620 204962 185632
rect 259546 185620 259552 185632
rect 204956 185592 259552 185620
rect 204956 185580 204962 185592
rect 259546 185580 259552 185592
rect 259604 185580 259610 185632
rect 37182 184152 37188 184204
rect 37240 184192 37246 184204
rect 151170 184192 151176 184204
rect 37240 184164 151176 184192
rect 37240 184152 37246 184164
rect 151170 184152 151176 184164
rect 151228 184152 151234 184204
rect 289078 184152 289084 184204
rect 289136 184192 289142 184204
rect 300854 184192 300860 184204
rect 289136 184164 300860 184192
rect 289136 184152 289142 184164
rect 300854 184152 300860 184164
rect 300912 184152 300918 184204
rect 2682 182792 2688 182844
rect 2740 182832 2746 182844
rect 166350 182832 166356 182844
rect 2740 182804 166356 182832
rect 2740 182792 2746 182804
rect 166350 182792 166356 182804
rect 166408 182792 166414 182844
rect 81526 180820 81532 180872
rect 81584 180860 81590 180872
rect 84838 180860 84844 180872
rect 81584 180832 84844 180860
rect 81584 180820 81590 180832
rect 84838 180820 84844 180832
rect 84896 180820 84902 180872
rect 5350 180072 5356 180124
rect 5408 180112 5414 180124
rect 156598 180112 156604 180124
rect 5408 180084 156604 180112
rect 5408 180072 5414 180084
rect 156598 180072 156604 180084
rect 156656 180072 156662 180124
rect 341518 179324 341524 179376
rect 341576 179364 341582 179376
rect 580166 179364 580172 179376
rect 341576 179336 580172 179364
rect 341576 179324 341582 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 28902 167628 28908 167680
rect 28960 167668 28966 167680
rect 184290 167668 184296 167680
rect 28960 167640 184296 167668
rect 28960 167628 28966 167640
rect 184290 167628 184296 167640
rect 184348 167628 184354 167680
rect 114462 164840 114468 164892
rect 114520 164880 114526 164892
rect 178770 164880 178776 164892
rect 114520 164852 178776 164880
rect 114520 164840 114526 164852
rect 178770 164840 178776 164852
rect 178828 164840 178834 164892
rect 20622 162120 20628 162172
rect 20680 162160 20686 162172
rect 187050 162160 187056 162172
rect 20680 162132 187056 162160
rect 20680 162120 20686 162132
rect 187050 162120 187056 162132
rect 187108 162120 187114 162172
rect 58986 160692 58992 160744
rect 59044 160732 59050 160744
rect 73798 160732 73804 160744
rect 59044 160704 73804 160732
rect 59044 160692 59050 160704
rect 73798 160692 73804 160704
rect 73856 160692 73862 160744
rect 66070 159332 66076 159384
rect 66128 159372 66134 159384
rect 273254 159372 273260 159384
rect 66128 159344 273260 159372
rect 66128 159332 66134 159344
rect 273254 159332 273260 159344
rect 273312 159332 273318 159384
rect 37090 157972 37096 158024
rect 37148 158012 37154 158024
rect 188430 158012 188436 158024
rect 37148 157984 188436 158012
rect 37148 157972 37154 157984
rect 188430 157972 188436 157984
rect 188488 157972 188494 158024
rect 84102 156680 84108 156732
rect 84160 156720 84166 156732
rect 102226 156720 102232 156732
rect 84160 156692 102232 156720
rect 84160 156680 84166 156692
rect 102226 156680 102232 156692
rect 102284 156680 102290 156732
rect 89070 156612 89076 156664
rect 89128 156652 89134 156664
rect 116578 156652 116584 156664
rect 89128 156624 116584 156652
rect 89128 156612 89134 156624
rect 116578 156612 116584 156624
rect 116636 156652 116642 156664
rect 316034 156652 316040 156664
rect 116636 156624 316040 156652
rect 116636 156612 116642 156624
rect 316034 156612 316040 156624
rect 316092 156612 316098 156664
rect 61746 155252 61752 155304
rect 61804 155292 61810 155304
rect 75178 155292 75184 155304
rect 61804 155264 75184 155292
rect 61804 155252 61810 155264
rect 75178 155252 75184 155264
rect 75236 155252 75242 155304
rect 43990 155184 43996 155236
rect 44048 155224 44054 155236
rect 180150 155224 180156 155236
rect 44048 155196 180156 155224
rect 44048 155184 44054 155196
rect 180150 155184 180156 155196
rect 180208 155184 180214 155236
rect 2958 149064 2964 149116
rect 3016 149104 3022 149116
rect 14458 149104 14464 149116
rect 3016 149076 14464 149104
rect 3016 149064 3022 149076
rect 14458 149064 14464 149076
rect 14516 149064 14522 149116
rect 313274 149104 313280 149116
rect 277366 149076 313280 149104
rect 63126 148996 63132 149048
rect 63184 149036 63190 149048
rect 276658 149036 276664 149048
rect 63184 149008 276664 149036
rect 63184 148996 63190 149008
rect 276658 148996 276664 149008
rect 276716 149036 276722 149048
rect 277366 149036 277394 149076
rect 313274 149064 313280 149076
rect 313332 149064 313338 149116
rect 276716 149008 277394 149036
rect 276716 148996 276722 149008
rect 39758 148316 39764 148368
rect 39816 148356 39822 148368
rect 73338 148356 73344 148368
rect 39816 148328 73344 148356
rect 39816 148316 39822 148328
rect 73338 148316 73344 148328
rect 73396 148316 73402 148368
rect 84562 147636 84568 147688
rect 84620 147676 84626 147688
rect 89070 147676 89076 147688
rect 84620 147648 89076 147676
rect 84620 147636 84626 147648
rect 89070 147636 89076 147648
rect 89128 147636 89134 147688
rect 76006 146072 76012 146124
rect 76064 146112 76070 146124
rect 79318 146112 79324 146124
rect 76064 146084 79324 146112
rect 76064 146072 76070 146084
rect 79318 146072 79324 146084
rect 79376 146072 79382 146124
rect 50798 145528 50804 145580
rect 50856 145568 50862 145580
rect 70486 145568 70492 145580
rect 50856 145540 70492 145568
rect 50856 145528 50862 145540
rect 70486 145528 70492 145540
rect 70544 145528 70550 145580
rect 84102 145528 84108 145580
rect 84160 145568 84166 145580
rect 116670 145568 116676 145580
rect 84160 145540 116676 145568
rect 84160 145528 84166 145540
rect 116670 145528 116676 145540
rect 116728 145528 116734 145580
rect 41230 144236 41236 144288
rect 41288 144276 41294 144288
rect 74810 144276 74816 144288
rect 41288 144248 74816 144276
rect 41288 144236 41294 144248
rect 74810 144236 74816 144248
rect 74868 144236 74874 144288
rect 53558 144168 53564 144220
rect 53616 144208 53622 144220
rect 170490 144208 170496 144220
rect 53616 144180 170496 144208
rect 53616 144168 53622 144180
rect 170490 144168 170496 144180
rect 170548 144168 170554 144220
rect 54846 142808 54852 142860
rect 54904 142848 54910 142860
rect 74534 142848 74540 142860
rect 54904 142820 74540 142848
rect 54904 142808 54910 142820
rect 74534 142808 74540 142820
rect 74592 142808 74598 142860
rect 85482 142808 85488 142860
rect 85540 142848 85546 142860
rect 94774 142848 94780 142860
rect 85540 142820 94780 142848
rect 85540 142808 85546 142820
rect 94774 142808 94780 142820
rect 94832 142808 94838 142860
rect 82814 142128 82820 142180
rect 82872 142168 82878 142180
rect 86218 142168 86224 142180
rect 82872 142140 86224 142168
rect 82872 142128 82878 142140
rect 86218 142128 86224 142140
rect 86276 142128 86282 142180
rect 88242 142128 88248 142180
rect 88300 142168 88306 142180
rect 100846 142168 100852 142180
rect 88300 142140 100852 142168
rect 88300 142128 88306 142140
rect 100846 142128 100852 142140
rect 100904 142128 100910 142180
rect 81342 141448 81348 141500
rect 81400 141488 81406 141500
rect 106366 141488 106372 141500
rect 81400 141460 106372 141488
rect 81400 141448 81406 141460
rect 106366 141448 106372 141460
rect 106424 141448 106430 141500
rect 3418 141380 3424 141432
rect 3476 141420 3482 141432
rect 88150 141420 88156 141432
rect 3476 141392 88156 141420
rect 3476 141380 3482 141392
rect 88150 141380 88156 141392
rect 88208 141380 88214 141432
rect 71682 140768 71688 140820
rect 71740 140808 71746 140820
rect 76558 140808 76564 140820
rect 71740 140780 76564 140808
rect 71740 140768 71746 140780
rect 76558 140768 76564 140780
rect 76616 140768 76622 140820
rect 106918 140768 106924 140820
rect 106976 140808 106982 140820
rect 114738 140808 114744 140820
rect 106976 140780 114744 140808
rect 106976 140768 106982 140780
rect 114738 140768 114744 140780
rect 114796 140768 114802 140820
rect 88150 140700 88156 140752
rect 88208 140740 88214 140752
rect 110506 140740 110512 140752
rect 88208 140712 110512 140740
rect 88208 140700 88214 140712
rect 110506 140700 110512 140712
rect 110564 140700 110570 140752
rect 56318 140088 56324 140140
rect 56376 140128 56382 140140
rect 78766 140128 78772 140140
rect 56376 140100 78772 140128
rect 56376 140088 56382 140100
rect 78766 140088 78772 140100
rect 78824 140088 78830 140140
rect 45370 140020 45376 140072
rect 45428 140060 45434 140072
rect 72326 140060 72332 140072
rect 45428 140032 72332 140060
rect 45428 140020 45434 140032
rect 72326 140020 72332 140032
rect 72384 140020 72390 140072
rect 91002 140020 91008 140072
rect 91060 140060 91066 140072
rect 102778 140060 102784 140072
rect 91060 140032 102784 140060
rect 91060 140020 91066 140032
rect 102778 140020 102784 140032
rect 102836 140020 102842 140072
rect 85482 139408 85488 139460
rect 85540 139448 85546 139460
rect 88978 139448 88984 139460
rect 85540 139420 88984 139448
rect 85540 139408 85546 139420
rect 88978 139408 88984 139420
rect 89036 139408 89042 139460
rect 14458 139340 14464 139392
rect 14516 139380 14522 139392
rect 88242 139380 88248 139392
rect 14516 139352 88248 139380
rect 14516 139340 14522 139352
rect 88242 139340 88248 139352
rect 88300 139340 88306 139392
rect 349798 139340 349804 139392
rect 349856 139380 349862 139392
rect 580166 139380 580172 139392
rect 349856 139352 580172 139380
rect 349856 139340 349862 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 94590 138728 94596 138780
rect 94648 138768 94654 138780
rect 113358 138768 113364 138780
rect 94648 138740 113364 138768
rect 94648 138728 94654 138740
rect 113358 138728 113364 138740
rect 113416 138728 113422 138780
rect 60366 138660 60372 138712
rect 60424 138700 60430 138712
rect 74626 138700 74632 138712
rect 60424 138672 74632 138700
rect 60424 138660 60430 138672
rect 74626 138660 74632 138672
rect 74684 138660 74690 138712
rect 79318 138660 79324 138712
rect 79376 138700 79382 138712
rect 111610 138700 111616 138712
rect 79376 138672 111616 138700
rect 79376 138660 79382 138672
rect 111610 138660 111616 138672
rect 111668 138700 111674 138712
rect 197998 138700 198004 138712
rect 111668 138672 198004 138700
rect 111668 138660 111674 138672
rect 197998 138660 198004 138672
rect 198056 138660 198062 138712
rect 75914 138048 75920 138100
rect 75972 138088 75978 138100
rect 76374 138088 76380 138100
rect 75972 138060 76380 138088
rect 75972 138048 75978 138060
rect 76374 138048 76380 138060
rect 76432 138048 76438 138100
rect 81434 138048 81440 138100
rect 81492 138088 81498 138100
rect 82078 138088 82084 138100
rect 81492 138060 82084 138088
rect 81492 138048 81498 138060
rect 82078 138048 82084 138060
rect 82136 138048 82142 138100
rect 89714 138048 89720 138100
rect 89772 138088 89778 138100
rect 90174 138088 90180 138100
rect 89772 138060 90180 138088
rect 89772 138048 89778 138060
rect 90174 138048 90180 138060
rect 90232 138048 90238 138100
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 39850 137952 39856 137964
rect 3292 137924 39856 137952
rect 3292 137912 3298 137924
rect 39850 137912 39856 137924
rect 39908 137912 39914 137964
rect 78490 137368 78496 137420
rect 78548 137408 78554 137420
rect 80422 137408 80428 137420
rect 78548 137380 80428 137408
rect 78548 137368 78554 137380
rect 80422 137368 80428 137380
rect 80480 137368 80486 137420
rect 88058 137300 88064 137352
rect 88116 137340 88122 137352
rect 102778 137340 102784 137352
rect 88116 137312 102784 137340
rect 88116 137300 88122 137312
rect 102778 137300 102784 137312
rect 102836 137300 102842 137352
rect 39850 137232 39856 137284
rect 39908 137272 39914 137284
rect 73154 137272 73160 137284
rect 39908 137244 73160 137272
rect 39908 137232 39914 137244
rect 73154 137232 73160 137244
rect 73212 137232 73218 137284
rect 79042 137232 79048 137284
rect 79100 137272 79106 137284
rect 86862 137272 86868 137284
rect 79100 137244 86868 137272
rect 79100 137232 79106 137244
rect 86862 137232 86868 137244
rect 86920 137232 86926 137284
rect 89070 137232 89076 137284
rect 89128 137272 89134 137284
rect 124858 137272 124864 137284
rect 89128 137244 124864 137272
rect 89128 137232 89134 137244
rect 124858 137232 124864 137244
rect 124916 137272 124922 137284
rect 170490 137272 170496 137284
rect 124916 137244 170496 137272
rect 124916 137232 124922 137244
rect 170490 137232 170496 137244
rect 170548 137232 170554 137284
rect 68278 136620 68284 136672
rect 68336 136660 68342 136672
rect 69934 136660 69940 136672
rect 68336 136632 69940 136660
rect 68336 136620 68342 136632
rect 69934 136620 69940 136632
rect 69992 136620 69998 136672
rect 74718 136620 74724 136672
rect 74776 136660 74782 136672
rect 76098 136660 76104 136672
rect 74776 136632 76104 136660
rect 74776 136620 74782 136632
rect 76098 136620 76104 136632
rect 76156 136620 76162 136672
rect 83642 136620 83648 136672
rect 83700 136660 83706 136672
rect 84102 136660 84108 136672
rect 83700 136632 84108 136660
rect 83700 136620 83706 136632
rect 84102 136620 84108 136632
rect 84160 136620 84166 136672
rect 85942 136620 85948 136672
rect 86000 136660 86006 136672
rect 88058 136660 88064 136672
rect 86000 136632 88064 136660
rect 86000 136620 86006 136632
rect 88058 136620 88064 136632
rect 88116 136620 88122 136672
rect 14458 135872 14464 135924
rect 14516 135912 14522 135924
rect 91002 135912 91008 135924
rect 14516 135884 91008 135912
rect 14516 135872 14522 135884
rect 91002 135872 91008 135884
rect 91060 135912 91066 135924
rect 91278 135912 91284 135924
rect 91060 135884 91284 135912
rect 91060 135872 91066 135884
rect 91278 135872 91284 135884
rect 91336 135872 91342 135924
rect 109126 135912 109132 135924
rect 99346 135884 109132 135912
rect 91186 135804 91192 135856
rect 91244 135844 91250 135856
rect 99346 135844 99374 135884
rect 109126 135872 109132 135884
rect 109184 135872 109190 135924
rect 91244 135816 99374 135844
rect 91244 135804 91250 135816
rect 44818 135260 44824 135312
rect 44876 135300 44882 135312
rect 91186 135300 91192 135312
rect 44876 135272 91192 135300
rect 44876 135260 44882 135272
rect 91186 135260 91192 135272
rect 91244 135260 91250 135312
rect 92290 135260 92296 135312
rect 92348 135300 92354 135312
rect 276014 135300 276020 135312
rect 92348 135272 276020 135300
rect 92348 135260 92354 135272
rect 276014 135260 276020 135272
rect 276072 135260 276078 135312
rect 35710 135192 35716 135244
rect 35768 135232 35774 135244
rect 66254 135232 66260 135244
rect 35768 135204 66260 135232
rect 35768 135192 35774 135204
rect 66254 135192 66260 135204
rect 66312 135192 66318 135244
rect 94774 135192 94780 135244
rect 94832 135232 94838 135244
rect 99374 135232 99380 135244
rect 94832 135204 99380 135232
rect 94832 135192 94838 135204
rect 99374 135192 99380 135204
rect 99432 135192 99438 135244
rect 40862 135124 40868 135176
rect 40920 135164 40926 135176
rect 41322 135164 41328 135176
rect 40920 135136 41328 135164
rect 40920 135124 40926 135136
rect 41322 135124 41328 135136
rect 41380 135164 41386 135176
rect 75454 135164 75460 135176
rect 41380 135136 75460 135164
rect 41380 135124 41386 135136
rect 75454 135124 75460 135136
rect 75512 135124 75518 135176
rect 68646 134784 68652 134836
rect 68704 134824 68710 134836
rect 69658 134824 69664 134836
rect 68704 134796 69664 134824
rect 68704 134784 68710 134796
rect 69658 134784 69664 134796
rect 69716 134784 69722 134836
rect 89254 134784 89260 134836
rect 89312 134784 89318 134836
rect 90358 134784 90364 134836
rect 90416 134824 90422 134836
rect 96062 134824 96068 134836
rect 90416 134796 96068 134824
rect 90416 134784 90422 134796
rect 96062 134784 96068 134796
rect 96120 134784 96126 134836
rect 89272 134756 89300 134784
rect 94866 134756 94872 134768
rect 89272 134728 94872 134756
rect 94866 134716 94872 134728
rect 94924 134716 94930 134768
rect 70486 134580 70492 134632
rect 70544 134620 70550 134632
rect 71222 134620 71228 134632
rect 70544 134592 71228 134620
rect 70544 134580 70550 134592
rect 71222 134580 71228 134592
rect 71280 134580 71286 134632
rect 3418 134512 3424 134564
rect 3476 134552 3482 134564
rect 40862 134552 40868 134564
rect 3476 134524 40868 134552
rect 3476 134512 3482 134524
rect 40862 134512 40868 134524
rect 40920 134512 40926 134564
rect 47854 133832 47860 133884
rect 47912 133872 47918 133884
rect 66254 133872 66260 133884
rect 47912 133844 66260 133872
rect 47912 133832 47918 133844
rect 66254 133832 66260 133844
rect 66312 133832 66318 133884
rect 96706 133832 96712 133884
rect 96764 133872 96770 133884
rect 122190 133872 122196 133884
rect 96764 133844 122196 133872
rect 96764 133832 96770 133844
rect 122190 133832 122196 133844
rect 122248 133832 122254 133884
rect 94958 133152 94964 133204
rect 95016 133192 95022 133204
rect 267826 133192 267832 133204
rect 95016 133164 267832 133192
rect 95016 133152 95022 133164
rect 267826 133152 267832 133164
rect 267884 133152 267890 133204
rect 44082 132404 44088 132456
rect 44140 132444 44146 132456
rect 66254 132444 66260 132456
rect 44140 132416 66260 132444
rect 44140 132404 44146 132416
rect 66254 132404 66260 132416
rect 66312 132404 66318 132456
rect 96614 132404 96620 132456
rect 96672 132444 96678 132456
rect 131758 132444 131764 132456
rect 96672 132416 131764 132444
rect 96672 132404 96678 132416
rect 131758 132404 131764 132416
rect 131816 132404 131822 132456
rect 53650 132336 53656 132388
rect 53708 132376 53714 132388
rect 66346 132376 66352 132388
rect 53708 132348 66352 132376
rect 53708 132336 53714 132348
rect 66346 132336 66352 132348
rect 66404 132336 66410 132388
rect 96706 129684 96712 129736
rect 96764 129724 96770 129736
rect 131206 129724 131212 129736
rect 96764 129696 131212 129724
rect 96764 129684 96770 129696
rect 131206 129684 131212 129696
rect 131264 129684 131270 129736
rect 97258 129616 97264 129668
rect 97316 129656 97322 129668
rect 127158 129656 127164 129668
rect 97316 129628 127164 129656
rect 97316 129616 97322 129628
rect 127158 129616 127164 129628
rect 127216 129616 127222 129668
rect 57882 129004 57888 129056
rect 57940 129044 57946 129056
rect 66438 129044 66444 129056
rect 57940 129016 66444 129044
rect 57940 129004 57946 129016
rect 66438 129004 66444 129016
rect 66496 129004 66502 129056
rect 32858 128256 32864 128308
rect 32916 128296 32922 128308
rect 66898 128296 66904 128308
rect 32916 128268 66904 128296
rect 32916 128256 32922 128268
rect 66898 128256 66904 128268
rect 66956 128256 66962 128308
rect 97534 128256 97540 128308
rect 97592 128296 97598 128308
rect 134702 128296 134708 128308
rect 97592 128268 134708 128296
rect 97592 128256 97598 128268
rect 134702 128256 134708 128268
rect 134760 128256 134766 128308
rect 59078 128188 59084 128240
rect 59136 128228 59142 128240
rect 66714 128228 66720 128240
rect 59136 128200 66720 128228
rect 59136 128188 59142 128200
rect 66714 128188 66720 128200
rect 66772 128188 66778 128240
rect 97166 128188 97172 128240
rect 97224 128228 97230 128240
rect 100846 128228 100852 128240
rect 97224 128200 100852 128228
rect 97224 128188 97230 128200
rect 100846 128188 100852 128200
rect 100904 128188 100910 128240
rect 97810 126896 97816 126948
rect 97868 126936 97874 126948
rect 135254 126936 135260 126948
rect 97868 126908 135260 126936
rect 97868 126896 97874 126908
rect 135254 126896 135260 126908
rect 135312 126896 135318 126948
rect 43898 126216 43904 126268
rect 43956 126256 43962 126268
rect 66898 126256 66904 126268
rect 43956 126228 66904 126256
rect 43956 126216 43962 126228
rect 66898 126216 66904 126228
rect 66956 126216 66962 126268
rect 101490 126216 101496 126268
rect 101548 126256 101554 126268
rect 106458 126256 106464 126268
rect 101548 126228 106464 126256
rect 101548 126216 101554 126228
rect 106458 126216 106464 126228
rect 106516 126216 106522 126268
rect 57790 125536 57796 125588
rect 57848 125576 57854 125588
rect 66254 125576 66260 125588
rect 57848 125548 66260 125576
rect 57848 125536 57854 125548
rect 66254 125536 66260 125548
rect 66312 125536 66318 125588
rect 97442 125536 97448 125588
rect 97500 125576 97506 125588
rect 122834 125576 122840 125588
rect 97500 125548 122840 125576
rect 97500 125536 97506 125548
rect 122834 125536 122840 125548
rect 122892 125536 122898 125588
rect 96798 124856 96804 124908
rect 96856 124896 96862 124908
rect 128446 124896 128452 124908
rect 96856 124868 128452 124896
rect 96856 124856 96862 124868
rect 128446 124856 128452 124868
rect 128504 124856 128510 124908
rect 59262 124108 59268 124160
rect 59320 124148 59326 124160
rect 63218 124148 63224 124160
rect 59320 124120 63224 124148
rect 59320 124108 59326 124120
rect 63218 124108 63224 124120
rect 63276 124108 63282 124160
rect 94682 124108 94688 124160
rect 94740 124148 94746 124160
rect 95142 124148 95148 124160
rect 94740 124120 95148 124148
rect 94740 124108 94746 124120
rect 95142 124108 95148 124120
rect 95200 124108 95206 124160
rect 97810 124108 97816 124160
rect 97868 124148 97874 124160
rect 130378 124148 130384 124160
rect 97868 124120 130384 124148
rect 97868 124108 97874 124120
rect 130378 124108 130384 124120
rect 130436 124148 130442 124160
rect 130562 124148 130568 124160
rect 130436 124120 130568 124148
rect 130436 124108 130442 124120
rect 130562 124108 130568 124120
rect 130620 124108 130626 124160
rect 96614 123972 96620 124024
rect 96672 124012 96678 124024
rect 98730 124012 98736 124024
rect 96672 123984 98736 124012
rect 96672 123972 96678 123984
rect 98730 123972 98736 123984
rect 98788 123972 98794 124024
rect 130562 123428 130568 123480
rect 130620 123468 130626 123480
rect 173250 123468 173256 123480
rect 130620 123440 173256 123468
rect 130620 123428 130626 123440
rect 173250 123428 173256 123440
rect 173308 123428 173314 123480
rect 63218 122884 63224 122936
rect 63276 122924 63282 122936
rect 66898 122924 66904 122936
rect 63276 122896 66904 122924
rect 63276 122884 63282 122896
rect 66898 122884 66904 122896
rect 66956 122884 66962 122936
rect 53374 122748 53380 122800
rect 53432 122788 53438 122800
rect 66898 122788 66904 122800
rect 53432 122760 66904 122788
rect 53432 122748 53438 122760
rect 66898 122748 66904 122760
rect 66956 122748 66962 122800
rect 97810 122748 97816 122800
rect 97868 122788 97874 122800
rect 135898 122788 135904 122800
rect 97868 122760 135904 122788
rect 97868 122748 97874 122760
rect 135898 122748 135904 122760
rect 135956 122748 135962 122800
rect 61654 122680 61660 122732
rect 61712 122720 61718 122732
rect 66714 122720 66720 122732
rect 61712 122692 66720 122720
rect 61712 122680 61718 122692
rect 66714 122680 66720 122692
rect 66772 122680 66778 122732
rect 96062 122272 96068 122324
rect 96120 122312 96126 122324
rect 97994 122312 98000 122324
rect 96120 122284 98000 122312
rect 96120 122272 96126 122284
rect 97994 122272 98000 122284
rect 98052 122272 98058 122324
rect 135898 122068 135904 122120
rect 135956 122108 135962 122120
rect 356054 122108 356060 122120
rect 135956 122080 356060 122108
rect 135956 122068 135962 122080
rect 356054 122068 356060 122080
rect 356112 122068 356118 122120
rect 32950 121388 32956 121440
rect 33008 121428 33014 121440
rect 65518 121428 65524 121440
rect 33008 121400 65524 121428
rect 33008 121388 33014 121400
rect 65518 121388 65524 121400
rect 65576 121388 65582 121440
rect 97810 121388 97816 121440
rect 97868 121428 97874 121440
rect 113266 121428 113272 121440
rect 97868 121400 113272 121428
rect 97868 121388 97874 121400
rect 113266 121388 113272 121400
rect 113324 121388 113330 121440
rect 60550 120164 60556 120216
rect 60608 120204 60614 120216
rect 66254 120204 66260 120216
rect 60608 120176 66260 120204
rect 60608 120164 60614 120176
rect 66254 120164 66260 120176
rect 66312 120164 66318 120216
rect 97810 120164 97816 120216
rect 97868 120204 97874 120216
rect 104894 120204 104900 120216
rect 97868 120176 104900 120204
rect 97868 120164 97874 120176
rect 104894 120164 104900 120176
rect 104952 120164 104958 120216
rect 54938 120028 54944 120080
rect 54996 120068 55002 120080
rect 66898 120068 66904 120080
rect 54996 120040 66904 120068
rect 54996 120028 55002 120040
rect 66898 120028 66904 120040
rect 66956 120028 66962 120080
rect 123570 119348 123576 119400
rect 123628 119388 123634 119400
rect 159450 119388 159456 119400
rect 123628 119360 159456 119388
rect 123628 119348 123634 119360
rect 159450 119348 159456 119360
rect 159508 119348 159514 119400
rect 97810 118600 97816 118652
rect 97868 118640 97874 118652
rect 122926 118640 122932 118652
rect 97868 118612 122932 118640
rect 97868 118600 97874 118612
rect 122926 118600 122932 118612
rect 122984 118600 122990 118652
rect 41138 118532 41144 118584
rect 41196 118572 41202 118584
rect 66898 118572 66904 118584
rect 41196 118544 66904 118572
rect 41196 118532 41202 118544
rect 66898 118532 66904 118544
rect 66956 118532 66962 118584
rect 50890 117240 50896 117292
rect 50948 117280 50954 117292
rect 66898 117280 66904 117292
rect 50948 117252 66904 117280
rect 50948 117240 50954 117252
rect 66898 117240 66904 117252
rect 66956 117240 66962 117292
rect 97810 117240 97816 117292
rect 97868 117280 97874 117292
rect 120074 117280 120080 117292
rect 97868 117252 120080 117280
rect 97868 117240 97874 117252
rect 120074 117240 120080 117252
rect 120132 117240 120138 117292
rect 96614 117036 96620 117088
rect 96672 117076 96678 117088
rect 98638 117076 98644 117088
rect 96672 117048 98644 117076
rect 96672 117036 96678 117048
rect 98638 117036 98644 117048
rect 98696 117036 98702 117088
rect 100018 116288 100024 116340
rect 100076 116328 100082 116340
rect 104986 116328 104992 116340
rect 100076 116300 104992 116328
rect 100076 116288 100082 116300
rect 104986 116288 104992 116300
rect 105044 116288 105050 116340
rect 47946 115880 47952 115932
rect 48004 115920 48010 115932
rect 66898 115920 66904 115932
rect 48004 115892 66904 115920
rect 48004 115880 48010 115892
rect 66898 115880 66904 115892
rect 66956 115880 66962 115932
rect 97718 115880 97724 115932
rect 97776 115920 97782 115932
rect 133138 115920 133144 115932
rect 97776 115892 133144 115920
rect 97776 115880 97782 115892
rect 133138 115880 133144 115892
rect 133196 115920 133202 115932
rect 133782 115920 133788 115932
rect 133196 115892 133788 115920
rect 133196 115880 133202 115892
rect 133782 115880 133788 115892
rect 133840 115880 133846 115932
rect 97810 115812 97816 115864
rect 97868 115852 97874 115864
rect 118786 115852 118792 115864
rect 97868 115824 118792 115852
rect 97868 115812 97874 115824
rect 118786 115812 118792 115824
rect 118844 115812 118850 115864
rect 133782 115200 133788 115252
rect 133840 115240 133846 115252
rect 187050 115240 187056 115252
rect 133840 115212 187056 115240
rect 133840 115200 133846 115212
rect 187050 115200 187056 115212
rect 187108 115200 187114 115252
rect 60642 114588 60648 114640
rect 60700 114628 60706 114640
rect 67174 114628 67180 114640
rect 60700 114600 67180 114628
rect 60700 114588 60706 114600
rect 67174 114588 67180 114600
rect 67232 114588 67238 114640
rect 8202 114452 8208 114504
rect 8260 114492 8266 114504
rect 66622 114492 66628 114504
rect 8260 114464 66628 114492
rect 8260 114452 8266 114464
rect 66622 114452 66628 114464
rect 66680 114452 66686 114504
rect 63494 114384 63500 114436
rect 63552 114424 63558 114436
rect 64598 114424 64604 114436
rect 63552 114396 64604 114424
rect 63552 114384 63558 114396
rect 64598 114384 64604 114396
rect 64656 114384 64662 114436
rect 96614 113840 96620 113892
rect 96672 113880 96678 113892
rect 109218 113880 109224 113892
rect 96672 113852 109224 113880
rect 96672 113840 96678 113852
rect 109218 113840 109224 113852
rect 109276 113840 109282 113892
rect 102778 113772 102784 113824
rect 102836 113812 102842 113824
rect 255314 113812 255320 113824
rect 102836 113784 255320 113812
rect 102836 113772 102842 113784
rect 255314 113772 255320 113784
rect 255372 113772 255378 113824
rect 34330 113092 34336 113144
rect 34388 113132 34394 113144
rect 66898 113132 66904 113144
rect 34388 113104 66904 113132
rect 34388 113092 34394 113104
rect 66898 113092 66904 113104
rect 66956 113092 66962 113144
rect 97810 113092 97816 113144
rect 97868 113132 97874 113144
rect 129734 113132 129740 113144
rect 97868 113104 129740 113132
rect 97868 113092 97874 113104
rect 129734 113092 129740 113104
rect 129792 113092 129798 113144
rect 102134 112412 102140 112464
rect 102192 112452 102198 112464
rect 125686 112452 125692 112464
rect 102192 112424 125692 112452
rect 102192 112412 102198 112424
rect 125686 112412 125692 112424
rect 125744 112412 125750 112464
rect 169110 112412 169116 112464
rect 169168 112452 169174 112464
rect 264238 112452 264244 112464
rect 169168 112424 264244 112452
rect 169168 112412 169174 112424
rect 264238 112412 264244 112424
rect 264296 112412 264302 112464
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 44818 111772 44824 111784
rect 3200 111744 44824 111772
rect 3200 111732 3206 111744
rect 44818 111732 44824 111744
rect 44876 111732 44882 111784
rect 56410 111732 56416 111784
rect 56468 111772 56474 111784
rect 66898 111772 66904 111784
rect 56468 111744 66904 111772
rect 56468 111732 56474 111744
rect 66898 111732 66904 111744
rect 66956 111732 66962 111784
rect 97902 111732 97908 111784
rect 97960 111772 97966 111784
rect 136726 111772 136732 111784
rect 97960 111744 136732 111772
rect 97960 111732 97966 111744
rect 136726 111732 136732 111744
rect 136784 111732 136790 111784
rect 101398 110984 101404 111036
rect 101456 111024 101462 111036
rect 104894 111024 104900 111036
rect 101456 110996 104900 111024
rect 101456 110984 101462 110996
rect 104894 110984 104900 110996
rect 104952 110984 104958 111036
rect 46750 110372 46756 110424
rect 46808 110412 46814 110424
rect 66898 110412 66904 110424
rect 46808 110384 66904 110412
rect 46808 110372 46814 110384
rect 66898 110372 66904 110384
rect 66956 110372 66962 110424
rect 97810 110372 97816 110424
rect 97868 110412 97874 110424
rect 133230 110412 133236 110424
rect 97868 110384 133236 110412
rect 97868 110372 97874 110384
rect 133230 110372 133236 110384
rect 133288 110372 133294 110424
rect 97902 110304 97908 110356
rect 97960 110344 97966 110356
rect 127066 110344 127072 110356
rect 97960 110316 127072 110344
rect 97960 110304 97966 110316
rect 127066 110304 127072 110316
rect 127124 110304 127130 110356
rect 45462 109692 45468 109744
rect 45520 109732 45526 109744
rect 57054 109732 57060 109744
rect 45520 109704 57060 109732
rect 45520 109692 45526 109704
rect 57054 109692 57060 109704
rect 57112 109692 57118 109744
rect 127066 109692 127072 109744
rect 127124 109732 127130 109744
rect 273898 109732 273904 109744
rect 127124 109704 273904 109732
rect 127124 109692 127130 109704
rect 273898 109692 273904 109704
rect 273956 109692 273962 109744
rect 56594 109012 56600 109064
rect 56652 109052 56658 109064
rect 57054 109052 57060 109064
rect 56652 109024 57060 109052
rect 56652 109012 56658 109024
rect 57054 109012 57060 109024
rect 57112 109052 57118 109064
rect 66254 109052 66260 109064
rect 57112 109024 66260 109052
rect 57112 109012 57118 109024
rect 66254 109012 66260 109024
rect 66312 109012 66318 109064
rect 52178 108944 52184 108996
rect 52236 108984 52242 108996
rect 66990 108984 66996 108996
rect 52236 108956 66996 108984
rect 52236 108944 52242 108956
rect 66990 108944 66996 108956
rect 67048 108944 67054 108996
rect 97902 108944 97908 108996
rect 97960 108984 97966 108996
rect 113174 108984 113180 108996
rect 97960 108956 113180 108984
rect 97960 108944 97966 108956
rect 113174 108944 113180 108956
rect 113232 108944 113238 108996
rect 57606 108876 57612 108928
rect 57664 108916 57670 108928
rect 66898 108916 66904 108928
rect 57664 108888 66904 108916
rect 57664 108876 57670 108888
rect 66898 108876 66904 108888
rect 66956 108876 66962 108928
rect 97718 108876 97724 108928
rect 97776 108916 97782 108928
rect 111978 108916 111984 108928
rect 97776 108888 111984 108916
rect 97776 108876 97782 108888
rect 111978 108876 111984 108888
rect 112036 108876 112042 108928
rect 41414 107584 41420 107636
rect 41472 107624 41478 107636
rect 42702 107624 42708 107636
rect 41472 107596 42708 107624
rect 41472 107584 41478 107596
rect 42702 107584 42708 107596
rect 42760 107624 42766 107636
rect 66898 107624 66904 107636
rect 42760 107596 66904 107624
rect 42760 107584 42766 107596
rect 66898 107584 66904 107596
rect 66956 107584 66962 107636
rect 49602 107516 49608 107568
rect 49660 107556 49666 107568
rect 66714 107556 66720 107568
rect 49660 107528 66720 107556
rect 49660 107516 49666 107528
rect 66714 107516 66720 107528
rect 66772 107516 66778 107568
rect 97534 107312 97540 107364
rect 97592 107352 97598 107364
rect 102134 107352 102140 107364
rect 97592 107324 102140 107352
rect 97592 107312 97598 107324
rect 102134 107312 102140 107324
rect 102192 107312 102198 107364
rect 7558 106904 7564 106956
rect 7616 106944 7622 106956
rect 41414 106944 41420 106956
rect 7616 106916 41420 106944
rect 7616 106904 7622 106916
rect 41414 106904 41420 106916
rect 41472 106904 41478 106956
rect 103422 106904 103428 106956
rect 103480 106944 103486 106956
rect 182818 106944 182824 106956
rect 103480 106916 182824 106944
rect 103480 106904 103486 106916
rect 182818 106904 182824 106916
rect 182876 106904 182882 106956
rect 49510 106224 49516 106276
rect 49568 106264 49574 106276
rect 66898 106264 66904 106276
rect 49568 106236 66904 106264
rect 49568 106224 49574 106236
rect 66898 106224 66904 106236
rect 66956 106224 66962 106276
rect 97626 106224 97632 106276
rect 97684 106264 97690 106276
rect 125778 106264 125784 106276
rect 97684 106236 125784 106264
rect 97684 106224 97690 106236
rect 125778 106224 125784 106236
rect 125836 106224 125842 106276
rect 97902 105544 97908 105596
rect 97960 105584 97966 105596
rect 180150 105584 180156 105596
rect 97960 105556 180156 105584
rect 97960 105544 97966 105556
rect 180150 105544 180156 105556
rect 180208 105544 180214 105596
rect 60458 104796 60464 104848
rect 60516 104836 60522 104848
rect 66254 104836 66260 104848
rect 60516 104808 66260 104836
rect 60516 104796 60522 104808
rect 66254 104796 66260 104808
rect 66312 104796 66318 104848
rect 97166 104796 97172 104848
rect 97224 104836 97230 104848
rect 107746 104836 107752 104848
rect 97224 104808 107752 104836
rect 97224 104796 97230 104808
rect 107746 104796 107752 104808
rect 107804 104796 107810 104848
rect 94774 104728 94780 104780
rect 94832 104768 94838 104780
rect 102318 104768 102324 104780
rect 94832 104740 102324 104768
rect 94832 104728 94838 104740
rect 102318 104728 102324 104740
rect 102376 104728 102382 104780
rect 61930 103436 61936 103488
rect 61988 103476 61994 103488
rect 66898 103476 66904 103488
rect 61988 103448 66904 103476
rect 61988 103436 61994 103448
rect 66898 103436 66904 103448
rect 66956 103436 66962 103488
rect 97166 103436 97172 103488
rect 97224 103476 97230 103488
rect 135346 103476 135352 103488
rect 97224 103448 135352 103476
rect 97224 103436 97230 103448
rect 135346 103436 135352 103448
rect 135404 103436 135410 103488
rect 97718 102756 97724 102808
rect 97776 102796 97782 102808
rect 120166 102796 120172 102808
rect 97776 102768 120172 102796
rect 97776 102756 97782 102768
rect 120166 102756 120172 102768
rect 120224 102756 120230 102808
rect 135346 102756 135352 102808
rect 135404 102796 135410 102808
rect 184290 102796 184296 102808
rect 135404 102768 184296 102796
rect 135404 102756 135410 102768
rect 184290 102756 184296 102768
rect 184348 102756 184354 102808
rect 64690 102076 64696 102128
rect 64748 102116 64754 102128
rect 66438 102116 66444 102128
rect 64748 102088 66444 102116
rect 64748 102076 64754 102088
rect 66438 102076 66444 102088
rect 66496 102076 66502 102128
rect 97902 102076 97908 102128
rect 97960 102116 97966 102128
rect 131298 102116 131304 102128
rect 97960 102088 131304 102116
rect 97960 102076 97966 102088
rect 131298 102076 131304 102088
rect 131356 102076 131362 102128
rect 97810 102008 97816 102060
rect 97868 102048 97874 102060
rect 124214 102048 124220 102060
rect 97868 102020 124220 102048
rect 97868 102008 97874 102020
rect 124214 102008 124220 102020
rect 124272 102008 124278 102060
rect 46842 101396 46848 101448
rect 46900 101436 46906 101448
rect 60734 101436 60740 101448
rect 46900 101408 60740 101436
rect 46900 101396 46906 101408
rect 60734 101396 60740 101408
rect 60792 101436 60798 101448
rect 66806 101436 66812 101448
rect 60792 101408 66812 101436
rect 60792 101396 60798 101408
rect 66806 101396 66812 101408
rect 66864 101396 66870 101448
rect 131298 101396 131304 101448
rect 131356 101436 131362 101448
rect 233142 101436 233148 101448
rect 131356 101408 233148 101436
rect 131356 101396 131362 101408
rect 233142 101396 233148 101408
rect 233200 101396 233206 101448
rect 61562 100648 61568 100700
rect 61620 100688 61626 100700
rect 66806 100688 66812 100700
rect 61620 100660 66812 100688
rect 61620 100648 61626 100660
rect 66806 100648 66812 100660
rect 66864 100648 66870 100700
rect 97902 100648 97908 100700
rect 97960 100688 97966 100700
rect 130194 100688 130200 100700
rect 97960 100660 130200 100688
rect 97960 100648 97966 100660
rect 130194 100648 130200 100660
rect 130252 100648 130258 100700
rect 130194 99968 130200 100020
rect 130252 100008 130258 100020
rect 131022 100008 131028 100020
rect 130252 99980 131028 100008
rect 130252 99968 130258 99980
rect 131022 99968 131028 99980
rect 131080 100008 131086 100020
rect 151170 100008 151176 100020
rect 131080 99980 151176 100008
rect 131080 99968 131086 99980
rect 151170 99968 151176 99980
rect 151228 99968 151234 100020
rect 168282 99968 168288 100020
rect 168340 100008 168346 100020
rect 198090 100008 198096 100020
rect 168340 99980 198096 100008
rect 168340 99968 168346 99980
rect 198090 99968 198096 99980
rect 198148 99968 198154 100020
rect 56502 99492 56508 99544
rect 56560 99532 56566 99544
rect 63402 99532 63408 99544
rect 56560 99504 63408 99532
rect 56560 99492 56566 99504
rect 63402 99492 63408 99504
rect 63460 99532 63466 99544
rect 66806 99532 66812 99544
rect 63460 99504 66812 99532
rect 63460 99492 63466 99504
rect 66806 99492 66812 99504
rect 66864 99492 66870 99544
rect 53466 99288 53472 99340
rect 53524 99328 53530 99340
rect 66806 99328 66812 99340
rect 53524 99300 66812 99328
rect 53524 99288 53530 99300
rect 66806 99288 66812 99300
rect 66864 99288 66870 99340
rect 97534 99288 97540 99340
rect 97592 99328 97598 99340
rect 134610 99328 134616 99340
rect 97592 99300 134616 99328
rect 97592 99288 97598 99300
rect 134610 99288 134616 99300
rect 134668 99328 134674 99340
rect 135162 99328 135168 99340
rect 134668 99300 135168 99328
rect 134668 99288 134674 99300
rect 135162 99288 135168 99300
rect 135220 99288 135226 99340
rect 135162 98608 135168 98660
rect 135220 98648 135226 98660
rect 220078 98648 220084 98660
rect 135220 98620 220084 98648
rect 135220 98608 135226 98620
rect 220078 98608 220084 98620
rect 220136 98608 220142 98660
rect 97902 97928 97908 97980
rect 97960 97968 97966 97980
rect 111886 97968 111892 97980
rect 97960 97940 111892 97968
rect 97960 97928 97966 97940
rect 111886 97928 111892 97940
rect 111944 97928 111950 97980
rect 97534 97860 97540 97912
rect 97592 97900 97598 97912
rect 106918 97900 106924 97912
rect 97592 97872 106924 97900
rect 97592 97860 97598 97872
rect 106918 97860 106924 97872
rect 106976 97860 106982 97912
rect 55122 97248 55128 97300
rect 55180 97288 55186 97300
rect 66806 97288 66812 97300
rect 55180 97260 66812 97288
rect 55180 97248 55186 97260
rect 66806 97248 66812 97260
rect 66864 97248 66870 97300
rect 3050 96636 3056 96688
rect 3108 96676 3114 96688
rect 65610 96676 65616 96688
rect 3108 96648 65616 96676
rect 3108 96636 3114 96648
rect 65610 96636 65616 96648
rect 65668 96636 65674 96688
rect 42610 96568 42616 96620
rect 42668 96608 42674 96620
rect 66254 96608 66260 96620
rect 42668 96580 66260 96608
rect 42668 96568 42674 96580
rect 66254 96568 66260 96580
rect 66312 96568 66318 96620
rect 97902 95956 97908 96008
rect 97960 95996 97966 96008
rect 99282 95996 99288 96008
rect 97960 95968 99288 95996
rect 97960 95956 97966 95968
rect 99282 95956 99288 95968
rect 99340 95996 99346 96008
rect 178770 95996 178776 96008
rect 99340 95968 178776 95996
rect 99340 95956 99346 95968
rect 178770 95956 178776 95968
rect 178828 95956 178834 96008
rect 175182 95888 175188 95940
rect 175240 95928 175246 95940
rect 276106 95928 276112 95940
rect 175240 95900 276112 95928
rect 175240 95888 175246 95900
rect 276106 95888 276112 95900
rect 276164 95888 276170 95940
rect 55030 95140 55036 95192
rect 55088 95180 55094 95192
rect 66438 95180 66444 95192
rect 55088 95152 66444 95180
rect 55088 95140 55094 95152
rect 66438 95140 66444 95152
rect 66496 95140 66502 95192
rect 97902 95140 97908 95192
rect 97960 95180 97966 95192
rect 110414 95180 110420 95192
rect 97960 95152 110420 95180
rect 97960 95140 97966 95152
rect 110414 95140 110420 95152
rect 110472 95140 110478 95192
rect 64782 93780 64788 93832
rect 64840 93820 64846 93832
rect 66806 93820 66812 93832
rect 64840 93792 66812 93820
rect 64840 93780 64846 93792
rect 66806 93780 66812 93792
rect 66864 93780 66870 93832
rect 97902 93780 97908 93832
rect 97960 93820 97966 93832
rect 128354 93820 128360 93832
rect 97960 93792 128360 93820
rect 97960 93780 97966 93792
rect 128354 93780 128360 93792
rect 128412 93780 128418 93832
rect 94682 93508 94688 93560
rect 94740 93548 94746 93560
rect 95878 93548 95884 93560
rect 94740 93520 95884 93548
rect 94740 93508 94746 93520
rect 95878 93508 95884 93520
rect 95936 93508 95942 93560
rect 95050 93100 95056 93152
rect 95108 93140 95114 93152
rect 103514 93140 103520 93152
rect 95108 93112 103520 93140
rect 95108 93100 95114 93112
rect 103514 93100 103520 93112
rect 103572 93100 103578 93152
rect 67634 92828 67640 92880
rect 67692 92868 67698 92880
rect 68646 92868 68652 92880
rect 67692 92840 68652 92868
rect 67692 92828 67698 92840
rect 68646 92828 68652 92840
rect 68704 92828 68710 92880
rect 54846 92760 54852 92812
rect 54904 92800 54910 92812
rect 54904 92772 64874 92800
rect 54904 92760 54910 92772
rect 64846 92732 64874 92772
rect 72832 92732 72838 92744
rect 64846 92704 72838 92732
rect 72832 92692 72838 92704
rect 72890 92692 72896 92744
rect 91784 92692 91790 92744
rect 91842 92732 91848 92744
rect 94774 92732 94780 92744
rect 91842 92704 94780 92732
rect 91842 92692 91848 92704
rect 94774 92692 94780 92704
rect 94832 92692 94838 92744
rect 68462 92624 68468 92676
rect 68520 92664 68526 92676
rect 71728 92664 71734 92676
rect 68520 92636 71734 92664
rect 68520 92624 68526 92636
rect 71728 92624 71734 92636
rect 71786 92624 71792 92676
rect 52362 92420 52368 92472
rect 52420 92460 52426 92472
rect 86034 92460 86040 92472
rect 52420 92432 86040 92460
rect 52420 92420 52426 92432
rect 86034 92420 86040 92432
rect 86092 92420 86098 92472
rect 89254 92420 89260 92472
rect 89312 92460 89318 92472
rect 106274 92460 106280 92472
rect 89312 92432 106280 92460
rect 89312 92420 89318 92432
rect 106274 92420 106280 92432
rect 106332 92420 106338 92472
rect 63310 92352 63316 92404
rect 63368 92392 63374 92404
rect 73338 92392 73344 92404
rect 63368 92364 73344 92392
rect 63368 92352 63374 92364
rect 73338 92352 73344 92364
rect 73396 92352 73402 92404
rect 86678 92352 86684 92404
rect 86736 92392 86742 92404
rect 98730 92392 98736 92404
rect 86736 92364 98736 92392
rect 86736 92352 86742 92364
rect 98730 92352 98736 92364
rect 98788 92352 98794 92404
rect 90174 90992 90180 91044
rect 90232 91032 90238 91044
rect 95234 91032 95240 91044
rect 90232 91004 95240 91032
rect 90232 90992 90238 91004
rect 95234 90992 95240 91004
rect 95292 91032 95298 91044
rect 96154 91032 96160 91044
rect 95292 91004 96160 91032
rect 95292 90992 95298 91004
rect 96154 90992 96160 91004
rect 96212 90992 96218 91044
rect 88242 90856 88248 90908
rect 88300 90896 88306 90908
rect 117958 90896 117964 90908
rect 88300 90868 117964 90896
rect 88300 90856 88306 90868
rect 117958 90856 117964 90868
rect 118016 90856 118022 90908
rect 74350 90720 74356 90772
rect 74408 90760 74414 90772
rect 75270 90760 75276 90772
rect 74408 90732 75276 90760
rect 74408 90720 74414 90732
rect 75270 90720 75276 90732
rect 75328 90720 75334 90772
rect 87598 90516 87604 90568
rect 87656 90556 87662 90568
rect 88242 90556 88248 90568
rect 87656 90528 88248 90556
rect 87656 90516 87662 90528
rect 88242 90516 88248 90528
rect 88300 90516 88306 90568
rect 82630 89904 82636 89956
rect 82688 89944 82694 89956
rect 86862 89944 86868 89956
rect 82688 89916 86868 89944
rect 82688 89904 82694 89916
rect 86862 89904 86868 89916
rect 86920 89904 86926 89956
rect 80974 89700 80980 89752
rect 81032 89740 81038 89752
rect 83458 89740 83464 89752
rect 81032 89712 83464 89740
rect 81032 89700 81038 89712
rect 83458 89700 83464 89712
rect 83516 89700 83522 89752
rect 85206 89700 85212 89752
rect 85264 89740 85270 89752
rect 89530 89740 89536 89752
rect 85264 89712 89536 89740
rect 85264 89700 85270 89712
rect 89530 89700 89536 89712
rect 89588 89700 89594 89752
rect 48038 89632 48044 89684
rect 48096 89672 48102 89684
rect 78306 89672 78312 89684
rect 48096 89644 78312 89672
rect 48096 89632 48102 89644
rect 78306 89632 78312 89644
rect 78364 89632 78370 89684
rect 92382 89632 92388 89684
rect 92440 89672 92446 89684
rect 118694 89672 118700 89684
rect 92440 89644 118700 89672
rect 92440 89632 92446 89644
rect 118694 89632 118700 89644
rect 118752 89632 118758 89684
rect 52270 89564 52276 89616
rect 52328 89604 52334 89616
rect 76282 89604 76288 89616
rect 52328 89576 76288 89604
rect 52328 89564 52334 89576
rect 76282 89564 76288 89576
rect 76340 89564 76346 89616
rect 84102 89564 84108 89616
rect 84160 89604 84166 89616
rect 100018 89604 100024 89616
rect 84160 89576 100024 89604
rect 84160 89564 84166 89576
rect 100018 89564 100024 89576
rect 100076 89564 100082 89616
rect 119982 88952 119988 89004
rect 120040 88992 120046 89004
rect 137278 88992 137284 89004
rect 120040 88964 137284 88992
rect 120040 88952 120046 88964
rect 137278 88952 137284 88964
rect 137336 88952 137342 89004
rect 59170 88272 59176 88324
rect 59228 88312 59234 88324
rect 76558 88312 76564 88324
rect 59228 88284 76564 88312
rect 59228 88272 59234 88284
rect 76558 88272 76564 88284
rect 76616 88312 76622 88324
rect 76834 88312 76840 88324
rect 76616 88284 76840 88312
rect 76616 88272 76622 88284
rect 76834 88272 76840 88284
rect 76892 88272 76898 88324
rect 80054 88272 80060 88324
rect 80112 88312 80118 88324
rect 111794 88312 111800 88324
rect 80112 88284 111800 88312
rect 80112 88272 80118 88284
rect 111794 88272 111800 88284
rect 111852 88272 111858 88324
rect 60366 88204 60372 88256
rect 60424 88244 60430 88256
rect 73798 88244 73804 88256
rect 60424 88216 73804 88244
rect 60424 88204 60430 88216
rect 73798 88204 73804 88216
rect 73856 88204 73862 88256
rect 87230 88204 87236 88256
rect 87288 88244 87294 88256
rect 115934 88244 115940 88256
rect 87288 88216 115940 88244
rect 87288 88204 87294 88216
rect 115934 88204 115940 88216
rect 115992 88204 115998 88256
rect 111794 87592 111800 87644
rect 111852 87632 111858 87644
rect 188430 87632 188436 87644
rect 111852 87604 188436 87632
rect 111852 87592 111858 87604
rect 188430 87592 188436 87604
rect 188488 87592 188494 87644
rect 65610 86912 65616 86964
rect 65668 86952 65674 86964
rect 96706 86952 96712 86964
rect 65668 86924 96712 86952
rect 65668 86912 65674 86924
rect 96706 86912 96712 86924
rect 96764 86912 96770 86964
rect 61746 86844 61752 86896
rect 61804 86884 61810 86896
rect 75178 86884 75184 86896
rect 61804 86856 75184 86884
rect 61804 86844 61810 86856
rect 75178 86844 75184 86856
rect 75236 86884 75242 86896
rect 75362 86884 75368 86896
rect 75236 86856 75368 86884
rect 75236 86844 75242 86856
rect 75362 86844 75368 86856
rect 75420 86844 75426 86896
rect 88150 86844 88156 86896
rect 88208 86884 88214 86896
rect 101490 86884 101496 86896
rect 88208 86856 101496 86884
rect 88208 86844 88214 86856
rect 101490 86844 101496 86856
rect 101548 86844 101554 86896
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 56594 85524 56600 85536
rect 3568 85496 56600 85524
rect 3568 85484 3574 85496
rect 56594 85484 56600 85496
rect 56652 85484 56658 85536
rect 86862 85484 86868 85536
rect 86920 85524 86926 85536
rect 97994 85524 98000 85536
rect 86920 85496 98000 85524
rect 86920 85484 86926 85496
rect 97994 85484 98000 85496
rect 98052 85484 98058 85536
rect 66070 84804 66076 84856
rect 66128 84844 66134 84856
rect 338206 84844 338212 84856
rect 66128 84816 338212 84844
rect 66128 84804 66134 84816
rect 338206 84804 338212 84816
rect 338264 84804 338270 84856
rect 56318 84124 56324 84176
rect 56376 84164 56382 84176
rect 78674 84164 78680 84176
rect 56376 84136 78680 84164
rect 56376 84124 56382 84136
rect 78674 84124 78680 84136
rect 78732 84124 78738 84176
rect 92474 84124 92480 84176
rect 92532 84164 92538 84176
rect 93762 84164 93768 84176
rect 92532 84136 93768 84164
rect 92532 84124 92538 84136
rect 93762 84124 93768 84136
rect 93820 84164 93826 84176
rect 128538 84164 128544 84176
rect 93820 84136 128544 84164
rect 93820 84124 93826 84136
rect 128538 84124 128544 84136
rect 128596 84124 128602 84176
rect 85574 84056 85580 84108
rect 85632 84096 85638 84108
rect 86770 84096 86776 84108
rect 85632 84068 86776 84096
rect 85632 84056 85638 84068
rect 86770 84056 86776 84068
rect 86828 84096 86834 84108
rect 99374 84096 99380 84108
rect 86828 84068 99380 84096
rect 86828 84056 86834 84068
rect 99374 84056 99380 84068
rect 99432 84056 99438 84108
rect 78674 82832 78680 82884
rect 78732 82872 78738 82884
rect 79318 82872 79324 82884
rect 78732 82844 79324 82872
rect 78732 82832 78738 82844
rect 79318 82832 79324 82844
rect 79376 82832 79382 82884
rect 83458 82764 83464 82816
rect 83516 82804 83522 82816
rect 84102 82804 84108 82816
rect 83516 82776 84108 82804
rect 83516 82764 83522 82776
rect 84102 82764 84108 82776
rect 84160 82804 84166 82816
rect 107654 82804 107660 82816
rect 84160 82776 107660 82804
rect 84160 82764 84166 82776
rect 107654 82764 107660 82776
rect 107712 82764 107718 82816
rect 63218 82084 63224 82136
rect 63276 82124 63282 82136
rect 327166 82124 327172 82136
rect 63276 82096 327172 82124
rect 63276 82084 63282 82096
rect 327166 82084 327172 82096
rect 327224 82084 327230 82136
rect 62022 80724 62028 80776
rect 62080 80764 62086 80776
rect 151078 80764 151084 80776
rect 62080 80736 151084 80764
rect 62080 80724 62086 80736
rect 151078 80724 151084 80736
rect 151136 80724 151142 80776
rect 96154 80656 96160 80708
rect 96212 80696 96218 80708
rect 349154 80696 349160 80708
rect 96212 80668 349160 80696
rect 96212 80656 96218 80668
rect 349154 80656 349160 80668
rect 349212 80656 349218 80708
rect 67174 79296 67180 79348
rect 67232 79336 67238 79348
rect 280154 79336 280160 79348
rect 67232 79308 280160 79336
rect 67232 79296 67238 79308
rect 280154 79296 280160 79308
rect 280212 79296 280218 79348
rect 75270 78616 75276 78668
rect 75328 78656 75334 78668
rect 100754 78656 100760 78668
rect 75328 78628 100760 78656
rect 75328 78616 75334 78628
rect 100754 78616 100760 78628
rect 100812 78656 100818 78668
rect 101122 78656 101128 78668
rect 100812 78628 101128 78656
rect 100812 78616 100818 78628
rect 101122 78616 101128 78628
rect 101180 78616 101186 78668
rect 48130 78004 48136 78056
rect 48188 78044 48194 78056
rect 123570 78044 123576 78056
rect 48188 78016 123576 78044
rect 48188 78004 48194 78016
rect 123570 78004 123576 78016
rect 123628 78004 123634 78056
rect 101122 77936 101128 77988
rect 101180 77976 101186 77988
rect 340874 77976 340880 77988
rect 101180 77948 340880 77976
rect 101180 77936 101186 77948
rect 340874 77936 340880 77948
rect 340932 77936 340938 77988
rect 63402 77188 63408 77240
rect 63460 77228 63466 77240
rect 252554 77228 252560 77240
rect 63460 77200 252560 77228
rect 63460 77188 63466 77200
rect 252554 77188 252560 77200
rect 252612 77228 252618 77240
rect 253198 77228 253204 77240
rect 252612 77200 253204 77228
rect 252612 77188 252618 77200
rect 253198 77188 253204 77200
rect 253256 77188 253262 77240
rect 79962 75148 79968 75200
rect 80020 75188 80026 75200
rect 184198 75188 184204 75200
rect 80020 75160 184204 75188
rect 80020 75148 80026 75160
rect 184198 75148 184204 75160
rect 184256 75148 184262 75200
rect 108942 73788 108948 73840
rect 109000 73828 109006 73840
rect 146938 73828 146944 73840
rect 109000 73800 146944 73828
rect 109000 73788 109006 73800
rect 146938 73788 146944 73800
rect 146996 73788 147002 73840
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 101398 71720 101404 71732
rect 3568 71692 101404 71720
rect 3568 71680 3574 71692
rect 101398 71680 101404 71692
rect 101456 71680 101462 71732
rect 96522 71000 96528 71052
rect 96580 71040 96586 71052
rect 155310 71040 155316 71052
rect 96580 71012 155316 71040
rect 96580 71000 96586 71012
rect 155310 71000 155316 71012
rect 155368 71000 155374 71052
rect 79318 69640 79324 69692
rect 79376 69680 79382 69692
rect 343634 69680 343640 69692
rect 79376 69652 343640 69680
rect 79376 69640 79382 69652
rect 343634 69640 343640 69652
rect 343692 69640 343698 69692
rect 66070 68348 66076 68400
rect 66128 68388 66134 68400
rect 162118 68388 162124 68400
rect 66128 68360 162124 68388
rect 66128 68348 66134 68360
rect 162118 68348 162124 68360
rect 162176 68348 162182 68400
rect 70302 68280 70308 68332
rect 70360 68320 70366 68332
rect 180058 68320 180064 68332
rect 70360 68292 180064 68320
rect 70360 68280 70366 68292
rect 180058 68280 180064 68292
rect 180116 68280 180122 68332
rect 65518 66852 65524 66904
rect 65576 66892 65582 66904
rect 332594 66892 332600 66904
rect 65576 66864 332600 66892
rect 65576 66852 65582 66864
rect 332594 66852 332600 66864
rect 332652 66852 332658 66904
rect 10962 65492 10968 65544
rect 11020 65532 11026 65544
rect 178678 65532 178684 65544
rect 11020 65504 178684 65532
rect 11020 65492 11026 65504
rect 178678 65492 178684 65504
rect 178736 65492 178742 65544
rect 68922 64132 68928 64184
rect 68980 64172 68986 64184
rect 189718 64172 189724 64184
rect 68980 64144 189724 64172
rect 68980 64132 68986 64144
rect 189718 64132 189724 64144
rect 189776 64132 189782 64184
rect 70210 62772 70216 62824
rect 70268 62812 70274 62824
rect 311894 62812 311900 62824
rect 70268 62784 311900 62812
rect 70268 62772 70274 62784
rect 311894 62772 311900 62784
rect 311952 62772 311958 62824
rect 95050 61412 95056 61464
rect 95108 61452 95114 61464
rect 141510 61452 141516 61464
rect 95108 61424 141516 61452
rect 95108 61412 95114 61424
rect 141510 61412 141516 61424
rect 141568 61412 141574 61464
rect 72418 61344 72424 61396
rect 72476 61384 72482 61396
rect 97258 61384 97264 61396
rect 72476 61356 97264 61384
rect 72476 61344 72482 61356
rect 97258 61344 97264 61356
rect 97316 61344 97322 61396
rect 128998 61344 129004 61396
rect 129056 61384 129062 61396
rect 206370 61384 206376 61396
rect 129056 61356 206376 61384
rect 129056 61344 129062 61356
rect 206370 61344 206376 61356
rect 206428 61344 206434 61396
rect 304258 60664 304264 60716
rect 304316 60704 304322 60716
rect 580166 60704 580172 60716
rect 304316 60676 580172 60704
rect 304316 60664 304322 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 67634 59984 67640 60036
rect 67692 60024 67698 60036
rect 291194 60024 291200 60036
rect 67692 59996 291200 60024
rect 67692 59984 67698 59996
rect 291194 59984 291200 59996
rect 291252 59984 291258 60036
rect 86770 58624 86776 58676
rect 86828 58664 86834 58676
rect 253198 58664 253204 58676
rect 86828 58636 253204 58664
rect 86828 58624 86834 58636
rect 253198 58624 253204 58636
rect 253256 58624 253262 58676
rect 71682 57264 71688 57316
rect 71740 57304 71746 57316
rect 173158 57304 173164 57316
rect 71740 57276 173164 57304
rect 71740 57264 71746 57276
rect 173158 57264 173164 57276
rect 173216 57264 173222 57316
rect 165522 57196 165528 57248
rect 165580 57236 165586 57248
rect 304258 57236 304264 57248
rect 165580 57208 304264 57236
rect 165580 57196 165586 57208
rect 304258 57196 304264 57208
rect 304316 57196 304322 57248
rect 67542 56516 67548 56568
rect 67600 56556 67606 56568
rect 269114 56556 269120 56568
rect 67600 56528 269120 56556
rect 67600 56516 67606 56528
rect 269114 56516 269120 56528
rect 269172 56516 269178 56568
rect 88150 54476 88156 54528
rect 88208 54516 88214 54528
rect 266354 54516 266360 54528
rect 88208 54488 266360 54516
rect 88208 54476 88214 54488
rect 266354 54476 266360 54488
rect 266412 54476 266418 54528
rect 75178 53048 75184 53100
rect 75236 53088 75242 53100
rect 224218 53088 224224 53100
rect 75236 53060 224224 53088
rect 75236 53048 75242 53060
rect 224218 53048 224224 53060
rect 224276 53048 224282 53100
rect 75822 51688 75828 51740
rect 75880 51728 75886 51740
rect 177298 51728 177304 51740
rect 75880 51700 177304 51728
rect 75880 51688 75886 51700
rect 177298 51688 177304 51700
rect 177356 51688 177362 51740
rect 193122 51688 193128 51740
rect 193180 51728 193186 51740
rect 242986 51728 242992 51740
rect 193180 51700 242992 51728
rect 193180 51688 193186 51700
rect 242986 51688 242992 51700
rect 243044 51688 243050 51740
rect 59262 50396 59268 50448
rect 59320 50436 59326 50448
rect 166258 50436 166264 50448
rect 59320 50408 166264 50436
rect 59320 50396 59326 50408
rect 166258 50396 166264 50408
rect 166316 50396 166322 50448
rect 89530 50328 89536 50380
rect 89588 50368 89594 50380
rect 289078 50368 289084 50380
rect 89588 50340 289084 50368
rect 89588 50328 89594 50340
rect 289078 50328 289084 50340
rect 289136 50328 289142 50380
rect 73798 48968 73804 49020
rect 73856 49008 73862 49020
rect 231118 49008 231124 49020
rect 73856 48980 231124 49008
rect 73856 48968 73862 48980
rect 231118 48968 231124 48980
rect 231176 48968 231182 49020
rect 248414 48492 248420 48544
rect 248472 48532 248478 48544
rect 252554 48532 252560 48544
rect 248472 48504 252560 48532
rect 248472 48492 248478 48504
rect 252554 48492 252560 48504
rect 252612 48492 252618 48544
rect 76558 46180 76564 46232
rect 76616 46220 76622 46232
rect 322198 46220 322204 46232
rect 76616 46192 322204 46220
rect 76616 46180 76622 46192
rect 322198 46180 322204 46192
rect 322256 46180 322262 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 60734 45540 60740 45552
rect 3476 45512 60740 45540
rect 3476 45500 3482 45512
rect 60734 45500 60740 45512
rect 60792 45500 60798 45552
rect 93762 44820 93768 44872
rect 93820 44860 93826 44872
rect 302326 44860 302332 44872
rect 93820 44832 302332 44860
rect 93820 44820 93826 44832
rect 302326 44820 302332 44832
rect 302384 44820 302390 44872
rect 84102 43392 84108 43444
rect 84160 43432 84166 43444
rect 274634 43432 274640 43444
rect 84160 43404 274640 43432
rect 84160 43392 84166 43404
rect 274634 43392 274640 43404
rect 274692 43392 274698 43444
rect 249058 42304 249064 42356
rect 249116 42344 249122 42356
rect 249794 42344 249800 42356
rect 249116 42316 249800 42344
rect 249116 42304 249122 42316
rect 249794 42304 249800 42316
rect 249852 42304 249858 42356
rect 88242 42032 88248 42084
rect 88300 42072 88306 42084
rect 284386 42072 284392 42084
rect 88300 42044 284392 42072
rect 88300 42032 88306 42044
rect 284386 42032 284392 42044
rect 284444 42032 284450 42084
rect 64598 40672 64604 40724
rect 64656 40712 64662 40724
rect 307846 40712 307852 40724
rect 64656 40684 307852 40712
rect 64656 40672 64662 40684
rect 307846 40672 307852 40684
rect 307904 40672 307910 40724
rect 197998 39312 198004 39364
rect 198056 39352 198062 39364
rect 262858 39352 262864 39364
rect 198056 39324 262864 39352
rect 198056 39312 198062 39324
rect 262858 39312 262864 39324
rect 262916 39312 262922 39364
rect 3970 37884 3976 37936
rect 4028 37924 4034 37936
rect 160830 37924 160836 37936
rect 4028 37896 160836 37924
rect 4028 37884 4034 37896
rect 160830 37884 160836 37896
rect 160888 37884 160894 37936
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 14458 33096 14464 33108
rect 3568 33068 14464 33096
rect 3568 33056 3574 33068
rect 14458 33056 14464 33068
rect 14516 33056 14522 33108
rect 82722 32376 82728 32428
rect 82780 32416 82786 32428
rect 147030 32416 147036 32428
rect 82780 32388 147036 32416
rect 82780 32376 82786 32388
rect 147030 32376 147036 32388
rect 147088 32376 147094 32428
rect 88978 26868 88984 26920
rect 89036 26908 89042 26920
rect 213178 26908 213184 26920
rect 89036 26880 213184 26908
rect 89036 26868 89042 26880
rect 213178 26868 213184 26880
rect 213236 26868 213242 26920
rect 280798 22720 280804 22772
rect 280856 22760 280862 22772
rect 292666 22760 292672 22772
rect 280856 22732 292672 22760
rect 280856 22720 280862 22732
rect 292666 22720 292672 22732
rect 292724 22720 292730 22772
rect 295978 22720 295984 22772
rect 296036 22760 296042 22772
rect 335354 22760 335360 22772
rect 296036 22732 335360 22760
rect 296036 22720 296042 22732
rect 335354 22720 335360 22732
rect 335412 22720 335418 22772
rect 151170 21360 151176 21412
rect 151228 21400 151234 21412
rect 277486 21400 277492 21412
rect 151228 21372 277492 21400
rect 151228 21360 151234 21372
rect 277486 21360 277492 21372
rect 277544 21360 277550 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 72418 20652 72424 20664
rect 3476 20624 72424 20652
rect 3476 20612 3482 20624
rect 72418 20612 72424 20624
rect 72476 20612 72482 20664
rect 78582 20000 78588 20052
rect 78640 20040 78646 20052
rect 175918 20040 175924 20052
rect 78640 20012 175924 20040
rect 78640 20000 78646 20012
rect 175918 20000 175924 20012
rect 175976 20000 175982 20052
rect 170490 19932 170496 19984
rect 170548 19972 170554 19984
rect 325694 19972 325700 19984
rect 170548 19944 325700 19972
rect 170548 19932 170554 19944
rect 325694 19932 325700 19944
rect 325752 19932 325758 19984
rect 88242 18640 88248 18692
rect 88300 18680 88306 18692
rect 206278 18680 206284 18692
rect 88300 18652 206284 18680
rect 88300 18640 88306 18652
rect 206278 18640 206284 18652
rect 206336 18640 206342 18692
rect 50982 18572 50988 18624
rect 51040 18612 51046 18624
rect 186958 18612 186964 18624
rect 51040 18584 186964 18612
rect 51040 18572 51046 18584
rect 186958 18572 186964 18584
rect 187016 18572 187022 18624
rect 220078 18572 220084 18624
rect 220136 18612 220142 18624
rect 331306 18612 331312 18624
rect 220136 18584 331312 18612
rect 220136 18572 220142 18584
rect 331306 18572 331312 18584
rect 331364 18572 331370 18624
rect 97902 17280 97908 17332
rect 97960 17320 97966 17332
rect 142798 17320 142804 17332
rect 97960 17292 142804 17320
rect 97960 17280 97966 17292
rect 142798 17280 142804 17292
rect 142856 17280 142862 17332
rect 65978 17212 65984 17264
rect 66036 17252 66042 17264
rect 125594 17252 125600 17264
rect 66036 17224 125600 17252
rect 66036 17212 66042 17224
rect 125594 17212 125600 17224
rect 125652 17212 125658 17264
rect 253198 17212 253204 17264
rect 253256 17252 253262 17264
rect 287146 17252 287152 17264
rect 253256 17224 287152 17252
rect 253256 17212 253262 17224
rect 287146 17212 287152 17224
rect 287204 17212 287210 17264
rect 307846 16192 307852 16244
rect 307904 16232 307910 16244
rect 309042 16232 309048 16244
rect 307904 16204 309048 16232
rect 307904 16192 307910 16204
rect 309042 16192 309048 16204
rect 309100 16192 309106 16244
rect 64782 15920 64788 15972
rect 64840 15960 64846 15972
rect 148318 15960 148324 15972
rect 64840 15932 148324 15960
rect 64840 15920 64846 15932
rect 148318 15920 148324 15932
rect 148376 15920 148382 15972
rect 86862 15852 86868 15904
rect 86920 15892 86926 15904
rect 322934 15892 322940 15904
rect 86920 15864 322940 15892
rect 86920 15852 86926 15864
rect 322934 15852 322940 15864
rect 322992 15852 322998 15904
rect 46658 14424 46664 14476
rect 46716 14464 46722 14476
rect 170398 14464 170404 14476
rect 46716 14436 170404 14464
rect 46716 14424 46722 14436
rect 170398 14424 170404 14436
rect 170456 14424 170462 14476
rect 173250 14424 173256 14476
rect 173308 14464 173314 14476
rect 337010 14464 337016 14476
rect 173308 14436 337016 14464
rect 173308 14424 173314 14436
rect 337010 14424 337016 14436
rect 337068 14424 337074 14476
rect 89530 13132 89536 13184
rect 89588 13172 89594 13184
rect 185578 13172 185584 13184
rect 89588 13144 185584 13172
rect 89588 13132 89594 13144
rect 185578 13132 185584 13144
rect 185636 13132 185642 13184
rect 45370 13064 45376 13116
rect 45428 13104 45434 13116
rect 160738 13104 160744 13116
rect 45428 13076 160744 13104
rect 45428 13064 45434 13076
rect 160738 13064 160744 13076
rect 160796 13064 160802 13116
rect 273898 13064 273904 13116
rect 273956 13104 273962 13116
rect 324866 13104 324872 13116
rect 273956 13076 324872 13104
rect 273956 13064 273962 13076
rect 324866 13064 324872 13076
rect 324924 13064 324930 13116
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 7558 12424 7564 12436
rect 3476 12396 7564 12424
rect 3476 12384 3482 12396
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 178770 11704 178776 11756
rect 178828 11744 178834 11756
rect 241698 11744 241704 11756
rect 178828 11716 241704 11744
rect 178828 11704 178834 11716
rect 241698 11704 241704 11716
rect 241756 11704 241762 11756
rect 262858 11704 262864 11756
rect 262916 11744 262922 11756
rect 302878 11744 302884 11756
rect 262916 11716 302884 11744
rect 262916 11704 262922 11716
rect 302878 11704 302884 11716
rect 302936 11704 302942 11756
rect 89622 10956 89628 11008
rect 89680 10996 89686 11008
rect 333974 10996 333980 11008
rect 89680 10968 333980 10996
rect 89680 10956 89686 10968
rect 333974 10956 333980 10968
rect 334032 10996 334038 11008
rect 334618 10996 334624 11008
rect 334032 10968 334624 10996
rect 334032 10956 334038 10968
rect 334618 10956 334624 10968
rect 334676 10956 334682 11008
rect 106 10276 112 10328
rect 164 10316 170 10328
rect 96614 10316 96620 10328
rect 164 10288 96620 10316
rect 164 10276 170 10288
rect 96614 10276 96620 10288
rect 96672 10276 96678 10328
rect 61930 8916 61936 8968
rect 61988 8956 61994 8968
rect 169018 8956 169024 8968
rect 61988 8928 169024 8956
rect 61988 8916 61994 8928
rect 169018 8916 169024 8928
rect 169076 8916 169082 8968
rect 180150 8916 180156 8968
rect 180208 8956 180214 8968
rect 346946 8956 346952 8968
rect 180208 8928 346952 8956
rect 180208 8916 180214 8928
rect 346946 8916 346952 8928
rect 347004 8916 347010 8968
rect 54938 7556 54944 7608
rect 54996 7596 55002 7608
rect 128998 7596 129004 7608
rect 54996 7568 129004 7596
rect 54996 7556 55002 7568
rect 128998 7556 129004 7568
rect 129056 7556 129062 7608
rect 184290 7556 184296 7608
rect 184348 7596 184354 7608
rect 317322 7596 317328 7608
rect 184348 7568 317328 7596
rect 184348 7556 184354 7568
rect 317322 7556 317328 7568
rect 317380 7556 317386 7608
rect 92474 6196 92480 6248
rect 92532 6236 92538 6248
rect 155218 6236 155224 6248
rect 92532 6208 155224 6236
rect 92532 6196 92538 6208
rect 155218 6196 155224 6208
rect 155276 6196 155282 6248
rect 83274 6128 83280 6180
rect 83332 6168 83338 6180
rect 159358 6168 159364 6180
rect 83332 6140 159364 6168
rect 83332 6128 83338 6140
rect 159358 6128 159364 6140
rect 159416 6128 159422 6180
rect 198090 6128 198096 6180
rect 198148 6168 198154 6180
rect 247586 6168 247592 6180
rect 198148 6140 247592 6168
rect 198148 6128 198154 6140
rect 247586 6128 247592 6140
rect 247644 6128 247650 6180
rect 261754 6128 261760 6180
rect 261812 6168 261818 6180
rect 270494 6168 270500 6180
rect 261812 6140 270500 6168
rect 261812 6128 261818 6140
rect 270494 6128 270500 6140
rect 270552 6128 270558 6180
rect 305638 6128 305644 6180
rect 305696 6168 305702 6180
rect 311434 6168 311440 6180
rect 305696 6140 311440 6168
rect 305696 6128 305702 6140
rect 311434 6128 311440 6140
rect 311492 6128 311498 6180
rect 310238 5516 310244 5568
rect 310296 5556 310302 5568
rect 313274 5556 313280 5568
rect 310296 5528 313280 5556
rect 310296 5516 310302 5528
rect 313274 5516 313280 5528
rect 313332 5516 313338 5568
rect 187050 4768 187056 4820
rect 187108 4808 187114 4820
rect 257062 4808 257068 4820
rect 187108 4780 257068 4808
rect 187108 4768 187114 4780
rect 257062 4768 257068 4780
rect 257120 4768 257126 4820
rect 264238 4768 264244 4820
rect 264296 4808 264302 4820
rect 279510 4808 279516 4820
rect 264296 4780 279516 4808
rect 264296 4768 264302 4780
rect 279510 4768 279516 4780
rect 279568 4768 279574 4820
rect 281902 4768 281908 4820
rect 281960 4808 281966 4820
rect 287054 4808 287060 4820
rect 281960 4780 287060 4808
rect 281960 4768 281966 4780
rect 287054 4768 287060 4780
rect 287112 4768 287118 4820
rect 122282 4088 122288 4140
rect 122340 4128 122346 4140
rect 123478 4128 123484 4140
rect 122340 4100 123484 4128
rect 122340 4088 122346 4100
rect 123478 4088 123484 4100
rect 123536 4088 123542 4140
rect 304258 3952 304264 4004
rect 304316 3992 304322 4004
rect 307938 3992 307944 4004
rect 304316 3964 307944 3992
rect 304316 3952 304322 3964
rect 307938 3952 307944 3964
rect 307996 3952 308002 4004
rect 342162 3680 342168 3732
rect 342220 3720 342226 3732
rect 345014 3720 345020 3732
rect 342220 3692 345020 3720
rect 342220 3680 342226 3692
rect 345014 3680 345020 3692
rect 345072 3680 345078 3732
rect 30098 3612 30104 3664
rect 30156 3652 30162 3664
rect 40678 3652 40684 3664
rect 30156 3624 40684 3652
rect 30156 3612 30162 3624
rect 40678 3612 40684 3624
rect 40736 3612 40742 3664
rect 108298 3652 108304 3664
rect 103486 3624 108304 3652
rect 13538 3584 13544 3596
rect 6886 3556 13544 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 6886 3516 6914 3556
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 53650 3584 53656 3596
rect 52604 3556 53656 3584
rect 52604 3544 52610 3556
rect 53650 3544 53656 3556
rect 53708 3544 53714 3596
rect 60826 3544 60832 3596
rect 60884 3584 60890 3596
rect 62022 3584 62028 3596
rect 60884 3556 62028 3584
rect 60884 3544 60890 3556
rect 62022 3544 62028 3556
rect 62080 3544 62086 3596
rect 72510 3584 72516 3596
rect 64846 3556 72516 3584
rect 5500 3488 6914 3516
rect 5500 3476 5506 3488
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12342 3516 12348 3528
rect 11204 3488 12348 3516
rect 11204 3476 11210 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16390 3516 16396 3528
rect 15988 3488 16396 3516
rect 15988 3476 15994 3488
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20530 3516 20536 3528
rect 19484 3488 20536 3516
rect 19484 3476 19490 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 21358 3516 21364 3528
rect 20680 3488 21364 3516
rect 20680 3476 20686 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 35986 3476 35992 3528
rect 36044 3516 36050 3528
rect 37090 3516 37096 3528
rect 36044 3488 37096 3516
rect 36044 3476 36050 3488
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41322 3516 41328 3528
rect 40736 3488 41328 3516
rect 40736 3476 40742 3488
rect 41322 3476 41328 3488
rect 41380 3476 41386 3528
rect 41874 3476 41880 3528
rect 41932 3516 41938 3528
rect 42702 3516 42708 3528
rect 41932 3488 42708 3516
rect 41932 3476 41938 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 43990 3516 43996 3528
rect 43128 3488 43996 3516
rect 43128 3476 43134 3488
rect 43990 3476 43996 3488
rect 44048 3476 44054 3528
rect 44266 3476 44272 3528
rect 44324 3516 44330 3528
rect 45370 3516 45376 3528
rect 44324 3488 45376 3516
rect 44324 3476 44330 3488
rect 45370 3476 45376 3488
rect 45428 3476 45434 3528
rect 48222 3476 48228 3528
rect 48280 3516 48286 3528
rect 48958 3516 48964 3528
rect 48280 3488 48964 3516
rect 48280 3476 48286 3488
rect 48958 3476 48964 3488
rect 49016 3476 49022 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50982 3516 50988 3528
rect 50212 3488 50988 3516
rect 50212 3476 50218 3488
rect 50982 3476 50988 3488
rect 51040 3476 51046 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 64846 3516 64874 3556
rect 72510 3544 72516 3556
rect 72568 3544 72574 3596
rect 92750 3544 92756 3596
rect 92808 3584 92814 3596
rect 103486 3584 103514 3624
rect 108298 3612 108304 3624
rect 108356 3612 108362 3664
rect 119338 3584 119344 3596
rect 92808 3556 103514 3584
rect 106844 3556 119344 3584
rect 92808 3544 92814 3556
rect 59688 3488 64874 3516
rect 59688 3476 59694 3488
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 70210 3516 70216 3528
rect 69164 3488 70216 3516
rect 69164 3476 69170 3488
rect 70210 3476 70216 3488
rect 70268 3476 70274 3528
rect 73798 3476 73804 3528
rect 73856 3516 73862 3528
rect 74442 3516 74448 3528
rect 73856 3488 74448 3516
rect 73856 3476 73862 3488
rect 74442 3476 74448 3488
rect 74500 3476 74506 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 82722 3516 82728 3528
rect 82136 3488 82728 3516
rect 82136 3476 82142 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 86862 3476 86868 3528
rect 86920 3516 86926 3528
rect 87598 3516 87604 3528
rect 86920 3488 87604 3516
rect 86920 3476 86926 3488
rect 87598 3476 87604 3488
rect 87656 3476 87662 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 92382 3516 92388 3528
rect 91612 3488 92388 3516
rect 91612 3476 91618 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 97902 3516 97908 3528
rect 97500 3488 97908 3516
rect 97500 3476 97506 3488
rect 97902 3476 97908 3488
rect 97960 3476 97966 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 106844 3516 106872 3556
rect 119338 3544 119344 3556
rect 119396 3544 119402 3596
rect 123478 3544 123484 3596
rect 123536 3584 123542 3596
rect 123536 3556 132494 3584
rect 123536 3544 123542 3556
rect 99892 3488 106872 3516
rect 99892 3476 99898 3488
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 121086 3476 121092 3528
rect 121144 3516 121150 3528
rect 122098 3516 122104 3528
rect 121144 3488 122104 3516
rect 121144 3476 121150 3488
rect 122098 3476 122104 3488
rect 122156 3476 122162 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 132466 3516 132494 3556
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277118 3584 277124 3596
rect 276072 3556 277124 3584
rect 276072 3544 276078 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 134518 3516 134524 3528
rect 132466 3488 134524 3516
rect 134518 3476 134524 3488
rect 134576 3476 134582 3528
rect 143534 3476 143540 3528
rect 143592 3516 143598 3528
rect 144822 3516 144828 3528
rect 143592 3488 144828 3516
rect 143592 3476 143598 3488
rect 144822 3476 144828 3488
rect 144880 3476 144886 3528
rect 224218 3476 224224 3528
rect 224276 3516 224282 3528
rect 246390 3516 246396 3528
rect 224276 3488 246396 3516
rect 224276 3476 224282 3488
rect 246390 3476 246396 3488
rect 246448 3476 246454 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 270586 3516 270592 3528
rect 264204 3488 270592 3516
rect 264204 3476 264210 3488
rect 270586 3476 270592 3488
rect 270644 3476 270650 3528
rect 282178 3476 282184 3528
rect 282236 3516 282242 3528
rect 283098 3516 283104 3528
rect 282236 3488 283104 3516
rect 282236 3476 282242 3488
rect 283098 3476 283104 3488
rect 283156 3476 283162 3528
rect 291838 3476 291844 3528
rect 291896 3516 291902 3528
rect 292574 3516 292580 3528
rect 291896 3488 292580 3516
rect 291896 3476 291902 3488
rect 292574 3476 292580 3488
rect 292632 3476 292638 3528
rect 297266 3476 297272 3528
rect 297324 3516 297330 3528
rect 299474 3516 299480 3528
rect 297324 3488 299480 3516
rect 297324 3476 297330 3488
rect 299474 3476 299480 3488
rect 299532 3476 299538 3528
rect 309778 3476 309784 3528
rect 309836 3516 309842 3528
rect 313826 3516 313832 3528
rect 309836 3488 313832 3516
rect 309836 3476 309842 3488
rect 313826 3476 313832 3488
rect 313884 3476 313890 3528
rect 322198 3476 322204 3528
rect 322256 3516 322262 3528
rect 324406 3516 324412 3528
rect 322256 3488 324412 3516
rect 322256 3476 322262 3488
rect 324406 3476 324412 3488
rect 324464 3476 324470 3528
rect 329190 3476 329196 3528
rect 329248 3516 329254 3528
rect 331214 3516 331220 3528
rect 329248 3488 331220 3516
rect 329248 3476 329254 3488
rect 331214 3476 331220 3488
rect 331272 3476 331278 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 582926 3516 582932 3528
rect 582248 3488 582932 3516
rect 582248 3476 582254 3488
rect 582926 3476 582932 3488
rect 582984 3476 582990 3528
rect 18598 3448 18604 3460
rect 12360 3420 18604 3448
rect 12360 3392 12388 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 50338 3448 50344 3460
rect 24268 3420 50344 3448
rect 24268 3408 24274 3420
rect 50338 3408 50344 3420
rect 50396 3408 50402 3460
rect 64322 3408 64328 3460
rect 64380 3448 64386 3460
rect 64782 3448 64788 3460
rect 64380 3420 64788 3448
rect 64380 3408 64386 3420
rect 64782 3408 64788 3420
rect 64840 3408 64846 3460
rect 72602 3408 72608 3460
rect 72660 3448 72666 3460
rect 92474 3448 92480 3460
rect 72660 3420 92480 3448
rect 72660 3408 72666 3420
rect 92474 3408 92480 3420
rect 92532 3408 92538 3460
rect 118786 3408 118792 3460
rect 118844 3448 118850 3460
rect 141418 3448 141424 3460
rect 118844 3420 141424 3448
rect 118844 3408 118850 3420
rect 141418 3408 141424 3420
rect 141476 3408 141482 3460
rect 188430 3408 188436 3460
rect 188488 3448 188494 3460
rect 242894 3448 242900 3460
rect 188488 3420 242900 3448
rect 188488 3408 188494 3420
rect 242894 3408 242900 3420
rect 242952 3408 242958 3460
rect 246298 3408 246304 3460
rect 246356 3448 246362 3460
rect 253474 3448 253480 3460
rect 246356 3420 253480 3448
rect 246356 3408 246362 3420
rect 253474 3408 253480 3420
rect 253532 3408 253538 3460
rect 256050 3408 256056 3460
rect 256108 3448 256114 3460
rect 265342 3448 265348 3460
rect 256108 3420 265348 3448
rect 256108 3408 256114 3420
rect 265342 3408 265348 3420
rect 265400 3408 265406 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 271230 3448 271236 3460
rect 267056 3420 271236 3448
rect 267056 3408 267062 3420
rect 271230 3408 271236 3420
rect 271288 3408 271294 3460
rect 315022 3408 315028 3460
rect 315080 3448 315086 3460
rect 327074 3448 327080 3460
rect 315080 3420 327080 3448
rect 315080 3408 315086 3420
rect 327074 3408 327080 3420
rect 327132 3408 327138 3460
rect 330386 3408 330392 3460
rect 330444 3448 330450 3460
rect 338114 3448 338120 3460
rect 330444 3420 338120 3448
rect 330444 3408 330450 3420
rect 338114 3408 338120 3420
rect 338172 3408 338178 3460
rect 351638 3408 351644 3460
rect 351696 3448 351702 3460
rect 357434 3448 357440 3460
rect 351696 3420 357440 3448
rect 351696 3408 351702 3420
rect 357434 3408 357440 3420
rect 357492 3408 357498 3460
rect 1302 3340 1308 3392
rect 1360 3380 1366 3392
rect 7650 3380 7656 3392
rect 1360 3352 7656 3380
rect 1360 3340 1366 3352
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 12342 3340 12348 3392
rect 12400 3340 12406 3392
rect 289078 3340 289084 3392
rect 289136 3380 289142 3392
rect 294874 3380 294880 3392
rect 289136 3352 294880 3380
rect 289136 3340 289142 3352
rect 294874 3340 294880 3352
rect 294932 3340 294938 3392
rect 345750 3340 345756 3392
rect 345808 3380 345814 3392
rect 351914 3380 351920 3392
rect 345808 3352 351920 3380
rect 345808 3340 345814 3352
rect 351914 3340 351920 3352
rect 351972 3340 351978 3392
rect 272426 3204 272432 3256
rect 272484 3244 272490 3256
rect 277394 3244 277400 3256
rect 272484 3216 277400 3244
rect 272484 3204 272490 3216
rect 277394 3204 277400 3216
rect 277452 3204 277458 3256
rect 56042 3136 56048 3188
rect 56100 3176 56106 3188
rect 58618 3176 58624 3188
rect 56100 3148 58624 3176
rect 56100 3136 56106 3148
rect 58618 3136 58624 3148
rect 58676 3136 58682 3188
rect 65518 3136 65524 3188
rect 65576 3176 65582 3188
rect 66070 3176 66076 3188
rect 65576 3148 66076 3176
rect 65576 3136 65582 3148
rect 66070 3136 66076 3148
rect 66128 3136 66134 3188
rect 80882 3136 80888 3188
rect 80940 3176 80946 3188
rect 83458 3176 83464 3188
rect 80940 3148 83464 3176
rect 80940 3136 80946 3148
rect 83458 3136 83464 3148
rect 83516 3136 83522 3188
rect 299658 3136 299664 3188
rect 299716 3176 299722 3188
rect 302234 3176 302240 3188
rect 299716 3148 302240 3176
rect 299716 3136 299722 3148
rect 302234 3136 302240 3148
rect 302292 3136 302298 3188
rect 302878 3068 302884 3120
rect 302936 3108 302942 3120
rect 305546 3108 305552 3120
rect 302936 3080 305552 3108
rect 302936 3068 302942 3080
rect 305546 3068 305552 3080
rect 305604 3068 305610 3120
rect 17034 3000 17040 3052
rect 17092 3040 17098 3052
rect 22738 3040 22744 3052
rect 17092 3012 22744 3040
rect 17092 3000 17098 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 29638 3040 29644 3052
rect 27764 3012 29644 3040
rect 27764 3000 27770 3012
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 93946 3000 93952 3052
rect 94004 3040 94010 3052
rect 95050 3040 95056 3052
rect 94004 3012 95056 3040
rect 94004 3000 94010 3012
rect 95050 3000 95056 3012
rect 95108 3000 95114 3052
rect 250438 3000 250444 3052
rect 250496 3040 250502 3052
rect 252370 3040 252376 3052
rect 250496 3012 252376 3040
rect 250496 3000 250502 3012
rect 252370 3000 252376 3012
rect 252428 3000 252434 3052
rect 580994 2864 581000 2916
rect 581052 2904 581058 2916
rect 583018 2904 583024 2916
rect 581052 2876 583024 2904
rect 581052 2864 581058 2876
rect 583018 2864 583024 2876
rect 583076 2864 583082 2916
rect 129366 2116 129372 2168
rect 129424 2156 129430 2168
rect 136634 2156 136640 2168
rect 129424 2128 136640 2156
rect 129424 2116 129430 2128
rect 136634 2116 136640 2128
rect 136692 2116 136698 2168
rect 51350 2048 51356 2100
rect 51408 2088 51414 2100
rect 195238 2088 195244 2100
rect 51408 2060 195244 2088
rect 51408 2048 51414 2060
rect 195238 2048 195244 2060
rect 195296 2048 195302 2100
rect 240778 2048 240784 2100
rect 240836 2088 240842 2100
rect 300762 2088 300768 2100
rect 240836 2060 300768 2088
rect 240836 2048 240842 2060
rect 300762 2048 300768 2060
rect 300820 2048 300826 2100
<< via1 >>
rect 70216 703264 70268 703316
rect 154120 703264 154172 703316
rect 89720 703196 89772 703248
rect 235172 703196 235224 703248
rect 119344 703128 119396 703180
rect 218980 703128 219032 703180
rect 271144 703128 271196 703180
rect 397460 703128 397512 703180
rect 67640 703060 67692 703112
rect 170312 703060 170364 703112
rect 276664 703060 276716 703112
rect 413652 703060 413704 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 84108 702992 84160 703044
rect 202788 702992 202840 703044
rect 268384 702992 268436 703044
rect 462320 702992 462372 703044
rect 101496 702924 101548 702976
rect 300124 702924 300176 702976
rect 61936 702856 61988 702908
rect 364984 702856 365036 702908
rect 116584 702788 116636 702840
rect 429844 702788 429896 702840
rect 24308 702720 24360 702772
rect 86224 702720 86276 702772
rect 99288 702720 99340 702772
rect 478512 702720 478564 702772
rect 79968 702652 80020 702704
rect 494796 702652 494848 702704
rect 8116 702584 8168 702636
rect 96620 702584 96672 702636
rect 106924 702584 106976 702636
rect 527180 702584 527232 702636
rect 57888 702516 57940 702568
rect 582472 702516 582524 702568
rect 66168 702448 66220 702500
rect 559656 702448 559708 702500
rect 71688 700272 71740 700324
rect 105452 700272 105504 700324
rect 269764 700272 269816 700324
rect 283840 700272 283892 700324
rect 286324 700272 286376 700324
rect 332508 700272 332560 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 3424 683136 3476 683188
rect 18604 683136 18656 683188
rect 2780 671032 2832 671084
rect 4804 671032 4856 671084
rect 3424 656888 3476 656940
rect 74540 656888 74592 656940
rect 309784 643084 309836 643136
rect 580172 643084 580224 643136
rect 3516 618264 3568 618316
rect 39304 618264 39356 618316
rect 3516 605820 3568 605872
rect 94780 605820 94832 605872
rect 83464 590656 83516 590708
rect 84108 590656 84160 590708
rect 132592 590656 132644 590708
rect 307024 590656 307076 590708
rect 579804 590656 579856 590708
rect 40040 589908 40092 589960
rect 96712 589908 96764 589960
rect 67732 587120 67784 587172
rect 71688 587120 71740 587172
rect 125600 587120 125652 587172
rect 78128 585760 78180 585812
rect 88340 585760 88392 585812
rect 121736 585760 121788 585812
rect 582564 585760 582616 585812
rect 55128 585148 55180 585200
rect 79324 585148 79376 585200
rect 87512 585148 87564 585200
rect 121460 585148 121512 585200
rect 121736 585148 121788 585200
rect 76288 583788 76340 583840
rect 107660 583788 107712 583840
rect 44088 583720 44140 583772
rect 92480 583720 92532 583772
rect 77208 583108 77260 583160
rect 79968 583108 80020 583160
rect 81808 582564 81860 582616
rect 83464 582564 83516 582616
rect 62028 582428 62080 582480
rect 73804 582428 73856 582480
rect 90272 582428 90324 582480
rect 95884 582428 95936 582480
rect 50988 582360 51040 582412
rect 69940 582360 69992 582412
rect 73528 582360 73580 582412
rect 110420 582360 110472 582412
rect 69664 581068 69716 581120
rect 80244 581068 80296 581120
rect 86592 581068 86644 581120
rect 126980 581068 127032 581120
rect 43996 581000 44048 581052
rect 89812 581000 89864 581052
rect 90548 581000 90600 581052
rect 93768 581000 93820 581052
rect 105544 581000 105596 581052
rect 46848 580252 46900 580304
rect 69664 580660 69716 580712
rect 85488 580660 85540 580712
rect 3332 579640 3384 579692
rect 46848 579640 46900 579692
rect 64696 579640 64748 579692
rect 66536 579640 66588 579692
rect 113364 579640 113416 579692
rect 94780 579572 94832 579624
rect 96804 579572 96856 579624
rect 97540 576852 97592 576904
rect 118700 576852 118752 576904
rect 97908 576716 97960 576768
rect 99196 576716 99248 576768
rect 101496 576716 101548 576768
rect 3424 576104 3476 576156
rect 33140 576104 33192 576156
rect 33140 575492 33192 575544
rect 34428 575492 34480 575544
rect 66444 575492 66496 575544
rect 97632 575424 97684 575476
rect 106924 575424 106976 575476
rect 97448 572704 97500 572756
rect 100852 572704 100904 572756
rect 99288 571956 99340 572008
rect 106924 571956 106976 572008
rect 64788 571344 64840 571396
rect 66720 571344 66772 571396
rect 97080 571344 97132 571396
rect 100024 571344 100076 571396
rect 56508 570596 56560 570648
rect 66628 570596 66680 570648
rect 97908 570596 97960 570648
rect 103428 570596 103480 570648
rect 582656 570596 582708 570648
rect 103428 569236 103480 569288
rect 114652 569236 114704 569288
rect 97908 569168 97960 569220
rect 133880 569168 133932 569220
rect 95884 567808 95936 567860
rect 103520 567808 103572 567860
rect 49608 565836 49660 565888
rect 67640 565836 67692 565888
rect 63408 564408 63460 564460
rect 66812 564408 66864 564460
rect 52368 564340 52420 564392
rect 57888 564340 57940 564392
rect 66536 564340 66588 564392
rect 35808 561688 35860 561740
rect 66812 561688 66864 561740
rect 96804 561688 96856 561740
rect 128360 561688 128412 561740
rect 48228 560260 48280 560312
rect 66812 560260 66864 560312
rect 60648 558900 60700 558952
rect 66812 558900 66864 558952
rect 96804 558900 96856 558952
rect 114560 558900 114612 558952
rect 97172 558696 97224 558748
rect 100760 558696 100812 558748
rect 53656 557540 53708 557592
rect 66812 557540 66864 557592
rect 57888 554752 57940 554804
rect 66720 554752 66772 554804
rect 3516 554004 3568 554056
rect 21364 554004 21416 554056
rect 57244 553392 57296 553444
rect 66812 553392 66864 553444
rect 96988 552032 97040 552084
rect 111800 552032 111852 552084
rect 97908 550604 97960 550656
rect 115940 550604 115992 550656
rect 97080 549312 97132 549364
rect 100116 549312 100168 549364
rect 41328 549244 41380 549296
rect 66812 549244 66864 549296
rect 50896 546456 50948 546508
rect 66536 546456 66588 546508
rect 65984 545096 66036 545148
rect 66168 545096 66220 545148
rect 55036 544348 55088 544400
rect 61936 544348 61988 544400
rect 66352 544348 66404 544400
rect 97356 543736 97408 543788
rect 108304 543736 108356 543788
rect 18604 542988 18656 543040
rect 66168 542988 66220 543040
rect 66628 542988 66680 543040
rect 95148 540880 95200 540932
rect 95516 540880 95568 540932
rect 67456 539860 67508 539912
rect 71780 539860 71832 539912
rect 87604 539792 87656 539844
rect 93860 539792 93912 539844
rect 48136 539588 48188 539640
rect 66628 539588 66680 539640
rect 75184 538840 75236 538892
rect 96896 538840 96948 538892
rect 3424 538228 3476 538280
rect 70952 538228 71004 538280
rect 89720 538228 89772 538280
rect 90180 538228 90232 538280
rect 136640 538228 136692 538280
rect 70952 537548 71004 537600
rect 79324 537548 79376 537600
rect 4804 537480 4856 537532
rect 96620 537480 96672 537532
rect 304264 536800 304316 536852
rect 580172 536800 580224 536852
rect 39304 536732 39356 536784
rect 73436 536732 73488 536784
rect 76564 536732 76616 536784
rect 78312 536596 78364 536648
rect 82176 536596 82228 536648
rect 21364 536052 21416 536104
rect 39856 536052 39908 536104
rect 69388 536052 69440 536104
rect 86684 536052 86736 536104
rect 91008 536052 91060 536104
rect 119344 536052 119396 536104
rect 80152 535780 80204 535832
rect 81348 535780 81400 535832
rect 82084 535440 82136 535492
rect 86224 535440 86276 535492
rect 90364 535440 90416 535492
rect 91836 535440 91888 535492
rect 3424 534080 3476 534132
rect 94504 534080 94556 534132
rect 68928 533332 68980 533384
rect 100024 533332 100076 533384
rect 82084 530612 82136 530664
rect 91192 530612 91244 530664
rect 61936 530544 61988 530596
rect 96804 530544 96856 530596
rect 88340 530136 88392 530188
rect 88892 530136 88944 530188
rect 3516 527824 3568 527876
rect 118700 527824 118752 527876
rect 83464 525036 83516 525088
rect 100852 525036 100904 525088
rect 88248 522248 88300 522300
rect 98000 522248 98052 522300
rect 76564 519528 76616 519580
rect 102232 519528 102284 519580
rect 3516 514768 3568 514820
rect 11704 514768 11756 514820
rect 48228 511232 48280 511284
rect 580172 511232 580224 511284
rect 82912 487772 82964 487824
rect 111064 487772 111116 487824
rect 65984 485052 66036 485104
rect 118792 485052 118844 485104
rect 82176 482264 82228 482316
rect 109684 482264 109736 482316
rect 64696 479476 64748 479528
rect 92572 479476 92624 479528
rect 86868 478116 86920 478168
rect 95332 478116 95384 478168
rect 64696 476756 64748 476808
rect 84200 476756 84252 476808
rect 2964 475668 3016 475720
rect 4068 475668 4120 475720
rect 4804 475668 4856 475720
rect 66076 475328 66128 475380
rect 98644 475328 98696 475380
rect 65984 474036 66036 474088
rect 75920 474036 75972 474088
rect 67732 473968 67784 474020
rect 120172 473968 120224 474020
rect 74448 471248 74500 471300
rect 112720 471248 112772 471300
rect 67732 469820 67784 469872
rect 96712 469820 96764 469872
rect 85580 468460 85632 468512
rect 116124 468460 116176 468512
rect 77116 467100 77168 467152
rect 89720 467100 89772 467152
rect 78680 465672 78732 465724
rect 100116 465672 100168 465724
rect 67824 464312 67876 464364
rect 118976 464312 119028 464364
rect 3240 462340 3292 462392
rect 29644 462340 29696 462392
rect 92480 461592 92532 461644
rect 125876 461592 125928 461644
rect 77208 459688 77260 459740
rect 77944 459688 77996 459740
rect 64788 458804 64840 458856
rect 107016 458804 107068 458856
rect 79324 457444 79376 457496
rect 121644 457444 121696 457496
rect 64788 456016 64840 456068
rect 86960 456016 87012 456068
rect 99196 456016 99248 456068
rect 117412 456016 117464 456068
rect 94504 452548 94556 452600
rect 96712 452548 96764 452600
rect 68468 451868 68520 451920
rect 90364 451868 90416 451920
rect 71872 450508 71924 450560
rect 120356 450508 120408 450560
rect 53656 449148 53708 449200
rect 85672 449148 85724 449200
rect 3148 448536 3200 448588
rect 21364 448536 21416 448588
rect 11704 448468 11756 448520
rect 103520 448468 103572 448520
rect 103704 448468 103756 448520
rect 66168 446360 66220 446412
rect 80336 446360 80388 446412
rect 67640 445136 67692 445188
rect 83096 445136 83148 445188
rect 82820 445000 82872 445052
rect 109040 445000 109092 445052
rect 65892 444728 65944 444780
rect 70492 444728 70544 444780
rect 81624 443640 81676 443692
rect 100760 443640 100812 443692
rect 50988 442212 51040 442264
rect 95240 442212 95292 442264
rect 102140 442008 102192 442060
rect 102784 442008 102836 442060
rect 102784 441600 102836 441652
rect 128452 441600 128504 441652
rect 52368 440852 52420 440904
rect 88708 440852 88760 440904
rect 108120 440308 108172 440360
rect 136732 440308 136784 440360
rect 46756 440240 46808 440292
rect 52368 440240 52420 440292
rect 94136 440240 94188 440292
rect 95148 440240 95200 440292
rect 125784 440240 125836 440292
rect 48228 439492 48280 439544
rect 74724 439492 74776 439544
rect 105544 439492 105596 439544
rect 116216 439492 116268 439544
rect 90088 438880 90140 438932
rect 122932 438880 122984 438932
rect 55036 438132 55088 438184
rect 83740 438132 83792 438184
rect 91008 438132 91060 438184
rect 106096 438132 106148 438184
rect 106648 437520 106700 437572
rect 118884 437520 118936 437572
rect 106096 437452 106148 437504
rect 123024 437452 123076 437504
rect 71136 437384 71188 437436
rect 75184 437384 75236 437436
rect 90456 437384 90508 437436
rect 94228 437384 94280 437436
rect 100116 437384 100168 437436
rect 104624 437384 104676 437436
rect 95240 437112 95292 437164
rect 95884 437112 95936 437164
rect 67088 436704 67140 436756
rect 74632 436704 74684 436756
rect 116032 436704 116084 436756
rect 582380 436704 582432 436756
rect 85120 436568 85172 436620
rect 87604 436568 87656 436620
rect 77392 436432 77444 436484
rect 82084 436432 82136 436484
rect 103796 436160 103848 436212
rect 104624 436160 104676 436212
rect 123484 436160 123536 436212
rect 18604 436092 18656 436144
rect 71136 436092 71188 436144
rect 95884 436092 95936 436144
rect 116032 436092 116084 436144
rect 69112 435208 69164 435260
rect 69940 435208 69992 435260
rect 50988 434800 51040 434852
rect 69112 434800 69164 434852
rect 4804 434732 4856 434784
rect 111800 434800 111852 434852
rect 112628 434800 112680 434852
rect 109684 434732 109736 434784
rect 114100 434732 114152 434784
rect 134524 434732 134576 434784
rect 71780 434528 71832 434580
rect 73022 434528 73074 434580
rect 68652 434188 68704 434240
rect 71780 434188 71832 434240
rect 53748 433984 53800 434036
rect 63224 433984 63276 434036
rect 66352 433984 66404 434036
rect 72608 433780 72660 433832
rect 73988 433712 74040 433764
rect 68284 433644 68336 433696
rect 69204 433644 69256 433696
rect 70860 433644 70912 433696
rect 67456 433236 67508 433288
rect 39948 432556 40000 432608
rect 111064 433780 111116 433832
rect 113180 433780 113232 433832
rect 111616 433644 111668 433696
rect 112812 433644 112864 433696
rect 132500 433304 132552 433356
rect 112812 433236 112864 433288
rect 120264 433236 120316 433288
rect 57520 431944 57572 431996
rect 66812 431944 66864 431996
rect 114744 431944 114796 431996
rect 124220 431944 124272 431996
rect 58900 430584 58952 430636
rect 66812 430584 66864 430636
rect 114744 430584 114796 430636
rect 135260 430584 135312 430636
rect 60556 429224 60608 429276
rect 66260 429224 66312 429276
rect 53656 429156 53708 429208
rect 66812 429156 66864 429208
rect 115388 427796 115440 427848
rect 118792 427796 118844 427848
rect 121552 427796 121604 427848
rect 56416 426436 56468 426488
rect 66812 426436 66864 426488
rect 114100 426436 114152 426488
rect 141424 426436 141476 426488
rect 118792 426368 118844 426420
rect 122840 426368 122892 426420
rect 45468 425688 45520 425740
rect 65892 425688 65944 425740
rect 66536 425688 66588 425740
rect 115848 425076 115900 425128
rect 118792 425076 118844 425128
rect 115848 424328 115900 424380
rect 142160 424328 142212 424380
rect 52368 423648 52420 423700
rect 66628 423648 66680 423700
rect 2780 423580 2832 423632
rect 4804 423580 4856 423632
rect 60740 423444 60792 423496
rect 61936 423444 61988 423496
rect 66812 423444 66864 423496
rect 37188 422900 37240 422952
rect 60740 422900 60792 422952
rect 115848 422900 115900 422952
rect 121644 422900 121696 422952
rect 144184 422900 144236 422952
rect 115848 421948 115900 422000
rect 118976 421948 119028 422000
rect 118976 421540 119028 421592
rect 151084 421540 151136 421592
rect 43996 420928 44048 420980
rect 48228 420928 48280 420980
rect 66812 420928 66864 420980
rect 66996 419568 67048 419620
rect 60464 419500 60516 419552
rect 66812 419500 66864 419552
rect 66812 419364 66864 419416
rect 43904 418140 43956 418192
rect 66812 418208 66864 418260
rect 64144 418140 64196 418192
rect 66996 418140 67048 418192
rect 34244 416780 34296 416832
rect 57244 416780 57296 416832
rect 115848 416780 115900 416832
rect 121644 416780 121696 416832
rect 66720 416712 66772 416764
rect 115204 415692 115256 415744
rect 116216 415692 116268 415744
rect 119344 415352 119396 415404
rect 120172 415352 120224 415404
rect 115848 414876 115900 414928
rect 119344 414876 119396 414928
rect 54852 414060 54904 414112
rect 66720 414060 66772 414112
rect 49516 413992 49568 414044
rect 67732 413992 67784 414044
rect 115204 413992 115256 414044
rect 143540 413992 143592 414044
rect 115848 413924 115900 413976
rect 128360 413924 128412 413976
rect 33048 413244 33100 413296
rect 59268 413244 59320 413296
rect 66260 413244 66312 413296
rect 128360 413244 128412 413296
rect 140780 413244 140832 413296
rect 115848 412020 115900 412072
rect 120356 412020 120408 412072
rect 129740 412020 129792 412072
rect 115848 410524 115900 410576
rect 117504 410524 117556 410576
rect 127072 410524 127124 410576
rect 2872 409844 2924 409896
rect 7564 409844 7616 409896
rect 49608 409844 49660 409896
rect 52276 409844 52328 409896
rect 66812 409844 66864 409896
rect 50804 408484 50856 408536
rect 66628 408484 66680 408536
rect 115848 408484 115900 408536
rect 147680 408484 147732 408536
rect 37096 407056 37148 407108
rect 41236 407056 41288 407108
rect 66812 407124 66864 407176
rect 115848 407124 115900 407176
rect 149060 407124 149112 407176
rect 115572 405628 115624 405680
rect 132592 405628 132644 405680
rect 133788 405628 133840 405680
rect 39856 404948 39908 405000
rect 59084 404948 59136 405000
rect 115848 404948 115900 405000
rect 126980 404948 127032 405000
rect 127440 404948 127492 405000
rect 133788 404948 133840 405000
rect 146300 404948 146352 405000
rect 64788 404336 64840 404388
rect 66812 404336 66864 404388
rect 66352 404268 66404 404320
rect 66904 404268 66956 404320
rect 127440 403588 127492 403640
rect 144920 403588 144972 403640
rect 115848 403248 115900 403300
rect 118608 403248 118660 403300
rect 39856 402976 39908 403028
rect 66352 403044 66404 403096
rect 63316 402976 63368 403028
rect 66812 402976 66864 403028
rect 118608 402228 118660 402280
rect 142804 402228 142856 402280
rect 35624 400868 35676 400920
rect 66444 400868 66496 400920
rect 115020 400392 115072 400444
rect 117504 400392 117556 400444
rect 56508 400188 56560 400240
rect 66812 400188 66864 400240
rect 115664 400188 115716 400240
rect 151820 400188 151872 400240
rect 55036 398828 55088 398880
rect 66812 398828 66864 398880
rect 114560 398080 114612 398132
rect 114928 398080 114980 398132
rect 115848 398080 115900 398132
rect 125692 398080 125744 398132
rect 3424 397468 3476 397520
rect 21456 397468 21508 397520
rect 42616 396720 42668 396772
rect 60648 396720 60700 396772
rect 66812 396720 66864 396772
rect 115848 396720 115900 396772
rect 124128 396720 124180 396772
rect 59084 396108 59136 396160
rect 66812 396108 66864 396160
rect 115848 396040 115900 396092
rect 131120 396040 131172 396092
rect 48044 395292 48096 395344
rect 64696 395292 64748 395344
rect 66812 395292 66864 395344
rect 115848 394680 115900 394732
rect 191104 394680 191156 394732
rect 64604 393320 64656 393372
rect 66812 393320 66864 393372
rect 115572 393320 115624 393372
rect 187700 393320 187752 393372
rect 115848 393116 115900 393168
rect 118700 393116 118752 393168
rect 118700 392028 118752 392080
rect 122840 392028 122892 392080
rect 57704 391960 57756 392012
rect 66812 391960 66864 392012
rect 115848 391960 115900 392012
rect 147772 391960 147824 392012
rect 63408 391280 63460 391332
rect 48136 391212 48188 391264
rect 87972 391008 88024 391060
rect 99472 391008 99524 391060
rect 106648 391008 106700 391060
rect 117412 391212 117464 391264
rect 128360 391212 128412 391264
rect 89904 390940 89956 390992
rect 92940 390940 92992 390992
rect 112168 390668 112220 390720
rect 112720 390668 112772 390720
rect 88248 390260 88300 390312
rect 88984 390260 89036 390312
rect 67640 390124 67692 390176
rect 68790 390124 68842 390176
rect 41328 389852 41380 389904
rect 53840 389852 53892 389904
rect 21364 389784 21416 389836
rect 99196 389784 99248 389836
rect 100760 389784 100812 389836
rect 104808 389784 104860 389836
rect 114928 389784 114980 389836
rect 53840 389172 53892 389224
rect 54760 389172 54812 389224
rect 83004 389172 83056 389224
rect 65984 389104 66036 389156
rect 72516 389104 72568 389156
rect 101680 389104 101732 389156
rect 106648 389104 106700 389156
rect 110144 389104 110196 389156
rect 121460 389104 121512 389156
rect 46664 388424 46716 388476
rect 65984 388424 66036 388476
rect 91100 388424 91152 388476
rect 100024 388424 100076 388476
rect 103704 388424 103756 388476
rect 232504 388424 232556 388476
rect 93400 388288 93452 388340
rect 95884 388288 95936 388340
rect 85396 387812 85448 387864
rect 90364 387812 90416 387864
rect 44088 387744 44140 387796
rect 55128 387744 55180 387796
rect 73988 387744 74040 387796
rect 74264 387744 74316 387796
rect 75276 387744 75328 387796
rect 79876 387744 79928 387796
rect 81532 387744 81584 387796
rect 120724 387744 120776 387796
rect 121460 387744 121512 387796
rect 76564 387608 76616 387660
rect 80060 387608 80112 387660
rect 86868 387064 86920 387116
rect 120724 387064 120776 387116
rect 69020 386996 69072 387048
rect 69756 386996 69808 387048
rect 77300 386996 77352 387048
rect 78036 386996 78088 387048
rect 93860 386996 93912 387048
rect 94780 386996 94832 387048
rect 111800 386996 111852 387048
rect 112260 386996 112312 387048
rect 46848 386316 46900 386368
rect 96620 386316 96672 386368
rect 97908 386316 97960 386368
rect 105176 386316 105228 386368
rect 133880 386316 133932 386368
rect 136640 386316 136692 386368
rect 80888 386248 80940 386300
rect 81348 386248 81400 386300
rect 115940 386248 115992 386300
rect 108672 384956 108724 385008
rect 125876 384956 125928 385008
rect 126888 384956 126940 385008
rect 101404 384344 101456 384396
rect 113180 384344 113232 384396
rect 57888 384276 57940 384328
rect 104900 384276 104952 384328
rect 35808 383596 35860 383648
rect 91836 383596 91888 383648
rect 77392 382984 77444 383036
rect 106924 382984 106976 383036
rect 97908 382916 97960 382968
rect 126980 382916 127032 382968
rect 91192 382440 91244 382492
rect 91836 382440 91888 382492
rect 34428 382168 34480 382220
rect 96712 382168 96764 382220
rect 96712 381556 96764 381608
rect 117412 381556 117464 381608
rect 73068 381488 73120 381540
rect 77484 381488 77536 381540
rect 107476 381488 107528 381540
rect 139400 381488 139452 381540
rect 38568 380128 38620 380180
rect 69112 380128 69164 380180
rect 93216 380128 93268 380180
rect 115940 380128 115992 380180
rect 103520 378836 103572 378888
rect 138020 378836 138072 378888
rect 21456 378768 21508 378820
rect 114468 378768 114520 378820
rect 116216 378768 116268 378820
rect 95148 378224 95200 378276
rect 102324 378224 102376 378276
rect 97908 377408 97960 377460
rect 120264 377408 120316 377460
rect 92388 376048 92440 376100
rect 97540 376048 97592 376100
rect 104256 376048 104308 376100
rect 123024 376048 123076 376100
rect 48136 375980 48188 376032
rect 76012 375980 76064 376032
rect 83464 375980 83516 376032
rect 105544 375980 105596 376032
rect 101956 374620 102008 374672
rect 113456 374620 113508 374672
rect 93952 373260 94004 373312
rect 124312 373260 124364 373312
rect 3424 371220 3476 371272
rect 106096 371220 106148 371272
rect 116124 371152 116176 371204
rect 93860 370472 93912 370524
rect 126244 370472 126296 370524
rect 86776 367752 86828 367804
rect 117320 367752 117372 367804
rect 90364 366324 90416 366376
rect 117964 366324 118016 366376
rect 88984 364964 89036 365016
rect 121460 364964 121512 365016
rect 93124 363604 93176 363656
rect 119068 363604 119120 363656
rect 95056 362176 95108 362228
rect 118884 362176 118936 362228
rect 89444 359456 89496 359508
rect 124404 359456 124456 359508
rect 3332 358708 3384 358760
rect 17224 358708 17276 358760
rect 84108 356668 84160 356720
rect 112444 356668 112496 356720
rect 85580 353948 85632 354000
rect 104164 353948 104216 354000
rect 113824 349120 113876 349172
rect 260104 349120 260156 349172
rect 93124 346400 93176 346452
rect 93676 346400 93728 346452
rect 272064 346400 272116 346452
rect 3332 345040 3384 345092
rect 11704 345040 11756 345092
rect 141424 345040 141476 345092
rect 270592 345040 270644 345092
rect 123484 343680 123536 343732
rect 269120 343680 269172 343732
rect 73804 343612 73856 343664
rect 240140 343612 240192 343664
rect 66996 342252 67048 342304
rect 67456 342252 67508 342304
rect 261484 342252 261536 342304
rect 151084 340960 151136 341012
rect 271972 340960 272024 341012
rect 75276 340892 75328 340944
rect 253296 340892 253348 340944
rect 142804 339532 142856 339584
rect 240416 339532 240468 339584
rect 45284 339464 45336 339516
rect 81440 339464 81492 339516
rect 83556 339464 83608 339516
rect 266452 339464 266504 339516
rect 81440 338716 81492 338768
rect 251180 338716 251232 338768
rect 97816 338104 97868 338156
rect 242164 338104 242216 338156
rect 69664 336812 69716 336864
rect 246396 336812 246448 336864
rect 53564 336744 53616 336796
rect 249800 336744 249852 336796
rect 39672 335996 39724 336048
rect 74632 335996 74684 336048
rect 238024 335996 238076 336048
rect 92388 335316 92440 335368
rect 191196 335316 191248 335368
rect 95240 334568 95292 334620
rect 122932 334568 122984 334620
rect 123852 334568 123904 334620
rect 123852 334024 123904 334076
rect 233884 334024 233936 334076
rect 88248 333956 88300 334008
rect 240784 333956 240836 334008
rect 89720 333208 89772 333260
rect 120172 333208 120224 333260
rect 120172 332596 120224 332648
rect 247684 332596 247736 332648
rect 80704 331304 80756 331356
rect 81256 331304 81308 331356
rect 241520 331304 241572 331356
rect 101496 331236 101548 331288
rect 101956 331236 102008 331288
rect 269212 331236 269264 331288
rect 42708 330488 42760 330540
rect 66996 330488 67048 330540
rect 99288 329876 99340 329928
rect 226984 329876 227036 329928
rect 53472 329808 53524 329860
rect 53656 329808 53708 329860
rect 267832 329808 267884 329860
rect 89720 329060 89772 329112
rect 123024 329060 123076 329112
rect 259644 329060 259696 329112
rect 100208 328448 100260 328500
rect 100668 328448 100720 328500
rect 242900 328448 242952 328500
rect 63224 328380 63276 328432
rect 63408 328380 63460 328432
rect 38476 328176 38528 328228
rect 39856 328176 39908 328228
rect 39856 327700 39908 327752
rect 67548 327700 67600 327752
rect 80244 327700 80296 327752
rect 89720 327700 89772 327752
rect 115204 327156 115256 327208
rect 246488 327156 246540 327208
rect 63408 327088 63460 327140
rect 266544 327088 266596 327140
rect 108856 326340 108908 326392
rect 116124 326340 116176 326392
rect 116124 325728 116176 325780
rect 254032 325728 254084 325780
rect 78036 325660 78088 325712
rect 84108 325660 84160 325712
rect 255412 325660 255464 325712
rect 129004 324912 129056 324964
rect 151084 324912 151136 324964
rect 192484 324368 192536 324420
rect 208676 324368 208728 324420
rect 49516 324300 49568 324352
rect 258172 324300 258224 324352
rect 291844 324300 291896 324352
rect 580172 324300 580224 324352
rect 96528 323552 96580 323604
rect 136732 323552 136784 323604
rect 260932 323552 260984 323604
rect 75368 322940 75420 322992
rect 75828 322940 75880 322992
rect 249064 322940 249116 322992
rect 119344 321920 119396 321972
rect 123484 321920 123536 321972
rect 88156 321716 88208 321768
rect 91192 321716 91244 321768
rect 125508 321648 125560 321700
rect 259552 321648 259604 321700
rect 108856 321580 108908 321632
rect 111892 321580 111944 321632
rect 265164 321580 265216 321632
rect 4804 320832 4856 320884
rect 18604 320832 18656 320884
rect 113916 320628 113968 320680
rect 114468 320628 114520 320680
rect 118884 320220 118936 320272
rect 267740 320220 267792 320272
rect 56232 320152 56284 320204
rect 88156 320152 88208 320204
rect 114468 320152 114520 320204
rect 263600 320152 263652 320204
rect 3884 319200 3936 319252
rect 4804 319200 4856 319252
rect 151084 318860 151136 318912
rect 250444 318860 250496 318912
rect 41144 318792 41196 318844
rect 63500 318792 63552 318844
rect 64144 318792 64196 318844
rect 72976 318792 73028 318844
rect 251824 318792 251876 318844
rect 100116 318112 100168 318164
rect 111892 318112 111944 318164
rect 63500 318044 63552 318096
rect 250536 318044 250588 318096
rect 111892 317432 111944 317484
rect 255504 317432 255556 317484
rect 63224 316684 63276 316736
rect 72884 316684 72936 316736
rect 256700 316684 256752 316736
rect 84200 316004 84252 316056
rect 85304 316004 85356 316056
rect 264980 316004 265032 316056
rect 106096 315256 106148 315308
rect 137100 315256 137152 315308
rect 134616 314712 134668 314764
rect 252744 314712 252796 314764
rect 136732 314644 136784 314696
rect 137100 314644 137152 314696
rect 258356 314644 258408 314696
rect 117780 313896 117832 313948
rect 125784 313896 125836 313948
rect 260840 313896 260892 313948
rect 71688 313284 71740 313336
rect 75184 313284 75236 313336
rect 75828 313284 75880 313336
rect 82912 313284 82964 313336
rect 117320 313284 117372 313336
rect 117780 313284 117832 313336
rect 186964 313284 187016 313336
rect 266636 313284 266688 313336
rect 160744 311924 160796 311976
rect 255320 311924 255372 311976
rect 144184 311856 144236 311908
rect 258080 311856 258132 311908
rect 94596 311108 94648 311160
rect 114468 311108 114520 311160
rect 160836 310564 160888 310616
rect 261024 310564 261076 310616
rect 114468 310496 114520 310548
rect 259736 310496 259788 310548
rect 78128 310428 78180 310480
rect 78588 310428 78640 310480
rect 180064 309816 180116 309868
rect 188344 309816 188396 309868
rect 78128 309748 78180 309800
rect 266360 309748 266412 309800
rect 189724 309136 189776 309188
rect 252836 309136 252888 309188
rect 79876 308388 79928 308440
rect 109316 308388 109368 308440
rect 233884 308388 233936 308440
rect 243912 308388 243964 308440
rect 245016 308388 245068 308440
rect 256976 308388 257028 308440
rect 123484 307844 123536 307896
rect 218244 307844 218296 307896
rect 109316 307776 109368 307828
rect 262496 307776 262548 307828
rect 123116 307708 123168 307760
rect 124220 307708 124272 307760
rect 240784 307708 240836 307760
rect 244464 307708 244516 307760
rect 250444 307708 250496 307760
rect 254124 307708 254176 307760
rect 250536 307640 250588 307692
rect 255596 307640 255648 307692
rect 176016 306416 176068 306468
rect 215944 306416 215996 306468
rect 100668 306348 100720 306400
rect 123116 306348 123168 306400
rect 137284 306348 137336 306400
rect 236368 306348 236420 306400
rect 246396 306348 246448 306400
rect 250352 306348 250404 306400
rect 122840 306280 122892 306332
rect 160744 306280 160796 306332
rect 249064 306008 249116 306060
rect 254216 306008 254268 306060
rect 84108 305600 84160 305652
rect 87052 305600 87104 305652
rect 111064 305600 111116 305652
rect 122840 305600 122892 305652
rect 214564 305600 214616 305652
rect 259460 305600 259512 305652
rect 126244 305396 126296 305448
rect 128544 305396 128596 305448
rect 232504 305124 232556 305176
rect 239864 305124 239916 305176
rect 182824 305056 182876 305108
rect 197268 305056 197320 305108
rect 96436 304988 96488 305040
rect 100208 304988 100260 305040
rect 155408 304988 155460 305040
rect 214196 304988 214248 305040
rect 260104 304988 260156 305040
rect 263876 304988 263928 305040
rect 62028 304920 62080 304972
rect 66904 304920 66956 304972
rect 160836 304920 160888 304972
rect 246304 304444 246356 304496
rect 249708 304444 249760 304496
rect 60372 304240 60424 304292
rect 151084 304240 151136 304292
rect 184204 303696 184256 303748
rect 160744 303628 160796 303680
rect 205456 303696 205508 303748
rect 211252 303696 211304 303748
rect 245108 303696 245160 303748
rect 289084 303696 289136 303748
rect 247408 303628 247460 303680
rect 248328 303628 248380 303680
rect 252652 303628 252704 303680
rect 336004 303628 336056 303680
rect 200304 303560 200356 303612
rect 201132 303560 201184 303612
rect 242808 302880 242860 302932
rect 273260 302880 273312 302932
rect 69756 302268 69808 302320
rect 75828 302268 75880 302320
rect 184296 302268 184348 302320
rect 200212 302268 200264 302320
rect 56508 302200 56560 302252
rect 120908 302200 120960 302252
rect 173164 302200 173216 302252
rect 249156 302200 249208 302252
rect 251824 302200 251876 302252
rect 252928 302200 252980 302252
rect 240140 302132 240192 302184
rect 240968 302132 241020 302184
rect 86868 301452 86920 301504
rect 100116 301452 100168 301504
rect 118056 301452 118108 301504
rect 142804 301452 142856 301504
rect 65984 301248 66036 301300
rect 69020 301248 69072 301300
rect 241336 301112 241388 301164
rect 262588 301112 262640 301164
rect 240784 301044 240836 301096
rect 160836 300908 160888 300960
rect 196348 300908 196400 300960
rect 66076 300840 66128 300892
rect 141424 300840 141476 300892
rect 53748 300772 53800 300824
rect 193496 300772 193548 300824
rect 250628 300976 250680 301028
rect 248052 300908 248104 300960
rect 193680 300092 193732 300144
rect 270500 300840 270552 300892
rect 253204 299684 253256 299736
rect 255688 299548 255740 299600
rect 274640 299548 274692 299600
rect 134524 299480 134576 299532
rect 193588 299480 193640 299532
rect 255872 299480 255924 299532
rect 282184 299480 282236 299532
rect 255780 299412 255832 299464
rect 263692 299412 263744 299464
rect 255688 299344 255740 299396
rect 258264 299344 258316 299396
rect 259368 299344 259420 299396
rect 85764 299072 85816 299124
rect 86776 299072 86828 299124
rect 100024 299004 100076 299056
rect 105636 299004 105688 299056
rect 186320 298868 186372 298920
rect 191748 298868 191800 298920
rect 259368 298732 259420 298784
rect 280896 298732 280948 298784
rect 71044 298596 71096 298648
rect 72608 298596 72660 298648
rect 86776 298120 86828 298172
rect 139492 298120 139544 298172
rect 263692 298120 263744 298172
rect 268476 298120 268528 298172
rect 298744 298120 298796 298172
rect 580172 298120 580224 298172
rect 255780 298052 255832 298104
rect 269212 298052 269264 298104
rect 270408 298052 270460 298104
rect 261484 297984 261536 298036
rect 262220 297984 262272 298036
rect 255688 297372 255740 297424
rect 262128 297372 262180 297424
rect 270408 297372 270460 297424
rect 282092 297372 282144 297424
rect 282184 297372 282236 297424
rect 317420 297372 317472 297424
rect 255688 296624 255740 296676
rect 267832 296624 267884 296676
rect 269028 296624 269080 296676
rect 57612 295944 57664 295996
rect 78588 295944 78640 295996
rect 191196 295944 191248 295996
rect 269028 295944 269080 295996
rect 287060 295944 287112 295996
rect 255412 295808 255464 295860
rect 255780 295808 255832 295860
rect 78680 295332 78732 295384
rect 79968 295332 80020 295384
rect 110604 295332 110656 295384
rect 170404 295332 170456 295384
rect 191748 295332 191800 295384
rect 255412 295332 255464 295384
rect 259368 295332 259420 295384
rect 259644 295332 259696 295384
rect 120816 294584 120868 294636
rect 191104 294584 191156 294636
rect 256792 294040 256844 294092
rect 257344 294040 257396 294092
rect 39856 293972 39908 294024
rect 75184 293972 75236 294024
rect 75368 293972 75420 294024
rect 93768 293972 93820 294024
rect 124864 293972 124916 294024
rect 191656 293972 191708 294024
rect 255412 293972 255464 294024
rect 263692 293972 263744 294024
rect 153108 293904 153160 293956
rect 191748 293904 191800 293956
rect 255688 293904 255740 293956
rect 263876 293904 263928 293956
rect 255412 293836 255464 293888
rect 262220 293836 262272 293888
rect 95884 293224 95936 293276
rect 104992 293224 105044 293276
rect 125508 293224 125560 293276
rect 151820 293224 151872 293276
rect 153108 293224 153160 293276
rect 41328 292612 41380 292664
rect 77852 292612 77904 292664
rect 78036 292612 78088 292664
rect 3516 292544 3568 292596
rect 14464 292544 14516 292596
rect 60464 292544 60516 292596
rect 60648 292544 60700 292596
rect 191472 292544 191524 292596
rect 255412 292068 255464 292120
rect 256976 292068 257028 292120
rect 159364 291864 159416 291916
rect 189816 291864 189868 291916
rect 77760 291796 77812 291848
rect 78128 291796 78180 291848
rect 85580 291796 85632 291848
rect 116032 291796 116084 291848
rect 120908 291796 120960 291848
rect 191104 291796 191156 291848
rect 37096 291320 37148 291372
rect 72424 291320 72476 291372
rect 41236 291252 41288 291304
rect 77760 291252 77812 291304
rect 72056 291184 72108 291236
rect 73068 291184 73120 291236
rect 131764 291184 131816 291236
rect 255688 291116 255740 291168
rect 271972 291116 272024 291168
rect 255412 290844 255464 290896
rect 258172 290844 258224 290896
rect 76196 290708 76248 290760
rect 76748 290708 76800 290760
rect 162124 290436 162176 290488
rect 192484 290436 192536 290488
rect 89536 289892 89588 289944
rect 120908 289892 120960 289944
rect 39764 289824 39816 289876
rect 76196 289824 76248 289876
rect 81992 289824 82044 289876
rect 82728 289824 82780 289876
rect 112076 289824 112128 289876
rect 191748 289824 191800 289876
rect 46756 289756 46808 289808
rect 52184 289756 52236 289808
rect 255688 289756 255740 289808
rect 270592 289756 270644 289808
rect 255412 289688 255464 289740
rect 260932 289688 260984 289740
rect 56324 288464 56376 288516
rect 83004 288464 83056 288516
rect 83464 288464 83516 288516
rect 101588 288464 101640 288516
rect 113824 288464 113876 288516
rect 52184 288396 52236 288448
rect 79968 288396 80020 288448
rect 95240 288396 95292 288448
rect 96528 288396 96580 288448
rect 109132 288396 109184 288448
rect 116584 288396 116636 288448
rect 191748 288396 191800 288448
rect 88616 288328 88668 288380
rect 89628 288328 89680 288380
rect 179420 288328 179472 288380
rect 190828 288328 190880 288380
rect 255412 288328 255464 288380
rect 269120 288328 269172 288380
rect 255688 288260 255740 288312
rect 265164 288260 265216 288312
rect 78680 287716 78732 287768
rect 79140 287716 79192 287768
rect 85672 287716 85724 287768
rect 86316 287716 86368 287768
rect 11704 287648 11756 287700
rect 34520 287648 34572 287700
rect 58992 287648 59044 287700
rect 71688 287648 71740 287700
rect 74540 287648 74592 287700
rect 110512 287648 110564 287700
rect 119344 287648 119396 287700
rect 169024 287648 169076 287700
rect 187056 287648 187108 287700
rect 93676 287104 93728 287156
rect 102232 287104 102284 287156
rect 34520 287036 34572 287088
rect 35716 287036 35768 287088
rect 70952 287036 71004 287088
rect 91468 287036 91520 287088
rect 110512 287036 110564 287088
rect 82912 286968 82964 287020
rect 85488 286968 85540 287020
rect 255504 286968 255556 287020
rect 265072 286968 265124 287020
rect 74080 286900 74132 286952
rect 76564 286900 76616 286952
rect 77392 286356 77444 286408
rect 77944 286356 77996 286408
rect 3424 286288 3476 286340
rect 15844 286288 15896 286340
rect 93032 286288 93084 286340
rect 93768 286288 93820 286340
rect 45376 285812 45428 285864
rect 75276 285812 75328 285864
rect 72516 285744 72568 285796
rect 148324 285744 148376 285796
rect 165528 285744 165580 285796
rect 191748 285744 191800 285796
rect 95608 285676 95660 285728
rect 107568 285676 107620 285728
rect 115848 285676 115900 285728
rect 190368 285676 190420 285728
rect 63224 285608 63276 285660
rect 64144 285608 64196 285660
rect 43904 284928 43956 284980
rect 60740 284928 60792 284980
rect 67548 284928 67600 284980
rect 68652 284928 68704 284980
rect 98368 284928 98420 284980
rect 151176 284928 151228 284980
rect 178776 284928 178828 284980
rect 255596 284928 255648 284980
rect 267740 284928 267792 284980
rect 255412 284520 255464 284572
rect 259552 284520 259604 284572
rect 52092 284316 52144 284368
rect 76656 284316 76708 284368
rect 173256 284316 173308 284368
rect 191748 284316 191800 284368
rect 255412 284248 255464 284300
rect 261024 284248 261076 284300
rect 75046 283704 75098 283756
rect 75276 283704 75328 283756
rect 39948 283568 40000 283620
rect 52460 283568 52512 283620
rect 91376 283568 91428 283620
rect 93124 283568 93176 283620
rect 99472 283568 99524 283620
rect 97908 283432 97960 283484
rect 98460 283432 98512 283484
rect 47860 282956 47912 283008
rect 69112 283092 69164 283144
rect 69848 283092 69900 283144
rect 68652 283024 68704 283076
rect 80244 283024 80296 283076
rect 68376 282956 68428 283008
rect 69204 282956 69256 283008
rect 69756 282956 69808 283008
rect 64512 282208 64564 282260
rect 84752 282956 84804 283008
rect 106372 282888 106424 282940
rect 126244 282888 126296 282940
rect 191748 282888 191800 282940
rect 98920 282820 98972 282872
rect 99380 282820 99432 282872
rect 255504 282820 255556 282872
rect 266636 282820 266688 282872
rect 255412 282752 255464 282804
rect 258356 282752 258408 282804
rect 52460 282140 52512 282192
rect 53656 282140 53708 282192
rect 69020 282140 69072 282192
rect 187148 282140 187200 282192
rect 120908 281528 120960 281580
rect 128452 281528 128504 281580
rect 48136 281460 48188 281512
rect 53104 281460 53156 281512
rect 98368 281460 98420 281512
rect 189724 281460 189776 281512
rect 255412 281460 255464 281512
rect 262496 281460 262548 281512
rect 99380 280780 99432 280832
rect 113364 280780 113416 280832
rect 134616 280780 134668 280832
rect 3424 280168 3476 280220
rect 67548 280168 67600 280220
rect 169116 280168 169168 280220
rect 191564 280168 191616 280220
rect 255504 280168 255556 280220
rect 271880 280168 271932 280220
rect 108948 280100 109000 280152
rect 186964 280100 187016 280152
rect 255320 280100 255372 280152
rect 263784 280100 263836 280152
rect 255412 280032 255464 280084
rect 259736 280032 259788 280084
rect 57888 279556 57940 279608
rect 66076 279556 66128 279608
rect 66628 279556 66680 279608
rect 4804 279420 4856 279472
rect 32864 279420 32916 279472
rect 60372 279420 60424 279472
rect 66812 279420 66864 279472
rect 99472 279420 99524 279472
rect 107844 279420 107896 279472
rect 175188 279420 175240 279472
rect 187700 279420 187752 279472
rect 191748 279488 191800 279540
rect 108304 279216 108356 279268
rect 108948 279216 109000 279268
rect 142988 278740 143040 278792
rect 175188 278740 175240 278792
rect 128452 278672 128504 278724
rect 191748 278672 191800 278724
rect 259368 278672 259420 278724
rect 259828 278672 259880 278724
rect 255412 278468 255464 278520
rect 258080 278468 258132 278520
rect 50988 277992 51040 278044
rect 59176 277992 59228 278044
rect 66812 277992 66864 278044
rect 102048 277992 102100 278044
rect 131212 277992 131264 278044
rect 151084 277992 151136 278044
rect 255412 277448 255464 277500
rect 258172 277448 258224 277500
rect 162216 277380 162268 277432
rect 191656 277380 191708 277432
rect 66076 277312 66128 277364
rect 68284 277312 68336 277364
rect 113824 276700 113876 276752
rect 127164 276700 127216 276752
rect 100024 276632 100076 276684
rect 118976 276632 119028 276684
rect 144828 276632 144880 276684
rect 182824 276632 182876 276684
rect 102140 276292 102192 276344
rect 102784 276292 102836 276344
rect 255504 276088 255556 276140
rect 263600 276088 263652 276140
rect 43904 276020 43956 276072
rect 52460 276020 52512 276072
rect 66812 276020 66864 276072
rect 136548 276020 136600 276072
rect 144184 276020 144236 276072
rect 255320 276020 255372 276072
rect 265256 276020 265308 276072
rect 63408 275952 63460 276004
rect 66904 275952 66956 276004
rect 255412 275952 255464 276004
rect 264980 275952 265032 276004
rect 261484 275340 261536 275392
rect 269120 275340 269172 275392
rect 100760 275272 100812 275324
rect 142160 275272 142212 275324
rect 142896 275272 142948 275324
rect 155224 275272 155276 275324
rect 188344 275272 188396 275324
rect 188988 274728 189040 274780
rect 191656 274728 191708 274780
rect 57796 274660 57848 274712
rect 63408 274660 63460 274712
rect 130568 274660 130620 274712
rect 168288 274660 168340 274712
rect 191748 274660 191800 274712
rect 58900 274592 58952 274644
rect 65892 274592 65944 274644
rect 66536 274592 66588 274644
rect 141424 274592 141476 274644
rect 193128 274592 193180 274644
rect 255412 274592 255464 274644
rect 260840 274592 260892 274644
rect 58900 274116 58952 274168
rect 59268 274116 59320 274168
rect 100760 273980 100812 274032
rect 128452 273980 128504 274032
rect 100852 273912 100904 273964
rect 135260 273912 135312 273964
rect 136548 273912 136600 273964
rect 255964 273912 256016 273964
rect 582472 273912 582524 273964
rect 128452 273844 128504 273896
rect 129004 273844 129056 273896
rect 104164 273164 104216 273216
rect 116860 273164 116912 273216
rect 116860 272484 116912 272536
rect 169116 272484 169168 272536
rect 62856 272076 62908 272128
rect 63224 272076 63276 272128
rect 66812 272076 66864 272128
rect 171784 271940 171836 271992
rect 191196 271940 191248 271992
rect 255504 271940 255556 271992
rect 269212 271940 269264 271992
rect 109684 271872 109736 271924
rect 112260 271872 112312 271924
rect 122840 271872 122892 271924
rect 160928 271872 160980 271924
rect 163596 271872 163648 271924
rect 191748 271872 191800 271924
rect 255412 271872 255464 271924
rect 265072 271872 265124 271924
rect 267004 271872 267056 271924
rect 580172 271872 580224 271924
rect 54944 271804 54996 271856
rect 56416 271804 56468 271856
rect 66812 271804 66864 271856
rect 255320 271804 255372 271856
rect 266544 271804 266596 271856
rect 255504 271600 255556 271652
rect 259460 271600 259512 271652
rect 101680 271124 101732 271176
rect 103428 271124 103480 271176
rect 130384 271124 130436 271176
rect 173164 271124 173216 271176
rect 100760 269900 100812 269952
rect 104440 269900 104492 269952
rect 135904 269764 135956 269816
rect 188436 269764 188488 269816
rect 255596 269764 255648 269816
rect 273352 269764 273404 269816
rect 103980 269084 104032 269136
rect 106832 269084 106884 269136
rect 135904 269084 135956 269136
rect 181444 269084 181496 269136
rect 191748 269084 191800 269136
rect 255412 269084 255464 269136
rect 260932 269084 260984 269136
rect 104900 269016 104952 269068
rect 109592 269016 109644 269068
rect 131764 269016 131816 269068
rect 192484 269016 192536 269068
rect 116676 268880 116728 268932
rect 118884 268880 118936 268932
rect 100760 268404 100812 268456
rect 104900 268404 104952 268456
rect 52368 268336 52420 268388
rect 66168 268336 66220 268388
rect 100852 268336 100904 268388
rect 113272 268336 113324 268388
rect 113916 268336 113968 268388
rect 178776 267724 178828 267776
rect 191656 267724 191708 267776
rect 255504 267724 255556 267776
rect 261116 267724 261168 267776
rect 53748 267656 53800 267708
rect 66260 267656 66312 267708
rect 255412 267656 255464 267708
rect 285680 267656 285732 267708
rect 104440 266976 104492 267028
rect 119436 266976 119488 267028
rect 141516 266976 141568 267028
rect 180156 266976 180208 267028
rect 255412 266976 255464 267028
rect 262220 266976 262272 267028
rect 3056 266364 3108 266416
rect 11704 266364 11756 266416
rect 66812 266364 66864 266416
rect 115388 266364 115440 266416
rect 120908 266364 120960 266416
rect 177396 266364 177448 266416
rect 191472 266364 191524 266416
rect 37188 266296 37240 266348
rect 50344 266296 50396 266348
rect 149060 266296 149112 266348
rect 162216 266296 162268 266348
rect 255320 266296 255372 266348
rect 276020 266296 276072 266348
rect 100116 265616 100168 265668
rect 107660 265616 107712 265668
rect 133788 265616 133840 265668
rect 149060 265616 149112 265668
rect 159456 265616 159508 265668
rect 185584 265616 185636 265668
rect 255964 265616 256016 265668
rect 583208 265616 583260 265668
rect 60648 265140 60700 265192
rect 66812 265140 66864 265192
rect 100852 264936 100904 264988
rect 133144 264936 133196 264988
rect 133788 264936 133840 264988
rect 182824 264936 182876 264988
rect 191748 264936 191800 264988
rect 41144 264188 41196 264240
rect 66628 264188 66680 264240
rect 100760 264188 100812 264240
rect 127072 264188 127124 264240
rect 255412 263644 255464 263696
rect 262220 263644 262272 263696
rect 36544 263576 36596 263628
rect 41144 263576 41196 263628
rect 100760 263576 100812 263628
rect 120080 263576 120132 263628
rect 147588 263576 147640 263628
rect 155316 263576 155368 263628
rect 191012 263576 191064 263628
rect 115020 263508 115072 263560
rect 118792 263508 118844 263560
rect 148324 263508 148376 263560
rect 255412 263508 255464 263560
rect 262312 263508 262364 263560
rect 100760 262896 100812 262948
rect 115020 262896 115072 262948
rect 33968 262828 34020 262880
rect 60740 262828 60792 262880
rect 66904 262828 66956 262880
rect 104164 262828 104216 262880
rect 124404 262828 124456 262880
rect 147588 262828 147640 262880
rect 174544 262828 174596 262880
rect 268384 262828 268436 262880
rect 580264 262828 580316 262880
rect 4804 262216 4856 262268
rect 33968 262216 34020 262268
rect 34336 262216 34388 262268
rect 185584 262216 185636 262268
rect 191012 262216 191064 262268
rect 63132 261536 63184 261588
rect 68284 261536 68336 261588
rect 56416 261468 56468 261520
rect 66720 261468 66772 261520
rect 100760 261468 100812 261520
rect 104808 261468 104860 261520
rect 109224 261468 109276 261520
rect 134524 261468 134576 261520
rect 268476 261468 268528 261520
rect 302240 261468 302292 261520
rect 104256 261060 104308 261112
rect 108304 261060 108356 261112
rect 49516 260788 49568 260840
rect 66444 260788 66496 260840
rect 113180 260720 113232 260772
rect 115204 260720 115256 260772
rect 45468 260108 45520 260160
rect 49516 260108 49568 260160
rect 135168 260108 135220 260160
rect 144920 260108 144972 260160
rect 182916 260108 182968 260160
rect 271788 260108 271840 260160
rect 582748 260108 582800 260160
rect 100852 259428 100904 259480
rect 133972 259428 134024 259480
rect 135168 259428 135220 259480
rect 188252 259428 188304 259480
rect 191748 259428 191800 259480
rect 255412 259428 255464 259480
rect 260840 259428 260892 259480
rect 100760 258748 100812 258800
rect 136732 258748 136784 258800
rect 266636 258748 266688 258800
rect 307024 258748 307076 258800
rect 100852 258680 100904 258732
rect 118056 258680 118108 258732
rect 133788 258680 133840 258732
rect 173348 258680 173400 258732
rect 267924 258680 267976 258732
rect 583300 258680 583352 258732
rect 45560 258136 45612 258188
rect 46204 258136 46256 258188
rect 66260 258136 66312 258188
rect 100852 258136 100904 258188
rect 177304 258136 177356 258188
rect 190644 258136 190696 258188
rect 42708 258068 42760 258120
rect 66352 258068 66404 258120
rect 100760 258068 100812 258120
rect 175924 258068 175976 258120
rect 190552 258068 190604 258120
rect 255412 258068 255464 258120
rect 266636 258068 266688 258120
rect 33048 258000 33100 258052
rect 45560 258000 45612 258052
rect 66260 258000 66312 258052
rect 68192 258000 68244 258052
rect 100852 258000 100904 258052
rect 125508 258000 125560 258052
rect 190460 258000 190512 258052
rect 193404 258000 193456 258052
rect 262680 258000 262732 258052
rect 304264 258000 304316 258052
rect 255412 257388 255464 257440
rect 262680 257388 262732 257440
rect 52276 257320 52328 257372
rect 66628 257320 66680 257372
rect 110420 257320 110472 257372
rect 130476 257320 130528 257372
rect 146944 257320 146996 257372
rect 176016 257320 176068 257372
rect 255688 257320 255740 257372
rect 583484 257320 583536 257372
rect 104348 256708 104400 256760
rect 110420 256708 110472 256760
rect 125508 256708 125560 256760
rect 127072 256708 127124 256760
rect 173164 256708 173216 256760
rect 191748 256708 191800 256760
rect 50804 256640 50856 256692
rect 66812 256640 66864 256692
rect 255504 256640 255556 256692
rect 258356 256640 258408 256692
rect 582840 256640 582892 256692
rect 100852 255960 100904 256012
rect 113180 255960 113232 256012
rect 142804 255960 142856 256012
rect 155408 255960 155460 256012
rect 255412 255960 255464 256012
rect 270776 255960 270828 256012
rect 270776 255484 270828 255536
rect 271788 255484 271840 255536
rect 49424 255280 49476 255332
rect 50804 255280 50856 255332
rect 100944 255280 100996 255332
rect 106096 255280 106148 255332
rect 133236 255280 133288 255332
rect 148324 255280 148376 255332
rect 191748 255280 191800 255332
rect 276020 254600 276072 254652
rect 298744 254600 298796 254652
rect 102784 254532 102836 254584
rect 123024 254532 123076 254584
rect 269028 254532 269080 254584
rect 583116 254532 583168 254584
rect 151084 253988 151136 254040
rect 191564 253988 191616 254040
rect 255412 253988 255464 254040
rect 267740 253988 267792 254040
rect 269028 253988 269080 254040
rect 49516 253920 49568 253972
rect 66812 253920 66864 253972
rect 106924 253920 106976 253972
rect 180248 253920 180300 253972
rect 255320 253920 255372 253972
rect 276020 253920 276072 253972
rect 15844 253852 15896 253904
rect 35256 253852 35308 253904
rect 35624 253852 35676 253904
rect 267004 253852 267056 253904
rect 268384 253852 268436 253904
rect 35256 253172 35308 253224
rect 66996 253172 67048 253224
rect 67364 253172 67416 253224
rect 129004 253172 129056 253224
rect 173256 253172 173308 253224
rect 271788 253172 271840 253224
rect 583392 253172 583444 253224
rect 188344 252628 188396 252680
rect 191012 252628 191064 252680
rect 255412 252628 255464 252680
rect 266452 252628 266504 252680
rect 267004 252628 267056 252680
rect 107752 252560 107804 252612
rect 111064 252560 111116 252612
rect 170496 252560 170548 252612
rect 191748 252560 191800 252612
rect 255504 252560 255556 252612
rect 270684 252560 270736 252612
rect 271788 252560 271840 252612
rect 100392 252492 100444 252544
rect 120816 252492 120868 252544
rect 109040 252424 109092 252476
rect 109684 252424 109736 252476
rect 263876 252288 263928 252340
rect 266912 252288 266964 252340
rect 163504 251880 163556 251932
rect 188252 251880 188304 251932
rect 38476 251812 38528 251864
rect 45928 251812 45980 251864
rect 135168 251812 135220 251864
rect 170404 251812 170456 251864
rect 255412 251540 255464 251592
rect 259736 251812 259788 251864
rect 582380 251812 582432 251864
rect 45928 251200 45980 251252
rect 46848 251200 46900 251252
rect 66812 251200 66864 251252
rect 109684 251200 109736 251252
rect 134616 251200 134668 251252
rect 135168 251200 135220 251252
rect 186964 251200 187016 251252
rect 191564 251200 191616 251252
rect 255504 251200 255556 251252
rect 262496 251200 262548 251252
rect 61568 250452 61620 250504
rect 66720 250452 66772 250504
rect 100852 250452 100904 250504
rect 107752 250452 107804 250504
rect 112444 250452 112496 250504
rect 114836 250452 114888 250504
rect 130568 250452 130620 250504
rect 133788 250452 133840 250504
rect 147772 250452 147824 250504
rect 192576 250452 192628 250504
rect 265164 250452 265216 250504
rect 582472 250452 582524 250504
rect 255320 249840 255372 249892
rect 265164 249840 265216 249892
rect 56508 249772 56560 249824
rect 100852 249772 100904 249824
rect 132592 249772 132644 249824
rect 133788 249772 133840 249824
rect 170404 249772 170456 249824
rect 191748 249772 191800 249824
rect 255412 249772 255464 249824
rect 266544 249772 266596 249824
rect 582380 249772 582432 249824
rect 61568 249704 61620 249756
rect 100944 249704 100996 249756
rect 111800 249704 111852 249756
rect 112352 249704 112404 249756
rect 112352 249092 112404 249144
rect 131304 249092 131356 249144
rect 100852 249024 100904 249076
rect 106648 249024 106700 249076
rect 122196 249024 122248 249076
rect 124312 249024 124364 249076
rect 187240 249024 187292 249076
rect 255320 248480 255372 248532
rect 268016 248480 268068 248532
rect 111616 248412 111668 248464
rect 114652 248412 114704 248464
rect 180156 248412 180208 248464
rect 190644 248412 190696 248464
rect 255688 248412 255740 248464
rect 271972 248412 272024 248464
rect 582564 248412 582616 248464
rect 100852 248344 100904 248396
rect 108948 248344 109000 248396
rect 42616 247664 42668 247716
rect 52460 247664 52512 247716
rect 108948 247664 109000 247716
rect 124220 247664 124272 247716
rect 254584 247664 254636 247716
rect 582472 247664 582524 247716
rect 62028 247052 62080 247104
rect 67456 247052 67508 247104
rect 188436 247052 188488 247104
rect 191748 247052 191800 247104
rect 255412 247052 255464 247104
rect 341524 247052 341576 247104
rect 100852 246916 100904 246968
rect 104348 246916 104400 246968
rect 100852 246304 100904 246356
rect 109040 246304 109092 246356
rect 120172 246304 120224 246356
rect 178684 246304 178736 246356
rect 59084 246100 59136 246152
rect 66996 246100 67048 246152
rect 67272 246100 67324 246152
rect 253204 245692 253256 245744
rect 313924 245692 313976 245744
rect 184296 245624 184348 245676
rect 191564 245624 191616 245676
rect 255412 245624 255464 245676
rect 258264 245624 258316 245676
rect 583300 245624 583352 245676
rect 100944 245556 100996 245608
rect 109684 245556 109736 245608
rect 254124 244944 254176 244996
rect 255596 244944 255648 244996
rect 55128 244876 55180 244928
rect 64604 244876 64656 244928
rect 66904 244876 66956 244928
rect 122104 244876 122156 244928
rect 142160 244876 142212 244928
rect 143448 244876 143500 244928
rect 255688 244332 255740 244384
rect 349804 244332 349856 244384
rect 100852 244264 100904 244316
rect 124312 244264 124364 244316
rect 143448 244264 143500 244316
rect 193036 244264 193088 244316
rect 260748 244264 260800 244316
rect 583392 244264 583444 244316
rect 103428 243584 103480 243636
rect 106280 243584 106332 243636
rect 105544 243516 105596 243568
rect 111800 243516 111852 243568
rect 163596 243516 163648 243568
rect 255504 243516 255556 243568
rect 262404 243516 262456 243568
rect 187056 242972 187108 243024
rect 191748 242972 191800 243024
rect 49608 242904 49660 242956
rect 55036 242904 55088 242956
rect 66812 242904 66864 242956
rect 98552 242904 98604 242956
rect 99288 242904 99340 242956
rect 103428 242904 103480 242956
rect 117964 242904 118016 242956
rect 193588 242904 193640 242956
rect 255412 242904 255464 242956
rect 261024 242972 261076 243024
rect 304264 242972 304316 243024
rect 262404 242904 262456 242956
rect 583116 242904 583168 242956
rect 253112 242836 253164 242888
rect 255688 242836 255740 242888
rect 100852 242700 100904 242752
rect 104256 242700 104308 242752
rect 54760 242156 54812 242208
rect 69020 242156 69072 242208
rect 118976 242156 119028 242208
rect 180340 242156 180392 242208
rect 255412 242156 255464 242208
rect 582748 242156 582800 242208
rect 251824 241884 251876 241936
rect 254124 241884 254176 241936
rect 250444 241816 250496 241868
rect 253112 241816 253164 241868
rect 69020 241748 69072 241800
rect 69848 241748 69900 241800
rect 94780 241748 94832 241800
rect 68560 241680 68612 241732
rect 69296 241680 69348 241732
rect 111064 241544 111116 241596
rect 193772 241544 193824 241596
rect 57612 241476 57664 241528
rect 77438 241476 77490 241528
rect 193680 241476 193732 241528
rect 213920 241476 213972 241528
rect 214748 241476 214800 241528
rect 255412 241476 255464 241528
rect 263784 241476 263836 241528
rect 291936 241476 291988 241528
rect 46664 241408 46716 241460
rect 71918 241408 71970 241460
rect 117228 241408 117280 241460
rect 255320 241408 255372 241460
rect 193036 241340 193088 241392
rect 199752 241340 199804 241392
rect 249248 241340 249300 241392
rect 253204 241340 253256 241392
rect 2780 241204 2832 241256
rect 4804 241204 4856 241256
rect 84660 240796 84712 240848
rect 112168 240796 112220 240848
rect 115940 240796 115992 240848
rect 117228 240796 117280 240848
rect 14464 240728 14516 240780
rect 88156 240728 88208 240780
rect 255320 240728 255372 240780
rect 580264 240728 580316 240780
rect 74540 240116 74592 240168
rect 74908 240116 74960 240168
rect 77300 240116 77352 240168
rect 78220 240116 78272 240168
rect 83096 240116 83148 240168
rect 83740 240116 83792 240168
rect 85580 240116 85632 240168
rect 85948 240116 86000 240168
rect 88340 240116 88392 240168
rect 88708 240116 88760 240168
rect 91100 240116 91152 240168
rect 92296 240116 92348 240168
rect 96620 240116 96672 240168
rect 96988 240116 97040 240168
rect 55956 240048 56008 240100
rect 56232 240048 56284 240100
rect 87052 240048 87104 240100
rect 93860 240048 93912 240100
rect 94228 240048 94280 240100
rect 103428 240048 103480 240100
rect 194784 240048 194836 240100
rect 250628 240048 250680 240100
rect 253020 240048 253072 240100
rect 64512 239980 64564 240032
rect 74632 239980 74684 240032
rect 83004 239980 83056 240032
rect 84016 239980 84068 240032
rect 128544 239980 128596 240032
rect 212264 239980 212316 240032
rect 80060 239436 80112 239488
rect 80428 239436 80480 239488
rect 252652 239436 252704 239488
rect 261116 239436 261168 239488
rect 11704 239368 11756 239420
rect 52368 239368 52420 239420
rect 55956 239368 56008 239420
rect 89628 239368 89680 239420
rect 106464 239368 106516 239420
rect 128544 239368 128596 239420
rect 243636 239368 243688 239420
rect 254584 239368 254636 239420
rect 38568 238688 38620 238740
rect 69112 238688 69164 238740
rect 69848 238688 69900 238740
rect 80152 238688 80204 238740
rect 83188 238688 83240 238740
rect 103520 238688 103572 238740
rect 192576 238688 192628 238740
rect 249156 238756 249208 238808
rect 258356 238756 258408 238808
rect 580356 238756 580408 238808
rect 53104 238620 53156 238672
rect 74540 238620 74592 238672
rect 88064 238620 88116 238672
rect 104992 238620 105044 238672
rect 180248 238620 180300 238672
rect 197268 238620 197320 238672
rect 87052 238076 87104 238128
rect 88064 238076 88116 238128
rect 104256 238008 104308 238060
rect 114744 238008 114796 238060
rect 119344 238008 119396 238060
rect 191288 238008 191340 238060
rect 232228 238008 232280 238060
rect 241520 238008 241572 238060
rect 243544 238008 243596 238060
rect 258172 238008 258224 238060
rect 69112 237396 69164 237448
rect 69664 237396 69716 237448
rect 80152 237396 80204 237448
rect 80704 237396 80756 237448
rect 82728 237396 82780 237448
rect 83188 237396 83240 237448
rect 39672 237328 39724 237380
rect 73252 237328 73304 237380
rect 88156 237328 88208 237380
rect 92572 237328 92624 237380
rect 102232 237328 102284 237380
rect 252836 237328 252888 237380
rect 111892 237260 111944 237312
rect 187240 237260 187292 237312
rect 224776 237260 224828 237312
rect 74724 236716 74776 236768
rect 89168 236716 89220 236768
rect 60464 236648 60516 236700
rect 76104 236648 76156 236700
rect 93124 236648 93176 236700
rect 102232 236648 102284 236700
rect 253204 236648 253256 236700
rect 263692 236648 263744 236700
rect 90824 235968 90876 236020
rect 91100 235968 91152 236020
rect 67364 235900 67416 235952
rect 111064 235900 111116 235952
rect 180340 235900 180392 235952
rect 202236 235900 202288 235952
rect 202788 235900 202840 235952
rect 50988 235832 51040 235884
rect 77300 235832 77352 235884
rect 94044 235492 94096 235544
rect 94504 235492 94556 235544
rect 102324 235492 102376 235544
rect 84108 235220 84160 235272
rect 89720 235220 89772 235272
rect 102784 235220 102836 235272
rect 107016 235220 107068 235272
rect 134708 235220 134760 235272
rect 142896 235220 142948 235272
rect 202788 235220 202840 235272
rect 246304 235220 246356 235272
rect 217324 234608 217376 234660
rect 267004 234608 267056 234660
rect 80060 234540 80112 234592
rect 111800 234540 111852 234592
rect 117688 234540 117740 234592
rect 117964 234540 118016 234592
rect 122196 234540 122248 234592
rect 182916 234540 182968 234592
rect 254032 234540 254084 234592
rect 193680 234472 193732 234524
rect 219716 234472 219768 234524
rect 68284 233928 68336 233980
rect 80428 233928 80480 233980
rect 4804 233860 4856 233912
rect 97816 233860 97868 233912
rect 114468 233860 114520 233912
rect 115940 233860 115992 233912
rect 122104 233860 122156 233912
rect 191104 233860 191156 233912
rect 100668 233248 100720 233300
rect 100852 233248 100904 233300
rect 103520 233248 103572 233300
rect 114652 233248 114704 233300
rect 138664 233248 138716 233300
rect 236644 233248 236696 233300
rect 237196 233248 237248 233300
rect 298100 233248 298152 233300
rect 76656 233180 76708 233232
rect 78680 233180 78732 233232
rect 80980 233180 81032 233232
rect 72792 233112 72844 233164
rect 75920 233112 75972 233164
rect 106924 233180 106976 233232
rect 193772 233180 193824 233232
rect 259552 233180 259604 233232
rect 74816 233044 74868 233096
rect 80980 232976 81032 233028
rect 109316 233112 109368 233164
rect 43812 232500 43864 232552
rect 71964 232500 72016 232552
rect 72792 232500 72844 232552
rect 199752 232500 199804 232552
rect 250444 232500 250496 232552
rect 255964 231820 256016 231872
rect 582564 231820 582616 231872
rect 174544 231752 174596 231804
rect 256792 231752 256844 231804
rect 207204 231684 207256 231736
rect 207664 231684 207716 231736
rect 39948 231072 40000 231124
rect 189816 231072 189868 231124
rect 207664 230460 207716 230512
rect 270592 230460 270644 230512
rect 133236 230392 133288 230444
rect 263876 230392 263928 230444
rect 80336 229780 80388 229832
rect 92388 229780 92440 229832
rect 114836 229780 114888 229832
rect 12348 229712 12400 229764
rect 191840 229712 191892 229764
rect 193220 229712 193272 229764
rect 251272 229712 251324 229764
rect 122748 229100 122800 229152
rect 123116 229100 123168 229152
rect 119436 228556 119488 228608
rect 120264 228556 120316 228608
rect 57704 228352 57756 228404
rect 70400 228352 70452 228404
rect 120264 228284 120316 228336
rect 252928 228352 252980 228404
rect 255504 228352 255556 228404
rect 583208 228352 583260 228404
rect 81440 227944 81492 227996
rect 85580 227944 85632 227996
rect 92204 227808 92256 227860
rect 88340 227740 88392 227792
rect 93124 227740 93176 227792
rect 94504 227740 94556 227792
rect 95976 227740 96028 227792
rect 100760 227740 100812 227792
rect 209780 227740 209832 227792
rect 256056 227740 256108 227792
rect 95148 227672 95200 227724
rect 129004 227672 129056 227724
rect 181536 227672 181588 227724
rect 244740 227672 244792 227724
rect 82084 227604 82136 227656
rect 103520 227604 103572 227656
rect 108304 226992 108356 227044
rect 191196 226992 191248 227044
rect 234620 226992 234672 227044
rect 291844 226992 291896 227044
rect 291936 226992 291988 227044
rect 582380 226992 582432 227044
rect 68928 226312 68980 226364
rect 71780 226312 71832 226364
rect 128544 226312 128596 226364
rect 129004 226312 129056 226364
rect 52184 226244 52236 226296
rect 77392 226244 77444 226296
rect 78588 226244 78640 226296
rect 125692 226244 125744 226296
rect 265072 226244 265124 226296
rect 88248 225632 88300 225684
rect 102140 225632 102192 225684
rect 101496 225564 101548 225616
rect 111984 225564 112036 225616
rect 125692 225564 125744 225616
rect 251916 224952 251968 225004
rect 351920 224952 351972 225004
rect 88432 224884 88484 224936
rect 115940 224884 115992 224936
rect 136548 224884 136600 224936
rect 255964 224884 256016 224936
rect 52276 224204 52328 224256
rect 76748 224204 76800 224256
rect 131764 224204 131816 224256
rect 135444 224204 135496 224256
rect 136548 224204 136600 224256
rect 89720 224136 89772 224188
rect 94780 224136 94832 224188
rect 229744 223592 229796 223644
rect 288440 223592 288492 223644
rect 130476 223524 130528 223576
rect 131028 223524 131080 223576
rect 222200 223524 222252 223576
rect 184388 223456 184440 223508
rect 265164 223456 265216 223508
rect 86868 222844 86920 222896
rect 112076 222844 112128 222896
rect 242256 222164 242308 222216
rect 306380 222164 306432 222216
rect 50344 222096 50396 222148
rect 50896 222096 50948 222148
rect 266544 222096 266596 222148
rect 126244 221416 126296 221468
rect 234712 221416 234764 221468
rect 244740 221416 244792 221468
rect 309784 221416 309836 221468
rect 98644 220804 98696 220856
rect 126888 220804 126940 220856
rect 69664 220736 69716 220788
rect 209780 220736 209832 220788
rect 247224 220736 247276 220788
rect 247684 220736 247736 220788
rect 58992 220056 59044 220108
rect 71780 220056 71832 220108
rect 247684 219444 247736 219496
rect 331220 219444 331272 219496
rect 41144 219376 41196 219428
rect 243636 219376 243688 219428
rect 268384 219376 268436 219428
rect 580172 219376 580224 219428
rect 107568 218696 107620 218748
rect 177396 218696 177448 218748
rect 213920 218696 213972 218748
rect 267924 218696 267976 218748
rect 53472 217948 53524 218000
rect 273444 217948 273496 218000
rect 104164 217404 104216 217456
rect 110420 217404 110472 217456
rect 125508 217268 125560 217320
rect 171784 217268 171836 217320
rect 280896 217268 280948 217320
rect 303620 217268 303672 217320
rect 73804 216588 73856 216640
rect 74448 216588 74500 216640
rect 267740 216588 267792 216640
rect 110604 216520 110656 216572
rect 242164 216520 242216 216572
rect 75920 215908 75972 215960
rect 110604 215908 110656 215960
rect 249156 215908 249208 215960
rect 338120 215908 338172 215960
rect 115756 215228 115808 215280
rect 261024 215228 261076 215280
rect 117228 215160 117280 215212
rect 241520 215160 241572 215212
rect 242164 215160 242216 215212
rect 88984 214616 89036 214668
rect 114560 214616 114612 214668
rect 115756 214616 115808 214668
rect 84844 214548 84896 214600
rect 116032 214548 116084 214600
rect 117228 214548 117280 214600
rect 3148 213936 3200 213988
rect 8208 213868 8260 213920
rect 36544 213868 36596 213920
rect 66812 213800 66864 213852
rect 67272 213800 67324 213852
rect 243544 213868 243596 213920
rect 139400 213800 139452 213852
rect 200764 213800 200816 213852
rect 100668 213188 100720 213240
rect 127256 213188 127308 213240
rect 139400 213188 139452 213240
rect 55128 212440 55180 212492
rect 247684 212440 247736 212492
rect 128636 212372 128688 212424
rect 250628 212372 250680 212424
rect 48044 211760 48096 211812
rect 76656 211760 76708 211812
rect 88064 211760 88116 211812
rect 116768 211760 116820 211812
rect 68468 211080 68520 211132
rect 68928 211080 68980 211132
rect 253940 211080 253992 211132
rect 54944 211012 54996 211064
rect 217324 211012 217376 211064
rect 92204 209108 92256 209160
rect 118700 209108 118752 209160
rect 271880 209108 271932 209160
rect 80704 209040 80756 209092
rect 103612 209040 103664 209092
rect 266452 209040 266504 209092
rect 61660 208292 61712 208344
rect 236644 208292 236696 208344
rect 136640 208224 136692 208276
rect 265256 208224 265308 208276
rect 96620 207612 96672 207664
rect 128360 207612 128412 207664
rect 136640 207612 136692 207664
rect 56416 206932 56468 206984
rect 207664 206932 207716 206984
rect 99196 206252 99248 206304
rect 240140 206184 240192 206236
rect 240784 206184 240836 206236
rect 98736 205640 98788 205692
rect 99196 205640 99248 205692
rect 61936 205572 61988 205624
rect 229744 205572 229796 205624
rect 126980 205504 127032 205556
rect 263600 205504 263652 205556
rect 91008 204892 91060 204944
rect 106280 204892 106332 204944
rect 126980 204892 127032 204944
rect 102968 204212 103020 204264
rect 103428 204212 103480 204264
rect 262404 204212 262456 204264
rect 82912 203532 82964 203584
rect 105084 203532 105136 203584
rect 138664 202784 138716 202836
rect 263784 202784 263836 202836
rect 3240 202104 3292 202156
rect 124220 202104 124272 202156
rect 105636 202036 105688 202088
rect 112168 202036 112220 202088
rect 129004 201492 129056 201544
rect 132592 201492 132644 201544
rect 122196 201424 122248 201476
rect 122748 201424 122800 201476
rect 271972 201424 272024 201476
rect 147036 200744 147088 200796
rect 163504 200744 163556 200796
rect 82728 199520 82780 199572
rect 90364 199520 90416 199572
rect 89812 199452 89864 199504
rect 102968 199452 103020 199504
rect 56324 199384 56376 199436
rect 80060 199384 80112 199436
rect 88156 199384 88208 199436
rect 102140 199384 102192 199436
rect 50988 198636 51040 198688
rect 249064 198636 249116 198688
rect 88156 197956 88208 198008
rect 115388 197956 115440 198008
rect 46756 197276 46808 197328
rect 276020 197276 276072 197328
rect 46204 196936 46256 196988
rect 46756 196936 46808 196988
rect 59176 196596 59228 196648
rect 77484 196596 77536 196648
rect 88064 196596 88116 196648
rect 107844 196596 107896 196648
rect 116768 195916 116820 195968
rect 269212 195916 269264 195968
rect 55036 194488 55088 194540
rect 267832 194488 267884 194540
rect 37096 193808 37148 193860
rect 68284 193808 68336 193860
rect 86776 193808 86828 193860
rect 114652 193808 114704 193860
rect 313924 193128 313976 193180
rect 580172 193128 580224 193180
rect 85580 191156 85632 191208
rect 142160 191156 142212 191208
rect 1308 191088 1360 191140
rect 157984 191088 158036 191140
rect 118608 189728 118660 189780
rect 181444 189728 181496 189780
rect 2780 188844 2832 188896
rect 4804 188844 4856 188896
rect 204904 185580 204956 185632
rect 259552 185580 259604 185632
rect 37188 184152 37240 184204
rect 151176 184152 151228 184204
rect 289084 184152 289136 184204
rect 300860 184152 300912 184204
rect 2688 182792 2740 182844
rect 166356 182792 166408 182844
rect 81532 180820 81584 180872
rect 84844 180820 84896 180872
rect 5356 180072 5408 180124
rect 156604 180072 156656 180124
rect 341524 179324 341576 179376
rect 580172 179324 580224 179376
rect 28908 167628 28960 167680
rect 184296 167628 184348 167680
rect 114468 164840 114520 164892
rect 178776 164840 178828 164892
rect 20628 162120 20680 162172
rect 187056 162120 187108 162172
rect 58992 160692 59044 160744
rect 73804 160692 73856 160744
rect 66076 159332 66128 159384
rect 273260 159332 273312 159384
rect 37096 157972 37148 158024
rect 188436 157972 188488 158024
rect 84108 156680 84160 156732
rect 102232 156680 102284 156732
rect 89076 156612 89128 156664
rect 116584 156612 116636 156664
rect 316040 156612 316092 156664
rect 61752 155252 61804 155304
rect 75184 155252 75236 155304
rect 43996 155184 44048 155236
rect 180156 155184 180208 155236
rect 2964 149064 3016 149116
rect 14464 149064 14516 149116
rect 63132 148996 63184 149048
rect 276664 148996 276716 149048
rect 313280 149064 313332 149116
rect 39764 148316 39816 148368
rect 73344 148316 73396 148368
rect 84568 147636 84620 147688
rect 89076 147636 89128 147688
rect 76012 146072 76064 146124
rect 79324 146072 79376 146124
rect 50804 145528 50856 145580
rect 70492 145528 70544 145580
rect 84108 145528 84160 145580
rect 116676 145528 116728 145580
rect 41236 144236 41288 144288
rect 74816 144236 74868 144288
rect 53564 144168 53616 144220
rect 170496 144168 170548 144220
rect 54852 142808 54904 142860
rect 74540 142808 74592 142860
rect 85488 142808 85540 142860
rect 94780 142808 94832 142860
rect 82820 142128 82872 142180
rect 86224 142128 86276 142180
rect 88248 142128 88300 142180
rect 100852 142128 100904 142180
rect 81348 141448 81400 141500
rect 106372 141448 106424 141500
rect 3424 141380 3476 141432
rect 88156 141380 88208 141432
rect 71688 140768 71740 140820
rect 76564 140768 76616 140820
rect 106924 140768 106976 140820
rect 114744 140768 114796 140820
rect 88156 140700 88208 140752
rect 110512 140700 110564 140752
rect 56324 140088 56376 140140
rect 78772 140088 78824 140140
rect 45376 140020 45428 140072
rect 72332 140020 72384 140072
rect 91008 140020 91060 140072
rect 102784 140020 102836 140072
rect 85488 139408 85540 139460
rect 88984 139408 89036 139460
rect 14464 139340 14516 139392
rect 88248 139340 88300 139392
rect 349804 139340 349856 139392
rect 580172 139340 580224 139392
rect 94596 138728 94648 138780
rect 113364 138728 113416 138780
rect 60372 138660 60424 138712
rect 74632 138660 74684 138712
rect 79324 138660 79376 138712
rect 111616 138660 111668 138712
rect 198004 138660 198056 138712
rect 75920 138048 75972 138100
rect 76380 138048 76432 138100
rect 81440 138048 81492 138100
rect 82084 138048 82136 138100
rect 89720 138048 89772 138100
rect 90180 138048 90232 138100
rect 3240 137912 3292 137964
rect 39856 137912 39908 137964
rect 78496 137368 78548 137420
rect 80428 137368 80480 137420
rect 88064 137300 88116 137352
rect 102784 137300 102836 137352
rect 39856 137232 39908 137284
rect 73160 137232 73212 137284
rect 79048 137232 79100 137284
rect 86868 137232 86920 137284
rect 89076 137232 89128 137284
rect 124864 137232 124916 137284
rect 170496 137232 170548 137284
rect 68284 136620 68336 136672
rect 69940 136620 69992 136672
rect 74724 136620 74776 136672
rect 76104 136620 76156 136672
rect 83648 136620 83700 136672
rect 84108 136620 84160 136672
rect 85948 136620 86000 136672
rect 88064 136620 88116 136672
rect 14464 135872 14516 135924
rect 91008 135872 91060 135924
rect 91284 135872 91336 135924
rect 91192 135804 91244 135856
rect 109132 135872 109184 135924
rect 44824 135260 44876 135312
rect 91192 135260 91244 135312
rect 92296 135260 92348 135312
rect 276020 135260 276072 135312
rect 35716 135192 35768 135244
rect 66260 135192 66312 135244
rect 94780 135192 94832 135244
rect 99380 135192 99432 135244
rect 40868 135124 40920 135176
rect 41328 135124 41380 135176
rect 75460 135124 75512 135176
rect 68652 134784 68704 134836
rect 69664 134784 69716 134836
rect 89260 134784 89312 134836
rect 90364 134784 90416 134836
rect 96068 134784 96120 134836
rect 94872 134716 94924 134768
rect 70492 134580 70544 134632
rect 71228 134580 71280 134632
rect 3424 134512 3476 134564
rect 40868 134512 40920 134564
rect 47860 133832 47912 133884
rect 66260 133832 66312 133884
rect 96712 133832 96764 133884
rect 122196 133832 122248 133884
rect 94964 133152 95016 133204
rect 267832 133152 267884 133204
rect 44088 132404 44140 132456
rect 66260 132404 66312 132456
rect 96620 132404 96672 132456
rect 131764 132404 131816 132456
rect 53656 132336 53708 132388
rect 66352 132336 66404 132388
rect 96712 129684 96764 129736
rect 131212 129684 131264 129736
rect 97264 129616 97316 129668
rect 127164 129616 127216 129668
rect 57888 129004 57940 129056
rect 66444 129004 66496 129056
rect 32864 128256 32916 128308
rect 66904 128256 66956 128308
rect 97540 128256 97592 128308
rect 134708 128256 134760 128308
rect 59084 128188 59136 128240
rect 66720 128188 66772 128240
rect 97172 128188 97224 128240
rect 100852 128188 100904 128240
rect 97816 126896 97868 126948
rect 135260 126896 135312 126948
rect 43904 126216 43956 126268
rect 66904 126216 66956 126268
rect 101496 126216 101548 126268
rect 106464 126216 106516 126268
rect 57796 125536 57848 125588
rect 66260 125536 66312 125588
rect 97448 125536 97500 125588
rect 122840 125536 122892 125588
rect 96804 124856 96856 124908
rect 128452 124856 128504 124908
rect 59268 124108 59320 124160
rect 63224 124108 63276 124160
rect 94688 124108 94740 124160
rect 95148 124108 95200 124160
rect 97816 124108 97868 124160
rect 130384 124108 130436 124160
rect 130568 124108 130620 124160
rect 96620 123972 96672 124024
rect 98736 123972 98788 124024
rect 130568 123428 130620 123480
rect 173256 123428 173308 123480
rect 63224 122884 63276 122936
rect 66904 122884 66956 122936
rect 53380 122748 53432 122800
rect 66904 122748 66956 122800
rect 97816 122748 97868 122800
rect 135904 122748 135956 122800
rect 61660 122680 61712 122732
rect 66720 122680 66772 122732
rect 96068 122272 96120 122324
rect 98000 122272 98052 122324
rect 135904 122068 135956 122120
rect 356060 122068 356112 122120
rect 32956 121388 33008 121440
rect 65524 121388 65576 121440
rect 97816 121388 97868 121440
rect 113272 121388 113324 121440
rect 60556 120164 60608 120216
rect 66260 120164 66312 120216
rect 97816 120164 97868 120216
rect 104900 120164 104952 120216
rect 54944 120028 54996 120080
rect 66904 120028 66956 120080
rect 123576 119348 123628 119400
rect 159456 119348 159508 119400
rect 97816 118600 97868 118652
rect 122932 118600 122984 118652
rect 41144 118532 41196 118584
rect 66904 118532 66956 118584
rect 50896 117240 50948 117292
rect 66904 117240 66956 117292
rect 97816 117240 97868 117292
rect 120080 117240 120132 117292
rect 96620 117036 96672 117088
rect 98644 117036 98696 117088
rect 100024 116288 100076 116340
rect 104992 116288 105044 116340
rect 47952 115880 48004 115932
rect 66904 115880 66956 115932
rect 97724 115880 97776 115932
rect 133144 115880 133196 115932
rect 133788 115880 133840 115932
rect 97816 115812 97868 115864
rect 118792 115812 118844 115864
rect 133788 115200 133840 115252
rect 187056 115200 187108 115252
rect 60648 114588 60700 114640
rect 67180 114588 67232 114640
rect 8208 114452 8260 114504
rect 66628 114452 66680 114504
rect 63500 114384 63552 114436
rect 64604 114384 64656 114436
rect 96620 113840 96672 113892
rect 109224 113840 109276 113892
rect 102784 113772 102836 113824
rect 255320 113772 255372 113824
rect 34336 113092 34388 113144
rect 66904 113092 66956 113144
rect 97816 113092 97868 113144
rect 129740 113092 129792 113144
rect 102140 112412 102192 112464
rect 125692 112412 125744 112464
rect 169116 112412 169168 112464
rect 264244 112412 264296 112464
rect 3148 111732 3200 111784
rect 44824 111732 44876 111784
rect 56416 111732 56468 111784
rect 66904 111732 66956 111784
rect 97908 111732 97960 111784
rect 136732 111732 136784 111784
rect 101404 110984 101456 111036
rect 104900 110984 104952 111036
rect 46756 110372 46808 110424
rect 66904 110372 66956 110424
rect 97816 110372 97868 110424
rect 133236 110372 133288 110424
rect 97908 110304 97960 110356
rect 127072 110304 127124 110356
rect 45468 109692 45520 109744
rect 57060 109692 57112 109744
rect 127072 109692 127124 109744
rect 273904 109692 273956 109744
rect 56600 109012 56652 109064
rect 57060 109012 57112 109064
rect 66260 109012 66312 109064
rect 52184 108944 52236 108996
rect 66996 108944 67048 108996
rect 97908 108944 97960 108996
rect 113180 108944 113232 108996
rect 57612 108876 57664 108928
rect 66904 108876 66956 108928
rect 97724 108876 97776 108928
rect 111984 108876 112036 108928
rect 41420 107584 41472 107636
rect 42708 107584 42760 107636
rect 66904 107584 66956 107636
rect 49608 107516 49660 107568
rect 66720 107516 66772 107568
rect 97540 107312 97592 107364
rect 102140 107312 102192 107364
rect 7564 106904 7616 106956
rect 41420 106904 41472 106956
rect 103428 106904 103480 106956
rect 182824 106904 182876 106956
rect 49516 106224 49568 106276
rect 66904 106224 66956 106276
rect 97632 106224 97684 106276
rect 125784 106224 125836 106276
rect 97908 105544 97960 105596
rect 180156 105544 180208 105596
rect 60464 104796 60516 104848
rect 66260 104796 66312 104848
rect 97172 104796 97224 104848
rect 107752 104796 107804 104848
rect 94780 104728 94832 104780
rect 102324 104728 102376 104780
rect 61936 103436 61988 103488
rect 66904 103436 66956 103488
rect 97172 103436 97224 103488
rect 135352 103436 135404 103488
rect 97724 102756 97776 102808
rect 120172 102756 120224 102808
rect 135352 102756 135404 102808
rect 184296 102756 184348 102808
rect 64696 102076 64748 102128
rect 66444 102076 66496 102128
rect 97908 102076 97960 102128
rect 131304 102076 131356 102128
rect 97816 102008 97868 102060
rect 124220 102008 124272 102060
rect 46848 101396 46900 101448
rect 60740 101396 60792 101448
rect 66812 101396 66864 101448
rect 131304 101396 131356 101448
rect 233148 101396 233200 101448
rect 61568 100648 61620 100700
rect 66812 100648 66864 100700
rect 97908 100648 97960 100700
rect 130200 100648 130252 100700
rect 130200 99968 130252 100020
rect 131028 99968 131080 100020
rect 151176 99968 151228 100020
rect 168288 99968 168340 100020
rect 198096 99968 198148 100020
rect 56508 99492 56560 99544
rect 63408 99492 63460 99544
rect 66812 99492 66864 99544
rect 53472 99288 53524 99340
rect 66812 99288 66864 99340
rect 97540 99288 97592 99340
rect 134616 99288 134668 99340
rect 135168 99288 135220 99340
rect 135168 98608 135220 98660
rect 220084 98608 220136 98660
rect 97908 97928 97960 97980
rect 111892 97928 111944 97980
rect 97540 97860 97592 97912
rect 106924 97860 106976 97912
rect 55128 97248 55180 97300
rect 66812 97248 66864 97300
rect 3056 96636 3108 96688
rect 65616 96636 65668 96688
rect 42616 96568 42668 96620
rect 66260 96568 66312 96620
rect 97908 95956 97960 96008
rect 99288 95956 99340 96008
rect 178776 95956 178828 96008
rect 175188 95888 175240 95940
rect 276112 95888 276164 95940
rect 55036 95140 55088 95192
rect 66444 95140 66496 95192
rect 97908 95140 97960 95192
rect 110420 95140 110472 95192
rect 64788 93780 64840 93832
rect 66812 93780 66864 93832
rect 97908 93780 97960 93832
rect 128360 93780 128412 93832
rect 94688 93508 94740 93560
rect 95884 93508 95936 93560
rect 95056 93100 95108 93152
rect 103520 93100 103572 93152
rect 67640 92828 67692 92880
rect 68652 92828 68704 92880
rect 54852 92760 54904 92812
rect 72838 92692 72890 92744
rect 91790 92692 91842 92744
rect 94780 92692 94832 92744
rect 68468 92624 68520 92676
rect 71734 92624 71786 92676
rect 52368 92420 52420 92472
rect 86040 92420 86092 92472
rect 89260 92420 89312 92472
rect 106280 92420 106332 92472
rect 63316 92352 63368 92404
rect 73344 92352 73396 92404
rect 86684 92352 86736 92404
rect 98736 92352 98788 92404
rect 90180 90992 90232 91044
rect 95240 90992 95292 91044
rect 96160 90992 96212 91044
rect 88248 90856 88300 90908
rect 117964 90856 118016 90908
rect 74356 90720 74408 90772
rect 75276 90720 75328 90772
rect 87604 90516 87656 90568
rect 88248 90516 88300 90568
rect 82636 89904 82688 89956
rect 86868 89904 86920 89956
rect 80980 89700 81032 89752
rect 83464 89700 83516 89752
rect 85212 89700 85264 89752
rect 89536 89700 89588 89752
rect 48044 89632 48096 89684
rect 78312 89632 78364 89684
rect 92388 89632 92440 89684
rect 118700 89632 118752 89684
rect 52276 89564 52328 89616
rect 76288 89564 76340 89616
rect 84108 89564 84160 89616
rect 100024 89564 100076 89616
rect 119988 88952 120040 89004
rect 137284 88952 137336 89004
rect 59176 88272 59228 88324
rect 76564 88272 76616 88324
rect 76840 88272 76892 88324
rect 80060 88272 80112 88324
rect 111800 88272 111852 88324
rect 60372 88204 60424 88256
rect 73804 88204 73856 88256
rect 87236 88204 87288 88256
rect 115940 88204 115992 88256
rect 111800 87592 111852 87644
rect 188436 87592 188488 87644
rect 65616 86912 65668 86964
rect 96712 86912 96764 86964
rect 61752 86844 61804 86896
rect 75184 86844 75236 86896
rect 75368 86844 75420 86896
rect 88156 86844 88208 86896
rect 101496 86844 101548 86896
rect 3516 85484 3568 85536
rect 56600 85484 56652 85536
rect 86868 85484 86920 85536
rect 98000 85484 98052 85536
rect 66076 84804 66128 84856
rect 338212 84804 338264 84856
rect 56324 84124 56376 84176
rect 78680 84124 78732 84176
rect 92480 84124 92532 84176
rect 93768 84124 93820 84176
rect 128544 84124 128596 84176
rect 85580 84056 85632 84108
rect 86776 84056 86828 84108
rect 99380 84056 99432 84108
rect 78680 82832 78732 82884
rect 79324 82832 79376 82884
rect 83464 82764 83516 82816
rect 84108 82764 84160 82816
rect 107660 82764 107712 82816
rect 63224 82084 63276 82136
rect 327172 82084 327224 82136
rect 62028 80724 62080 80776
rect 151084 80724 151136 80776
rect 96160 80656 96212 80708
rect 349160 80656 349212 80708
rect 67180 79296 67232 79348
rect 280160 79296 280212 79348
rect 75276 78616 75328 78668
rect 100760 78616 100812 78668
rect 101128 78616 101180 78668
rect 48136 78004 48188 78056
rect 123576 78004 123628 78056
rect 101128 77936 101180 77988
rect 340880 77936 340932 77988
rect 63408 77188 63460 77240
rect 252560 77188 252612 77240
rect 253204 77188 253256 77240
rect 79968 75148 80020 75200
rect 184204 75148 184256 75200
rect 108948 73788 109000 73840
rect 146944 73788 146996 73840
rect 3516 71680 3568 71732
rect 101404 71680 101456 71732
rect 96528 71000 96580 71052
rect 155316 71000 155368 71052
rect 79324 69640 79376 69692
rect 343640 69640 343692 69692
rect 66076 68348 66128 68400
rect 162124 68348 162176 68400
rect 70308 68280 70360 68332
rect 180064 68280 180116 68332
rect 65524 66852 65576 66904
rect 332600 66852 332652 66904
rect 10968 65492 11020 65544
rect 178684 65492 178736 65544
rect 68928 64132 68980 64184
rect 189724 64132 189776 64184
rect 70216 62772 70268 62824
rect 311900 62772 311952 62824
rect 95056 61412 95108 61464
rect 141516 61412 141568 61464
rect 72424 61344 72476 61396
rect 97264 61344 97316 61396
rect 129004 61344 129056 61396
rect 206376 61344 206428 61396
rect 304264 60664 304316 60716
rect 580172 60664 580224 60716
rect 67640 59984 67692 60036
rect 291200 59984 291252 60036
rect 86776 58624 86828 58676
rect 253204 58624 253256 58676
rect 71688 57264 71740 57316
rect 173164 57264 173216 57316
rect 165528 57196 165580 57248
rect 304264 57196 304316 57248
rect 67548 56516 67600 56568
rect 269120 56516 269172 56568
rect 88156 54476 88208 54528
rect 266360 54476 266412 54528
rect 75184 53048 75236 53100
rect 224224 53048 224276 53100
rect 75828 51688 75880 51740
rect 177304 51688 177356 51740
rect 193128 51688 193180 51740
rect 242992 51688 243044 51740
rect 59268 50396 59320 50448
rect 166264 50396 166316 50448
rect 89536 50328 89588 50380
rect 289084 50328 289136 50380
rect 73804 48968 73856 49020
rect 231124 48968 231176 49020
rect 248420 48492 248472 48544
rect 252560 48492 252612 48544
rect 76564 46180 76616 46232
rect 322204 46180 322256 46232
rect 3424 45500 3476 45552
rect 60740 45500 60792 45552
rect 93768 44820 93820 44872
rect 302332 44820 302384 44872
rect 84108 43392 84160 43444
rect 274640 43392 274692 43444
rect 249064 42304 249116 42356
rect 249800 42304 249852 42356
rect 88248 42032 88300 42084
rect 284392 42032 284444 42084
rect 64604 40672 64656 40724
rect 307852 40672 307904 40724
rect 198004 39312 198056 39364
rect 262864 39312 262916 39364
rect 3976 37884 4028 37936
rect 160836 37884 160888 37936
rect 3516 33056 3568 33108
rect 14464 33056 14516 33108
rect 82728 32376 82780 32428
rect 147036 32376 147088 32428
rect 88984 26868 89036 26920
rect 213184 26868 213236 26920
rect 280804 22720 280856 22772
rect 292672 22720 292724 22772
rect 295984 22720 296036 22772
rect 335360 22720 335412 22772
rect 151176 21360 151228 21412
rect 277492 21360 277544 21412
rect 3424 20612 3476 20664
rect 72424 20612 72476 20664
rect 78588 20000 78640 20052
rect 175924 20000 175976 20052
rect 170496 19932 170548 19984
rect 325700 19932 325752 19984
rect 88248 18640 88300 18692
rect 206284 18640 206336 18692
rect 50988 18572 51040 18624
rect 186964 18572 187016 18624
rect 220084 18572 220136 18624
rect 331312 18572 331364 18624
rect 97908 17280 97960 17332
rect 142804 17280 142856 17332
rect 65984 17212 66036 17264
rect 125600 17212 125652 17264
rect 253204 17212 253256 17264
rect 287152 17212 287204 17264
rect 307852 16192 307904 16244
rect 309048 16192 309100 16244
rect 64788 15920 64840 15972
rect 148324 15920 148376 15972
rect 86868 15852 86920 15904
rect 322940 15852 322992 15904
rect 46664 14424 46716 14476
rect 170404 14424 170456 14476
rect 173256 14424 173308 14476
rect 337016 14424 337068 14476
rect 89536 13132 89588 13184
rect 185584 13132 185636 13184
rect 45376 13064 45428 13116
rect 160744 13064 160796 13116
rect 273904 13064 273956 13116
rect 324872 13064 324924 13116
rect 3424 12384 3476 12436
rect 7564 12384 7616 12436
rect 178776 11704 178828 11756
rect 241704 11704 241756 11756
rect 262864 11704 262916 11756
rect 302884 11704 302936 11756
rect 89628 10956 89680 11008
rect 333980 10956 334032 11008
rect 334624 10956 334676 11008
rect 112 10276 164 10328
rect 96620 10276 96672 10328
rect 61936 8916 61988 8968
rect 169024 8916 169076 8968
rect 180156 8916 180208 8968
rect 346952 8916 347004 8968
rect 54944 7556 54996 7608
rect 129004 7556 129056 7608
rect 184296 7556 184348 7608
rect 317328 7556 317380 7608
rect 92480 6196 92532 6248
rect 155224 6196 155276 6248
rect 83280 6128 83332 6180
rect 159364 6128 159416 6180
rect 198096 6128 198148 6180
rect 247592 6128 247644 6180
rect 261760 6128 261812 6180
rect 270500 6128 270552 6180
rect 305644 6128 305696 6180
rect 311440 6128 311492 6180
rect 310244 5516 310296 5568
rect 313280 5516 313332 5568
rect 187056 4768 187108 4820
rect 257068 4768 257120 4820
rect 264244 4768 264296 4820
rect 279516 4768 279568 4820
rect 281908 4768 281960 4820
rect 287060 4768 287112 4820
rect 122288 4088 122340 4140
rect 123484 4088 123536 4140
rect 304264 3952 304316 4004
rect 307944 3952 307996 4004
rect 342168 3680 342220 3732
rect 345020 3680 345072 3732
rect 30104 3612 30156 3664
rect 40684 3612 40736 3664
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 5448 3476 5500 3528
rect 13544 3544 13596 3596
rect 52552 3544 52604 3596
rect 53656 3544 53708 3596
rect 60832 3544 60884 3596
rect 62028 3544 62080 3596
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12348 3476 12400 3528
rect 15936 3476 15988 3528
rect 16396 3476 16448 3528
rect 19432 3476 19484 3528
rect 20536 3476 20588 3528
rect 20628 3476 20680 3528
rect 21364 3476 21416 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 35992 3476 36044 3528
rect 37096 3476 37148 3528
rect 40684 3476 40736 3528
rect 41328 3476 41380 3528
rect 41880 3476 41932 3528
rect 42708 3476 42760 3528
rect 43076 3476 43128 3528
rect 43996 3476 44048 3528
rect 44272 3476 44324 3528
rect 45376 3476 45428 3528
rect 48228 3476 48280 3528
rect 48964 3476 49016 3528
rect 50160 3476 50212 3528
rect 50988 3476 51040 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 72516 3544 72568 3596
rect 92756 3544 92808 3596
rect 108304 3612 108356 3664
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 69112 3476 69164 3528
rect 70216 3476 70268 3528
rect 73804 3476 73856 3528
rect 74448 3476 74500 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 82084 3476 82136 3528
rect 82728 3476 82780 3528
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 86868 3476 86920 3528
rect 87604 3476 87656 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 92388 3476 92440 3528
rect 97448 3476 97500 3528
rect 97908 3476 97960 3528
rect 99840 3476 99892 3528
rect 119344 3544 119396 3596
rect 123484 3544 123536 3596
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 121092 3476 121144 3528
rect 122104 3476 122156 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 276020 3544 276072 3596
rect 277124 3544 277176 3596
rect 134524 3476 134576 3528
rect 143540 3476 143592 3528
rect 144828 3476 144880 3528
rect 224224 3476 224276 3528
rect 246396 3476 246448 3528
rect 264152 3476 264204 3528
rect 270592 3476 270644 3528
rect 282184 3476 282236 3528
rect 283104 3476 283156 3528
rect 291844 3476 291896 3528
rect 292580 3476 292632 3528
rect 297272 3476 297324 3528
rect 299480 3476 299532 3528
rect 309784 3476 309836 3528
rect 313832 3476 313884 3528
rect 322204 3476 322256 3528
rect 324412 3476 324464 3528
rect 329196 3476 329248 3528
rect 331220 3476 331272 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 582196 3476 582248 3528
rect 582932 3476 582984 3528
rect 18604 3408 18656 3460
rect 24216 3408 24268 3460
rect 50344 3408 50396 3460
rect 64328 3408 64380 3460
rect 64788 3408 64840 3460
rect 72608 3408 72660 3460
rect 92480 3408 92532 3460
rect 118792 3408 118844 3460
rect 141424 3408 141476 3460
rect 188436 3408 188488 3460
rect 242900 3408 242952 3460
rect 246304 3408 246356 3460
rect 253480 3408 253532 3460
rect 256056 3408 256108 3460
rect 265348 3408 265400 3460
rect 267004 3408 267056 3460
rect 271236 3408 271288 3460
rect 315028 3408 315080 3460
rect 327080 3408 327132 3460
rect 330392 3408 330444 3460
rect 338120 3408 338172 3460
rect 351644 3408 351696 3460
rect 357440 3408 357492 3460
rect 1308 3340 1360 3392
rect 7656 3340 7708 3392
rect 12348 3340 12400 3392
rect 289084 3340 289136 3392
rect 294880 3340 294932 3392
rect 345756 3340 345808 3392
rect 351920 3340 351972 3392
rect 272432 3204 272484 3256
rect 277400 3204 277452 3256
rect 56048 3136 56100 3188
rect 58624 3136 58676 3188
rect 65524 3136 65576 3188
rect 66076 3136 66128 3188
rect 80888 3136 80940 3188
rect 83464 3136 83516 3188
rect 299664 3136 299716 3188
rect 302240 3136 302292 3188
rect 302884 3068 302936 3120
rect 305552 3068 305604 3120
rect 17040 3000 17092 3052
rect 22744 3000 22796 3052
rect 27712 3000 27764 3052
rect 29644 3000 29696 3052
rect 93952 3000 94004 3052
rect 95056 3000 95108 3052
rect 250444 3000 250496 3052
rect 252376 3000 252428 3052
rect 581000 2864 581052 2916
rect 583024 2864 583076 2916
rect 129372 2116 129424 2168
rect 136640 2116 136692 2168
rect 51356 2048 51408 2100
rect 195244 2048 195296 2100
rect 240784 2048 240836 2100
rect 300768 2048 300820 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702642 8156 703520
rect 24320 702778 24348 703520
rect 24308 702772 24360 702778
rect 24308 702714 24360 702720
rect 8116 702636 8168 702642
rect 8116 702578 8168 702584
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 18604 683188 18656 683194
rect 18604 683130 18656 683136
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 2792 671090 2820 671191
rect 2780 671084 2832 671090
rect 2780 671026 2832 671032
rect 4804 671084 4856 671090
rect 4804 671026 4856 671032
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3436 576162 3464 632023
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3424 576156 3476 576162
rect 3424 576098 3476 576104
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 554062 3556 566879
rect 3516 554056 3568 554062
rect 3516 553998 3568 554004
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 538286 3464 553823
rect 4816 541113 4844 671026
rect 18616 543046 18644 683130
rect 39304 618316 39356 618322
rect 39304 618258 39356 618264
rect 33140 576156 33192 576162
rect 33140 576098 33192 576104
rect 33152 575550 33180 576098
rect 33140 575544 33192 575550
rect 33140 575486 33192 575492
rect 34428 575544 34480 575550
rect 34428 575486 34480 575492
rect 21364 554056 21416 554062
rect 21364 553998 21416 554004
rect 18604 543040 18656 543046
rect 18604 542982 18656 542988
rect 4802 541104 4858 541113
rect 4802 541039 4858 541048
rect 3424 538280 3476 538286
rect 3424 538222 3476 538228
rect 4804 537532 4856 537538
rect 4804 537474 4856 537480
rect 3424 534132 3476 534138
rect 3424 534074 3476 534080
rect 3436 501809 3464 534074
rect 3514 527912 3570 527921
rect 3514 527847 3516 527856
rect 3568 527847 3570 527856
rect 3516 527818 3568 527824
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 4816 475726 4844 537474
rect 21376 536110 21404 553998
rect 21364 536104 21416 536110
rect 21364 536046 21416 536052
rect 11704 514820 11756 514826
rect 11704 514762 11756 514768
rect 2964 475720 3016 475726
rect 2962 475688 2964 475697
rect 4068 475720 4120 475726
rect 3016 475688 3018 475697
rect 4068 475662 4120 475668
rect 4804 475720 4856 475726
rect 4804 475662 4856 475668
rect 2962 475623 3018 475632
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 2780 423632 2832 423638
rect 2778 423600 2780 423609
rect 2832 423600 2834 423609
rect 2778 423535 2834 423544
rect 2870 410544 2926 410553
rect 2870 410479 2926 410488
rect 2884 409902 2912 410479
rect 2872 409896 2924 409902
rect 2872 409838 2924 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 4080 392193 4108 475662
rect 11716 448526 11744 514762
rect 29644 462392 29696 462398
rect 29644 462334 29696 462340
rect 21364 448588 21416 448594
rect 21364 448530 21416 448536
rect 11704 448520 11756 448526
rect 11704 448462 11756 448468
rect 18604 436144 18656 436150
rect 18604 436086 18656 436092
rect 4804 434784 4856 434790
rect 4804 434726 4856 434732
rect 4816 423638 4844 434726
rect 4804 423632 4856 423638
rect 4804 423574 4856 423580
rect 7564 409896 7616 409902
rect 7564 409838 7616 409844
rect 4066 392184 4122 392193
rect 4066 392119 4122 392128
rect 7576 391921 7604 409838
rect 17222 397488 17278 397497
rect 17222 397423 17278 397432
rect 7562 391912 7618 391921
rect 7562 391847 7618 391856
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 17236 358766 17264 397423
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 17224 358760 17276 358766
rect 17224 358702 17276 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 11704 345092 11756 345098
rect 11704 345034 11756 345040
rect 4804 320884 4856 320890
rect 4804 320826 4856 320832
rect 3882 319288 3938 319297
rect 4816 319258 4844 320826
rect 3882 319223 3884 319232
rect 3936 319223 3938 319232
rect 4804 319252 4856 319258
rect 3884 319194 3936 319200
rect 4804 319194 4856 319200
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3436 286346 3464 306167
rect 3514 293176 3570 293185
rect 3514 293111 3570 293120
rect 3528 292602 3556 293111
rect 3516 292596 3568 292602
rect 3516 292538 3568 292544
rect 3424 286340 3476 286346
rect 3424 286282 3476 286288
rect 3424 280220 3476 280226
rect 3424 280162 3476 280168
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3436 254153 3464 280162
rect 4816 279478 4844 319194
rect 11716 287706 11744 345034
rect 18616 320890 18644 436086
rect 21376 389842 21404 448530
rect 21456 397520 21508 397526
rect 21456 397462 21508 397468
rect 21364 389836 21416 389842
rect 21364 389778 21416 389784
rect 21468 378826 21496 397462
rect 29656 388793 29684 462334
rect 34244 416832 34296 416838
rect 34244 416774 34296 416780
rect 33048 413296 33100 413302
rect 33048 413238 33100 413244
rect 29642 388784 29698 388793
rect 29642 388719 29698 388728
rect 21456 378820 21508 378826
rect 21456 378762 21508 378768
rect 18604 320884 18656 320890
rect 18604 320826 18656 320832
rect 17222 314800 17278 314809
rect 17222 314735 17278 314744
rect 16486 310584 16542 310593
rect 16486 310519 16542 310528
rect 14464 292596 14516 292602
rect 14464 292538 14516 292544
rect 11704 287700 11756 287706
rect 11704 287642 11756 287648
rect 4804 279472 4856 279478
rect 4804 279414 4856 279420
rect 11704 266416 11756 266422
rect 11704 266358 11756 266364
rect 4804 262268 4856 262274
rect 4804 262210 4856 262216
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 4816 241262 4844 262210
rect 2780 241256 2832 241262
rect 2780 241198 2832 241204
rect 4804 241256 4856 241262
rect 4804 241198 4856 241204
rect 2792 241097 2820 241198
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 11716 239426 11744 266358
rect 14476 240786 14504 292538
rect 15844 286340 15896 286346
rect 15844 286282 15896 286288
rect 15856 253910 15884 286282
rect 15844 253904 15896 253910
rect 15844 253846 15896 253852
rect 14464 240780 14516 240786
rect 14464 240722 14516 240728
rect 11704 239420 11756 239426
rect 11704 239362 11756 239368
rect 15106 235240 15162 235249
rect 15106 235175 15162 235184
rect 4804 233912 4856 233918
rect 4804 233854 4856 233860
rect 4066 222864 4122 222873
rect 4066 222799 4122 222808
rect 3146 214976 3202 214985
rect 3146 214911 3202 214920
rect 3160 213994 3188 214911
rect 3148 213988 3200 213994
rect 3148 213930 3200 213936
rect 3240 202156 3292 202162
rect 3240 202098 3292 202104
rect 3252 201929 3280 202098
rect 3238 201920 3294 201929
rect 3238 201855 3294 201864
rect 1308 191140 1360 191146
rect 1308 191082 1360 191088
rect 112 10328 164 10334
rect 112 10270 164 10276
rect 124 490 152 10270
rect 1320 3398 1348 191082
rect 2780 188896 2832 188902
rect 2778 188864 2780 188873
rect 2832 188864 2834 188873
rect 2778 188799 2834 188808
rect 2688 182844 2740 182850
rect 2688 182786 2740 182792
rect 2700 3534 2728 182786
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 2962 149832 3018 149841
rect 2962 149767 3018 149776
rect 2976 149122 3004 149767
rect 2964 149116 3016 149122
rect 2964 149058 3016 149064
rect 3436 141438 3464 162823
rect 3424 141432 3476 141438
rect 3424 141374 3476 141380
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 134564 3476 134570
rect 3424 134506 3476 134512
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3054 97608 3110 97617
rect 3054 97543 3110 97552
rect 3068 96694 3096 97543
rect 3056 96688 3108 96694
rect 3056 96630 3108 96636
rect 3436 58585 3464 134506
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3976 37936 4028 37942
rect 3976 37878 4028 37884
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3436 6497 3464 12378
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3988 3534 4016 37878
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 1308 3392 1360 3398
rect 1308 3334 1360 3340
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 3470
rect 2884 480 2912 3470
rect 4080 480 4108 222799
rect 4816 188902 4844 233854
rect 12348 229764 12400 229770
rect 12348 229706 12400 229712
rect 8208 213920 8260 213926
rect 8208 213862 8260 213868
rect 4804 188896 4856 188902
rect 4804 188838 4856 188844
rect 5446 188320 5502 188329
rect 5446 188255 5502 188264
rect 5356 180124 5408 180130
rect 5356 180066 5408 180072
rect 5368 6914 5396 180066
rect 5276 6886 5396 6914
rect 5276 480 5304 6886
rect 5460 3534 5488 188255
rect 8220 114510 8248 213862
rect 8208 114504 8260 114510
rect 8208 114446 8260 114452
rect 7564 106956 7616 106962
rect 7564 106898 7616 106904
rect 6826 39264 6882 39273
rect 6826 39199 6882 39208
rect 6840 6914 6868 39199
rect 7576 12442 7604 106898
rect 10968 65544 11020 65550
rect 10968 65486 11020 65492
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 6472 6886 6868 6914
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 6472 480 6500 6886
rect 10980 3534 11008 65486
rect 12360 3534 12388 229706
rect 14464 149116 14516 149122
rect 14464 149058 14516 149064
rect 14476 139398 14504 149058
rect 14464 139392 14516 139398
rect 14464 139334 14516 139340
rect 14464 135924 14516 135930
rect 14464 135866 14516 135872
rect 14476 33114 14504 135866
rect 14464 33108 14516 33114
rect 14464 33050 14516 33056
rect 15120 6914 15148 235175
rect 16394 151056 16450 151065
rect 16394 150991 16450 151000
rect 14752 6886 15148 6914
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 8758 3360 8814 3369
rect 7668 480 7696 3334
rect 8758 3295 8814 3304
rect 8772 480 8800 3295
rect 9968 480 9996 3470
rect 11164 480 11192 3470
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12360 480 12388 3334
rect 13556 480 13584 3538
rect 14752 480 14780 6886
rect 16408 3534 16436 150991
rect 16500 4049 16528 310519
rect 16486 4040 16542 4049
rect 16486 3975 16542 3984
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 15948 480 15976 3470
rect 17236 3369 17264 314735
rect 22742 311944 22798 311953
rect 22742 311879 22798 311888
rect 18602 310720 18658 310729
rect 18602 310655 18658 310664
rect 18234 4040 18290 4049
rect 18234 3975 18290 3984
rect 17222 3360 17278 3369
rect 17222 3295 17278 3304
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 17052 480 17080 2994
rect 18248 480 18276 3975
rect 18616 3466 18644 310655
rect 22006 298752 22062 298761
rect 22006 298687 22062 298696
rect 21362 185600 21418 185609
rect 21362 185535 21418 185544
rect 20628 162172 20680 162178
rect 20628 162114 20680 162120
rect 20640 6914 20668 162114
rect 20548 6886 20668 6914
rect 20548 3534 20576 6886
rect 21376 3534 21404 185535
rect 22020 6914 22048 298687
rect 21836 6886 22048 6914
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 19444 480 19472 3470
rect 20640 480 20668 3470
rect 21836 480 21864 6886
rect 22756 3058 22784 311879
rect 29642 309224 29698 309233
rect 29642 309159 29698 309168
rect 26146 306504 26202 306513
rect 26146 306439 26202 306448
rect 23386 33824 23442 33833
rect 23386 33759 23442 33768
rect 23400 6914 23428 33759
rect 23032 6886 23428 6914
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 23032 480 23060 6886
rect 26160 3534 26188 306439
rect 28908 167680 28960 167686
rect 28908 167622 28960 167628
rect 27526 21312 27582 21321
rect 27526 21247 27582 21256
rect 27540 3534 27568 21247
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3470
rect 26528 480 26556 3470
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 480 27752 2994
rect 28920 480 28948 167622
rect 29656 3058 29684 309159
rect 32864 279472 32916 279478
rect 32864 279414 32916 279420
rect 32876 128314 32904 279414
rect 32954 275224 33010 275233
rect 32954 275159 33010 275168
rect 32864 128308 32916 128314
rect 32864 128250 32916 128256
rect 32968 121446 32996 275159
rect 33060 258058 33088 413238
rect 33968 262880 34020 262886
rect 33968 262822 34020 262828
rect 33980 262274 34008 262822
rect 33968 262268 34020 262274
rect 33968 262210 34020 262216
rect 34256 261497 34284 416774
rect 34440 382226 34468 575486
rect 35808 561740 35860 561746
rect 35808 561682 35860 561688
rect 35624 400920 35676 400926
rect 35624 400862 35676 400868
rect 34428 382220 34480 382226
rect 34428 382162 34480 382168
rect 34426 313304 34482 313313
rect 34426 313239 34482 313248
rect 34336 262268 34388 262274
rect 34336 262210 34388 262216
rect 34242 261488 34298 261497
rect 34242 261423 34298 261432
rect 33048 258052 33100 258058
rect 33048 257994 33100 258000
rect 33046 232520 33102 232529
rect 33046 232455 33102 232464
rect 32956 121440 33008 121446
rect 32956 121382 33008 121388
rect 30104 3664 30156 3670
rect 30104 3606 30156 3612
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 30116 480 30144 3606
rect 33060 3534 33088 232455
rect 34348 113150 34376 262210
rect 34336 113144 34388 113150
rect 34336 113086 34388 113092
rect 34440 3534 34468 313239
rect 34520 287700 34572 287706
rect 34520 287642 34572 287648
rect 34532 287094 34560 287642
rect 34520 287088 34572 287094
rect 34520 287030 34572 287036
rect 35636 253910 35664 400862
rect 35820 383654 35848 561682
rect 39316 536790 39344 618258
rect 40052 589966 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 70216 703316 70268 703322
rect 70216 703258 70268 703264
rect 67640 703112 67692 703118
rect 67640 703054 67692 703060
rect 61936 702908 61988 702914
rect 61936 702850 61988 702856
rect 57888 702568 57940 702574
rect 57888 702510 57940 702516
rect 40040 589960 40092 589966
rect 40040 589902 40092 589908
rect 55128 585200 55180 585206
rect 55128 585142 55180 585148
rect 44088 583772 44140 583778
rect 44088 583714 44140 583720
rect 43996 581052 44048 581058
rect 43996 580994 44048 581000
rect 41328 549296 41380 549302
rect 41328 549238 41380 549244
rect 39304 536784 39356 536790
rect 39304 536726 39356 536732
rect 39856 536104 39908 536110
rect 39856 536046 39908 536052
rect 37094 531992 37150 532001
rect 37094 531927 37150 531936
rect 37108 407114 37136 531927
rect 37188 422952 37240 422958
rect 37188 422894 37240 422900
rect 37096 407108 37148 407114
rect 37096 407050 37148 407056
rect 35808 383648 35860 383654
rect 35808 383590 35860 383596
rect 35806 316160 35862 316169
rect 35806 316095 35862 316104
rect 35716 287088 35768 287094
rect 35716 287030 35768 287036
rect 35256 253904 35308 253910
rect 35256 253846 35308 253852
rect 35624 253904 35676 253910
rect 35624 253846 35676 253852
rect 35268 253230 35296 253846
rect 35256 253224 35308 253230
rect 35256 253166 35308 253172
rect 35728 135250 35756 287030
rect 35716 135244 35768 135250
rect 35716 135186 35768 135192
rect 35820 3534 35848 316095
rect 37096 291372 37148 291378
rect 37096 291314 37148 291320
rect 36544 263628 36596 263634
rect 36544 263570 36596 263576
rect 36556 213926 36584 263570
rect 36544 213920 36596 213926
rect 36544 213862 36596 213868
rect 37108 193866 37136 291314
rect 37200 266354 37228 422894
rect 39868 405006 39896 536046
rect 39948 432608 40000 432614
rect 39948 432550 40000 432556
rect 39856 405000 39908 405006
rect 39856 404942 39908 404948
rect 39856 403028 39908 403034
rect 39856 402970 39908 402976
rect 38568 380180 38620 380186
rect 38568 380122 38620 380128
rect 38476 328228 38528 328234
rect 38476 328170 38528 328176
rect 37188 266348 37240 266354
rect 37188 266290 37240 266296
rect 38488 251870 38516 328170
rect 38476 251864 38528 251870
rect 38476 251806 38528 251812
rect 38580 238746 38608 380122
rect 39672 336048 39724 336054
rect 39672 335990 39724 335996
rect 38568 238740 38620 238746
rect 38568 238682 38620 238688
rect 39684 237386 39712 335990
rect 39868 328234 39896 402970
rect 39856 328228 39908 328234
rect 39856 328170 39908 328176
rect 39868 327758 39896 328170
rect 39856 327752 39908 327758
rect 39856 327694 39908 327700
rect 39856 294024 39908 294030
rect 39856 293966 39908 293972
rect 39764 289876 39816 289882
rect 39764 289818 39816 289824
rect 39672 237380 39724 237386
rect 39672 237322 39724 237328
rect 38566 214568 38622 214577
rect 38566 214503 38622 214512
rect 37096 193860 37148 193866
rect 37096 193802 37148 193808
rect 37188 184204 37240 184210
rect 37188 184146 37240 184152
rect 37096 158024 37148 158030
rect 37096 157966 37148 157972
rect 37108 3534 37136 157966
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 35992 3528 36044 3534
rect 35992 3470 36044 3476
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 31298 3360 31354 3369
rect 31298 3295 31354 3304
rect 31312 480 31340 3295
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 36004 480 36032 3470
rect 37200 480 37228 184146
rect 38580 6914 38608 214503
rect 39776 148374 39804 289818
rect 39764 148368 39816 148374
rect 39764 148310 39816 148316
rect 39868 137970 39896 293966
rect 39960 283626 39988 432550
rect 41236 407108 41288 407114
rect 41236 407050 41288 407056
rect 41248 407017 41276 407050
rect 41234 407008 41290 407017
rect 41234 406943 41290 406952
rect 41340 389910 41368 549238
rect 44008 420986 44036 580994
rect 43996 420980 44048 420986
rect 43996 420922 44048 420928
rect 43904 418192 43956 418198
rect 43904 418134 43956 418140
rect 42616 396772 42668 396778
rect 42616 396714 42668 396720
rect 41328 389904 41380 389910
rect 41328 389846 41380 389852
rect 41144 318844 41196 318850
rect 41144 318786 41196 318792
rect 39948 283620 40000 283626
rect 39948 283562 40000 283568
rect 41050 267880 41106 267889
rect 41050 267815 41106 267824
rect 39948 231124 40000 231130
rect 39948 231066 40000 231072
rect 39856 137964 39908 137970
rect 39856 137906 39908 137912
rect 39868 137290 39896 137906
rect 39856 137284 39908 137290
rect 39856 137226 39908 137232
rect 39960 6914 39988 231066
rect 41064 229094 41092 267815
rect 41156 264246 41184 318786
rect 41328 292664 41380 292670
rect 41328 292606 41380 292612
rect 41236 291304 41288 291310
rect 41236 291246 41288 291252
rect 41144 264240 41196 264246
rect 41144 264182 41196 264188
rect 41156 263634 41184 264182
rect 41144 263628 41196 263634
rect 41144 263570 41196 263576
rect 41064 229066 41184 229094
rect 41156 219434 41184 229066
rect 41144 219428 41196 219434
rect 41144 219370 41196 219376
rect 40682 153776 40738 153785
rect 40682 153711 40738 153720
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 40696 3670 40724 153711
rect 40868 135176 40920 135182
rect 40868 135118 40920 135124
rect 40880 134570 40908 135118
rect 40868 134564 40920 134570
rect 40868 134506 40920 134512
rect 41156 118590 41184 219370
rect 41248 144294 41276 291246
rect 41236 144288 41288 144294
rect 41236 144230 41288 144236
rect 41340 135182 41368 292606
rect 42628 247722 42656 396714
rect 43810 338736 43866 338745
rect 43810 338671 43866 338680
rect 42708 330540 42760 330546
rect 42708 330482 42760 330488
rect 42720 258126 42748 330482
rect 42708 258120 42760 258126
rect 42708 258062 42760 258068
rect 42616 247716 42668 247722
rect 42616 247658 42668 247664
rect 42614 216608 42670 216617
rect 42614 216543 42670 216552
rect 41328 135176 41380 135182
rect 41328 135118 41380 135124
rect 41144 118584 41196 118590
rect 41144 118526 41196 118532
rect 41420 107636 41472 107642
rect 41420 107578 41472 107584
rect 41432 106962 41460 107578
rect 41420 106956 41472 106962
rect 41420 106898 41472 106904
rect 42628 96626 42656 216543
rect 42720 107642 42748 258062
rect 43824 232558 43852 338671
rect 43916 321609 43944 418134
rect 44100 387802 44128 583714
rect 50988 582412 51040 582418
rect 50988 582354 51040 582360
rect 46848 580304 46900 580310
rect 46848 580246 46900 580252
rect 46860 579698 46888 580246
rect 46848 579692 46900 579698
rect 46848 579634 46900 579640
rect 46756 440292 46808 440298
rect 46756 440234 46808 440240
rect 45468 425740 45520 425746
rect 45468 425682 45520 425688
rect 44088 387796 44140 387802
rect 44088 387738 44140 387744
rect 43994 384296 44050 384305
rect 43994 384231 44050 384240
rect 43902 321600 43958 321609
rect 43902 321535 43958 321544
rect 43916 284986 43944 321535
rect 43904 284980 43956 284986
rect 43904 284922 43956 284928
rect 43904 276072 43956 276078
rect 43904 276014 43956 276020
rect 43812 232552 43864 232558
rect 43812 232494 43864 232500
rect 43916 126274 43944 276014
rect 44008 239873 44036 384231
rect 45284 339516 45336 339522
rect 45284 339458 45336 339464
rect 44086 284880 44142 284889
rect 44086 284815 44142 284824
rect 43994 239864 44050 239873
rect 43994 239799 44050 239808
rect 43996 155236 44048 155242
rect 43996 155178 44048 155184
rect 43904 126268 43956 126274
rect 43904 126210 43956 126216
rect 42708 107636 42760 107642
rect 42708 107578 42760 107584
rect 42616 96620 42668 96626
rect 42616 96562 42668 96568
rect 42706 35184 42762 35193
rect 42706 35119 42762 35128
rect 41326 22672 41382 22681
rect 41326 22607 41382 22616
rect 40684 3664 40736 3670
rect 40684 3606 40736 3612
rect 41340 3534 41368 22607
rect 42720 3534 42748 35119
rect 44008 3534 44036 155178
rect 44100 132462 44128 284815
rect 45296 234569 45324 339458
rect 45376 285864 45428 285870
rect 45376 285806 45428 285812
rect 45282 234560 45338 234569
rect 45282 234495 45338 234504
rect 45388 140078 45416 285806
rect 45480 267889 45508 425682
rect 46664 388476 46716 388482
rect 46664 388418 46716 388424
rect 45466 267880 45522 267889
rect 45466 267815 45522 267824
rect 45468 260160 45520 260166
rect 45468 260102 45520 260108
rect 45376 140072 45428 140078
rect 45376 140014 45428 140020
rect 44824 135312 44876 135318
rect 44824 135254 44876 135260
rect 44088 132456 44140 132462
rect 44088 132398 44140 132404
rect 44836 111790 44864 135254
rect 44824 111784 44876 111790
rect 44824 111726 44876 111732
rect 45480 109750 45508 260102
rect 45560 258188 45612 258194
rect 45560 258130 45612 258136
rect 46204 258188 46256 258194
rect 46204 258130 46256 258136
rect 45572 258058 45600 258130
rect 45560 258052 45612 258058
rect 45560 257994 45612 258000
rect 45928 251864 45980 251870
rect 45928 251806 45980 251812
rect 45940 251258 45968 251806
rect 45928 251252 45980 251258
rect 45928 251194 45980 251200
rect 46216 196994 46244 258130
rect 46676 241466 46704 388418
rect 46768 289814 46796 440234
rect 46860 386374 46888 579634
rect 49608 565888 49660 565894
rect 49608 565830 49660 565836
rect 48228 560312 48280 560318
rect 48228 560254 48280 560260
rect 48136 539640 48188 539646
rect 48136 539582 48188 539588
rect 48044 395344 48096 395350
rect 48044 395286 48096 395292
rect 46848 386368 46900 386374
rect 46848 386310 46900 386316
rect 46756 289808 46808 289814
rect 46756 289750 46808 289756
rect 47860 283008 47912 283014
rect 47860 282950 47912 282956
rect 46848 251252 46900 251258
rect 46848 251194 46900 251200
rect 46664 241460 46716 241466
rect 46664 241402 46716 241408
rect 46756 197328 46808 197334
rect 46756 197270 46808 197276
rect 46768 196994 46796 197270
rect 46204 196988 46256 196994
rect 46204 196930 46256 196936
rect 46756 196988 46808 196994
rect 46756 196930 46808 196936
rect 46768 110430 46796 196930
rect 46756 110424 46808 110430
rect 46756 110366 46808 110372
rect 45468 109744 45520 109750
rect 45468 109686 45520 109692
rect 46860 101454 46888 251194
rect 47872 133890 47900 282950
rect 48056 244497 48084 395286
rect 48148 391270 48176 539582
rect 48240 511290 48268 560254
rect 48228 511284 48280 511290
rect 48228 511226 48280 511232
rect 48240 439550 48268 511226
rect 48228 439544 48280 439550
rect 48228 439486 48280 439492
rect 48228 420980 48280 420986
rect 48228 420922 48280 420928
rect 48136 391264 48188 391270
rect 48136 391206 48188 391212
rect 48136 376032 48188 376038
rect 48136 375974 48188 375980
rect 48148 281518 48176 375974
rect 48136 281512 48188 281518
rect 48136 281454 48188 281460
rect 48240 265033 48268 420922
rect 49516 414044 49568 414050
rect 49516 413986 49568 413992
rect 49528 324358 49556 413986
rect 49620 409902 49648 565830
rect 50896 546508 50948 546514
rect 50896 546450 50948 546456
rect 49608 409896 49660 409902
rect 49608 409838 49660 409844
rect 50804 408536 50856 408542
rect 50804 408478 50856 408484
rect 49606 393544 49662 393553
rect 49606 393479 49662 393488
rect 49516 324352 49568 324358
rect 49516 324294 49568 324300
rect 48226 265024 48282 265033
rect 48226 264959 48282 264968
rect 48042 244488 48098 244497
rect 48042 244423 48098 244432
rect 47950 237416 48006 237425
rect 47950 237351 48006 237360
rect 47860 133884 47912 133890
rect 47860 133826 47912 133832
rect 47964 115938 47992 237351
rect 48056 216617 48084 244423
rect 48240 238649 48268 264959
rect 49528 260846 49556 324294
rect 49516 260840 49568 260846
rect 49516 260782 49568 260788
rect 49528 260166 49556 260782
rect 49516 260160 49568 260166
rect 49516 260102 49568 260108
rect 49424 255332 49476 255338
rect 49424 255274 49476 255280
rect 48226 238640 48282 238649
rect 48226 238575 48282 238584
rect 48240 237425 48268 238575
rect 48226 237416 48282 237425
rect 48226 237351 48282 237360
rect 49436 223553 49464 255274
rect 49514 254552 49570 254561
rect 49514 254487 49570 254496
rect 49528 253978 49556 254487
rect 49516 253972 49568 253978
rect 49516 253914 49568 253920
rect 49422 223544 49478 223553
rect 49422 223479 49478 223488
rect 48042 216608 48098 216617
rect 48042 216543 48098 216552
rect 48044 211812 48096 211818
rect 48044 211754 48096 211760
rect 47952 115932 48004 115938
rect 47952 115874 48004 115880
rect 46848 101448 46900 101454
rect 46848 101390 46900 101396
rect 48056 89690 48084 211754
rect 49528 209681 49556 253914
rect 49620 242962 49648 393479
rect 50710 285832 50766 285841
rect 50710 285767 50766 285776
rect 50344 266348 50396 266354
rect 50344 266290 50396 266296
rect 49608 242956 49660 242962
rect 49608 242898 49660 242904
rect 49606 223544 49662 223553
rect 49606 223479 49662 223488
rect 49514 209672 49570 209681
rect 49514 209607 49570 209616
rect 48226 146976 48282 146985
rect 48226 146911 48282 146920
rect 48044 89684 48096 89690
rect 48044 89626 48096 89632
rect 48136 78056 48188 78062
rect 48136 77998 48188 78004
rect 45466 36544 45522 36553
rect 45466 36479 45522 36488
rect 45376 13116 45428 13122
rect 45376 13058 45428 13064
rect 45388 3534 45416 13058
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41328 3528 41380 3534
rect 41328 3470 41380 3476
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 43996 3528 44048 3534
rect 43996 3470 44048 3476
rect 44272 3528 44324 3534
rect 44272 3470 44324 3476
rect 45376 3528 45428 3534
rect 45376 3470 45428 3476
rect 40696 480 40724 3470
rect 41892 480 41920 3470
rect 43088 480 43116 3470
rect 44284 480 44312 3470
rect 45480 480 45508 36479
rect 46664 14476 46716 14482
rect 46664 14418 46716 14424
rect 46676 480 46704 14418
rect 48148 6914 48176 77998
rect 47872 6886 48176 6914
rect 47872 480 47900 6886
rect 48240 3534 48268 146911
rect 49528 106282 49556 209607
rect 49620 107574 49648 223479
rect 50356 222154 50384 266290
rect 50344 222148 50396 222154
rect 50344 222090 50396 222096
rect 50724 220833 50752 285767
rect 50816 256698 50844 408478
rect 50908 389201 50936 546450
rect 51000 442270 51028 582354
rect 53746 578912 53802 578921
rect 53746 578847 53802 578856
rect 52368 564392 52420 564398
rect 52368 564334 52420 564340
rect 50988 442264 51040 442270
rect 50988 442206 51040 442212
rect 52380 440910 52408 564334
rect 53656 557592 53708 557598
rect 53656 557534 53708 557540
rect 53668 449206 53696 557534
rect 53656 449200 53708 449206
rect 53656 449142 53708 449148
rect 52368 440904 52420 440910
rect 52368 440846 52420 440852
rect 52380 440298 52408 440846
rect 52368 440292 52420 440298
rect 52368 440234 52420 440240
rect 52182 436248 52238 436257
rect 52182 436183 52238 436192
rect 50988 434852 51040 434858
rect 50988 434794 51040 434800
rect 50894 389192 50950 389201
rect 50894 389127 50950 389136
rect 50894 387696 50950 387705
rect 50894 387631 50950 387640
rect 50804 256692 50856 256698
rect 50804 256634 50856 256640
rect 50816 255338 50844 256634
rect 50804 255332 50856 255338
rect 50804 255274 50856 255280
rect 50908 248414 50936 387631
rect 51000 278050 51028 434794
rect 52196 306377 52224 436183
rect 53760 434042 53788 578847
rect 55036 544400 55088 544406
rect 55036 544342 55088 544348
rect 55048 438190 55076 544342
rect 55036 438184 55088 438190
rect 55036 438126 55088 438132
rect 53748 434036 53800 434042
rect 53748 433978 53800 433984
rect 53562 433664 53618 433673
rect 53562 433599 53618 433608
rect 52368 423700 52420 423706
rect 52368 423642 52420 423648
rect 52276 409896 52328 409902
rect 52276 409838 52328 409844
rect 52182 306368 52238 306377
rect 52182 306303 52238 306312
rect 52196 305017 52224 306303
rect 52182 305008 52238 305017
rect 52182 304943 52238 304952
rect 52184 289808 52236 289814
rect 52184 289750 52236 289756
rect 52196 288454 52224 289750
rect 52184 288448 52236 288454
rect 52184 288390 52236 288396
rect 52092 284368 52144 284374
rect 52092 284310 52144 284316
rect 50988 278044 51040 278050
rect 50988 277986 51040 277992
rect 50908 248386 51028 248414
rect 51000 235890 51028 248386
rect 50988 235884 51040 235890
rect 50988 235826 51040 235832
rect 50896 222148 50948 222154
rect 50896 222090 50948 222096
rect 50710 220824 50766 220833
rect 50710 220759 50766 220768
rect 50724 219434 50752 220759
rect 50724 219406 50844 219434
rect 50342 149696 50398 149705
rect 50342 149631 50398 149640
rect 49608 107568 49660 107574
rect 49608 107510 49660 107516
rect 49516 106276 49568 106282
rect 49516 106218 49568 106224
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 50356 3466 50384 149631
rect 50816 145586 50844 219406
rect 50804 145580 50856 145586
rect 50804 145522 50856 145528
rect 50908 117298 50936 222090
rect 51000 198694 51028 235826
rect 52104 228993 52132 284310
rect 52090 228984 52146 228993
rect 52090 228919 52146 228928
rect 50988 198688 51040 198694
rect 50988 198630 51040 198636
rect 50896 117292 50948 117298
rect 50896 117234 50948 117240
rect 51000 90817 51028 198630
rect 52104 137329 52132 228919
rect 52196 226302 52224 288390
rect 52288 257378 52316 409838
rect 52380 268394 52408 423642
rect 53576 336802 53604 433599
rect 53656 429208 53708 429214
rect 53656 429150 53708 429156
rect 53564 336796 53616 336802
rect 53564 336738 53616 336744
rect 53472 329860 53524 329866
rect 53472 329802 53524 329808
rect 52460 283620 52512 283626
rect 52460 283562 52512 283568
rect 52472 282198 52500 283562
rect 52460 282192 52512 282198
rect 52460 282134 52512 282140
rect 53104 281512 53156 281518
rect 53104 281454 53156 281460
rect 52458 276176 52514 276185
rect 52458 276111 52514 276120
rect 52472 276078 52500 276111
rect 52460 276072 52512 276078
rect 52460 276014 52512 276020
rect 52368 268388 52420 268394
rect 52368 268330 52420 268336
rect 52276 257372 52328 257378
rect 52276 257314 52328 257320
rect 52184 226296 52236 226302
rect 52184 226238 52236 226244
rect 52182 224904 52238 224913
rect 52288 224890 52316 257314
rect 52460 247716 52512 247722
rect 52460 247658 52512 247664
rect 52472 247217 52500 247658
rect 52458 247208 52514 247217
rect 52458 247143 52514 247152
rect 52368 239420 52420 239426
rect 52368 239362 52420 239368
rect 52238 224862 52316 224890
rect 52182 224839 52238 224848
rect 52090 137320 52146 137329
rect 52090 137255 52146 137264
rect 52196 109002 52224 224839
rect 52276 224256 52328 224262
rect 52276 224198 52328 224204
rect 52184 108996 52236 109002
rect 52184 108938 52236 108944
rect 50986 90808 51042 90817
rect 50986 90743 51042 90752
rect 52288 89622 52316 224198
rect 52380 92478 52408 239362
rect 53116 238678 53144 281454
rect 53484 271969 53512 329802
rect 53576 282169 53604 336738
rect 53668 329866 53696 429150
rect 53746 420200 53802 420209
rect 53746 420135 53802 420144
rect 53656 329860 53708 329866
rect 53656 329802 53708 329808
rect 53760 300830 53788 420135
rect 54852 414112 54904 414118
rect 54852 414054 54904 414060
rect 53840 389904 53892 389910
rect 53840 389846 53892 389852
rect 53852 389230 53880 389846
rect 53840 389224 53892 389230
rect 53840 389166 53892 389172
rect 54760 389224 54812 389230
rect 54760 389166 54812 389172
rect 53748 300824 53800 300830
rect 53748 300766 53800 300772
rect 53656 282192 53708 282198
rect 53562 282160 53618 282169
rect 53656 282134 53708 282140
rect 53562 282095 53618 282104
rect 53470 271960 53526 271969
rect 53470 271895 53526 271904
rect 53484 258074 53512 271895
rect 53392 258046 53512 258074
rect 53104 238672 53156 238678
rect 53104 238614 53156 238620
rect 53392 122806 53420 258046
rect 53562 247208 53618 247217
rect 53562 247143 53618 247152
rect 53576 219434 53604 247143
rect 53484 219406 53604 219434
rect 53484 218006 53512 219406
rect 53472 218000 53524 218006
rect 53472 217942 53524 217948
rect 53380 122800 53432 122806
rect 53380 122742 53432 122748
rect 53484 99346 53512 217942
rect 53564 144220 53616 144226
rect 53564 144162 53616 144168
rect 53472 99340 53524 99346
rect 53472 99282 53524 99288
rect 52368 92472 52420 92478
rect 52368 92414 52420 92420
rect 52276 89616 52328 89622
rect 52276 89558 52328 89564
rect 50988 18624 51040 18630
rect 50988 18566 51040 18572
rect 51000 3534 51028 18566
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 50344 3460 50396 3466
rect 50344 3402 50396 3408
rect 51356 2100 51408 2106
rect 51356 2042 51408 2048
rect 51368 480 51396 2042
rect 52564 480 52592 3538
rect 53576 3482 53604 144162
rect 53668 132394 53696 282134
rect 53760 267714 53788 300766
rect 53748 267708 53800 267714
rect 53748 267650 53800 267656
rect 54772 242214 54800 389166
rect 54864 264217 54892 414054
rect 55036 398880 55088 398886
rect 55036 398822 55088 398828
rect 54944 271856 54996 271862
rect 54944 271798 54996 271804
rect 54850 264208 54906 264217
rect 54850 264143 54906 264152
rect 54760 242208 54812 242214
rect 54760 242150 54812 242156
rect 54956 211070 54984 271798
rect 55048 248418 55076 398822
rect 55140 387977 55168 585142
rect 56508 570648 56560 570654
rect 56508 570590 56560 570596
rect 56416 426488 56468 426494
rect 56416 426430 56468 426436
rect 55126 387968 55182 387977
rect 55126 387903 55182 387912
rect 55128 387796 55180 387802
rect 55128 387738 55180 387744
rect 55140 386481 55168 387738
rect 55126 386472 55182 386481
rect 55126 386407 55182 386416
rect 56232 320204 56284 320210
rect 56232 320146 56284 320152
rect 55218 248432 55274 248441
rect 55048 248390 55218 248418
rect 55218 248367 55274 248376
rect 55128 244928 55180 244934
rect 55128 244870 55180 244876
rect 55036 242956 55088 242962
rect 55036 242898 55088 242904
rect 54944 211064 54996 211070
rect 54944 211006 54996 211012
rect 54852 142860 54904 142866
rect 54852 142802 54904 142808
rect 53656 132388 53708 132394
rect 53656 132330 53708 132336
rect 54864 92818 54892 142802
rect 54956 120086 54984 211006
rect 55048 194546 55076 242898
rect 55140 212498 55168 244870
rect 56244 240106 56272 320146
rect 56324 288516 56376 288522
rect 56324 288458 56376 288464
rect 55956 240100 56008 240106
rect 55956 240042 56008 240048
rect 56232 240100 56284 240106
rect 56232 240042 56284 240048
rect 55968 239426 55996 240042
rect 55956 239420 56008 239426
rect 55956 239362 56008 239368
rect 55128 212492 55180 212498
rect 55128 212434 55180 212440
rect 55036 194540 55088 194546
rect 55036 194482 55088 194488
rect 54944 120080 54996 120086
rect 54944 120022 54996 120028
rect 55048 95198 55076 194482
rect 55140 97306 55168 212434
rect 56336 199442 56364 288458
rect 56428 271862 56456 426430
rect 56520 406994 56548 570590
rect 57900 564398 57928 702510
rect 59266 581088 59322 581097
rect 59266 581023 59322 581032
rect 57888 564392 57940 564398
rect 57888 564334 57940 564340
rect 57888 554804 57940 554810
rect 57888 554746 57940 554752
rect 57244 553444 57296 553450
rect 57244 553386 57296 553392
rect 57256 416838 57284 553386
rect 57520 431996 57572 432002
rect 57520 431938 57572 431944
rect 57244 416832 57296 416838
rect 57244 416774 57296 416780
rect 56598 407008 56654 407017
rect 56520 406966 56598 406994
rect 56598 406943 56654 406952
rect 56508 400240 56560 400246
rect 56508 400182 56560 400188
rect 56520 302258 56548 400182
rect 56508 302252 56560 302258
rect 56508 302194 56560 302200
rect 56416 271856 56468 271862
rect 56416 271798 56468 271804
rect 56414 264208 56470 264217
rect 56414 264143 56470 264152
rect 56428 261526 56456 264143
rect 56416 261520 56468 261526
rect 56416 261462 56468 261468
rect 56428 206990 56456 261462
rect 56520 249830 56548 302194
rect 57532 275913 57560 431938
rect 57704 392012 57756 392018
rect 57704 391954 57756 391960
rect 57716 331265 57744 391954
rect 57900 384334 57928 554746
rect 58990 533352 59046 533361
rect 58990 533287 59046 533296
rect 58900 430636 58952 430642
rect 58900 430578 58952 430584
rect 57888 384328 57940 384334
rect 57888 384270 57940 384276
rect 57702 331256 57758 331265
rect 57702 331191 57758 331200
rect 57612 295996 57664 296002
rect 57612 295938 57664 295944
rect 57518 275904 57574 275913
rect 57518 275839 57574 275848
rect 57532 275233 57560 275839
rect 57518 275224 57574 275233
rect 57518 275159 57574 275168
rect 56508 249824 56560 249830
rect 56508 249766 56560 249772
rect 56506 248432 56562 248441
rect 56506 248367 56562 248376
rect 56416 206984 56468 206990
rect 56416 206926 56468 206932
rect 56324 199436 56376 199442
rect 56324 199378 56376 199384
rect 56324 140140 56376 140146
rect 56324 140082 56376 140088
rect 55128 97300 55180 97306
rect 55128 97242 55180 97248
rect 55036 95192 55088 95198
rect 55036 95134 55088 95140
rect 54852 92812 54904 92818
rect 54852 92754 54904 92760
rect 54482 91760 54538 91769
rect 54482 91695 54538 91704
rect 53746 24168 53802 24177
rect 53746 24103 53802 24112
rect 53760 6914 53788 24103
rect 53668 6886 53788 6914
rect 53668 3602 53696 6886
rect 53656 3596 53708 3602
rect 53656 3538 53708 3544
rect 53576 3454 53788 3482
rect 53760 480 53788 3454
rect 54496 3369 54524 91695
rect 56336 84182 56364 140082
rect 56428 111790 56456 206926
rect 56416 111784 56468 111790
rect 56416 111726 56468 111732
rect 56520 99550 56548 248367
rect 57624 241534 57652 295938
rect 57716 246265 57744 331191
rect 57888 279608 57940 279614
rect 57888 279550 57940 279556
rect 57796 274712 57848 274718
rect 57796 274654 57848 274660
rect 57702 246256 57758 246265
rect 57702 246191 57758 246200
rect 57612 241528 57664 241534
rect 57612 241470 57664 241476
rect 57704 228404 57756 228410
rect 57704 228346 57756 228352
rect 57610 222184 57666 222193
rect 57610 222119 57666 222128
rect 57060 109744 57112 109750
rect 57060 109686 57112 109692
rect 57072 109070 57100 109686
rect 56600 109064 56652 109070
rect 56600 109006 56652 109012
rect 57060 109064 57112 109070
rect 57060 109006 57112 109012
rect 56508 99544 56560 99550
rect 56508 99486 56560 99492
rect 56612 85542 56640 109006
rect 57624 108934 57652 222119
rect 57716 205601 57744 228346
rect 57702 205592 57758 205601
rect 57702 205527 57758 205536
rect 57612 108928 57664 108934
rect 57612 108870 57664 108876
rect 57716 90953 57744 205527
rect 57808 125594 57836 274654
rect 57900 129062 57928 279550
rect 58912 274650 58940 430578
rect 59004 393553 59032 533287
rect 59280 413302 59308 581023
rect 60648 558952 60700 558958
rect 60648 558894 60700 558900
rect 60556 429276 60608 429282
rect 60556 429218 60608 429224
rect 60464 419552 60516 419558
rect 60464 419494 60516 419500
rect 59268 413296 59320 413302
rect 59268 413238 59320 413244
rect 59084 405000 59136 405006
rect 59084 404942 59136 404948
rect 59096 396166 59124 404942
rect 59084 396160 59136 396166
rect 59084 396102 59136 396108
rect 58990 393544 59046 393553
rect 58990 393479 59046 393488
rect 58992 287700 59044 287706
rect 58992 287642 59044 287648
rect 58900 274644 58952 274650
rect 58900 274586 58952 274592
rect 58912 274174 58940 274586
rect 58900 274168 58952 274174
rect 58900 274110 58952 274116
rect 59004 220114 59032 287642
rect 59096 246158 59124 396102
rect 60372 304292 60424 304298
rect 60372 304234 60424 304240
rect 60384 279478 60412 304234
rect 60476 292602 60504 419494
rect 60464 292596 60516 292602
rect 60464 292538 60516 292544
rect 60462 283520 60518 283529
rect 60462 283455 60518 283464
rect 60372 279472 60424 279478
rect 60372 279414 60424 279420
rect 59176 278044 59228 278050
rect 59176 277986 59228 277992
rect 59084 246152 59136 246158
rect 59084 246094 59136 246100
rect 59188 238754 59216 277986
rect 59268 274168 59320 274174
rect 59268 274110 59320 274116
rect 59096 238726 59216 238754
rect 59096 237289 59124 238726
rect 59082 237280 59138 237289
rect 59082 237215 59138 237224
rect 58992 220108 59044 220114
rect 58992 220050 59044 220056
rect 58992 160744 59044 160750
rect 58992 160686 59044 160692
rect 57888 129056 57940 129062
rect 57888 128998 57940 129004
rect 57796 125588 57848 125594
rect 57796 125530 57848 125536
rect 57702 90944 57758 90953
rect 57702 90879 57758 90888
rect 58622 89040 58678 89049
rect 58622 88975 58678 88984
rect 57886 86320 57942 86329
rect 57886 86255 57942 86264
rect 56600 85536 56652 85542
rect 56600 85478 56652 85484
rect 56324 84176 56376 84182
rect 56324 84118 56376 84124
rect 54944 7608 54996 7614
rect 54944 7550 54996 7556
rect 54482 3360 54538 3369
rect 54482 3295 54538 3304
rect 54956 480 54984 7550
rect 57900 3534 57928 86255
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 56048 3188 56100 3194
rect 56048 3130 56100 3136
rect 56060 480 56088 3130
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 58636 3194 58664 88975
rect 59004 88233 59032 160686
rect 59096 128246 59124 237215
rect 59176 196648 59228 196654
rect 59176 196590 59228 196596
rect 59084 128240 59136 128246
rect 59084 128182 59136 128188
rect 59188 88330 59216 196590
rect 59280 124166 59308 274110
rect 60370 254008 60426 254017
rect 60370 253943 60426 253952
rect 60384 229094 60412 253943
rect 60476 236706 60504 283455
rect 60568 273329 60596 429218
rect 60660 396778 60688 558894
rect 61948 544406 61976 702850
rect 66168 702500 66220 702506
rect 66168 702442 66220 702448
rect 62028 582480 62080 582486
rect 62028 582422 62080 582428
rect 61936 544400 61988 544406
rect 61936 544342 61988 544348
rect 61936 530596 61988 530602
rect 61936 530538 61988 530544
rect 61948 423502 61976 530538
rect 60740 423496 60792 423502
rect 60740 423438 60792 423444
rect 61936 423496 61988 423502
rect 61936 423438 61988 423444
rect 60752 422958 60780 423438
rect 60740 422952 60792 422958
rect 60740 422894 60792 422900
rect 61934 418296 61990 418305
rect 61934 418231 61990 418240
rect 60648 396772 60700 396778
rect 60648 396714 60700 396720
rect 61842 318064 61898 318073
rect 61842 317999 61898 318008
rect 60648 292596 60700 292602
rect 60648 292538 60700 292544
rect 60554 273320 60610 273329
rect 60554 273255 60610 273264
rect 60554 269240 60610 269249
rect 60554 269175 60610 269184
rect 60464 236700 60516 236706
rect 60464 236642 60516 236648
rect 60384 229066 60504 229094
rect 60476 226273 60504 229066
rect 60462 226264 60518 226273
rect 60462 226199 60518 226208
rect 60372 138712 60424 138718
rect 60372 138654 60424 138660
rect 59268 124160 59320 124166
rect 59268 124102 59320 124108
rect 59176 88324 59228 88330
rect 59176 88266 59228 88272
rect 60384 88262 60412 138654
rect 60476 104854 60504 226199
rect 60568 120222 60596 269175
rect 60660 265198 60688 292538
rect 60740 284980 60792 284986
rect 60740 284922 60792 284928
rect 60648 265192 60700 265198
rect 60648 265134 60700 265140
rect 60556 120216 60608 120222
rect 60556 120158 60608 120164
rect 60660 114646 60688 265134
rect 60752 262886 60780 284922
rect 61856 284889 61884 317999
rect 61948 295361 61976 418231
rect 62040 389337 62068 582422
rect 64696 579692 64748 579698
rect 64696 579634 64748 579640
rect 63408 564460 63460 564466
rect 63408 564402 63460 564408
rect 63224 434036 63276 434042
rect 63224 433978 63276 433984
rect 62026 389328 62082 389337
rect 62026 389263 62082 389272
rect 63236 328438 63264 433978
rect 63316 403028 63368 403034
rect 63316 402970 63368 402976
rect 63224 328432 63276 328438
rect 63224 328374 63276 328380
rect 63224 316736 63276 316742
rect 63224 316678 63276 316684
rect 62028 304972 62080 304978
rect 62028 304914 62080 304920
rect 61934 295352 61990 295361
rect 61934 295287 61990 295296
rect 61842 284880 61898 284889
rect 61842 284815 61898 284824
rect 61750 270736 61806 270745
rect 61750 270671 61806 270680
rect 60740 262880 60792 262886
rect 60740 262822 60792 262828
rect 61568 250504 61620 250510
rect 61568 250446 61620 250452
rect 61580 249762 61608 250446
rect 61568 249756 61620 249762
rect 61568 249698 61620 249704
rect 60648 114640 60700 114646
rect 60648 114582 60700 114588
rect 60464 104848 60516 104854
rect 60464 104790 60516 104796
rect 60740 101448 60792 101454
rect 60740 101390 60792 101396
rect 60372 88256 60424 88262
rect 58990 88224 59046 88233
rect 60372 88198 60424 88204
rect 58990 88159 59046 88168
rect 59268 50448 59320 50454
rect 59268 50390 59320 50396
rect 59280 3534 59308 50390
rect 60752 45558 60780 101390
rect 61580 100706 61608 249698
rect 61764 209774 61792 270671
rect 61948 263673 61976 295287
rect 61934 263664 61990 263673
rect 61934 263599 61990 263608
rect 61842 252784 61898 252793
rect 61842 252719 61898 252728
rect 61672 209746 61792 209774
rect 61856 209774 61884 252719
rect 62040 247110 62068 304914
rect 63130 287328 63186 287337
rect 63130 287263 63186 287272
rect 62854 273184 62910 273193
rect 62854 273119 62910 273128
rect 62868 272134 62896 273119
rect 62856 272128 62908 272134
rect 62856 272070 62908 272076
rect 63144 261594 63172 287263
rect 63236 285666 63264 316678
rect 63224 285660 63276 285666
rect 63224 285602 63276 285608
rect 63224 272128 63276 272134
rect 63224 272070 63276 272076
rect 63132 261588 63184 261594
rect 63132 261530 63184 261536
rect 62028 247104 62080 247110
rect 62028 247046 62080 247052
rect 61856 209746 61976 209774
rect 61672 208350 61700 209746
rect 61660 208344 61712 208350
rect 61660 208286 61712 208292
rect 61672 122738 61700 208286
rect 61948 205630 61976 209746
rect 61936 205624 61988 205630
rect 61936 205566 61988 205572
rect 61752 155304 61804 155310
rect 61752 155246 61804 155252
rect 61660 122732 61712 122738
rect 61660 122674 61712 122680
rect 61568 100700 61620 100706
rect 61568 100642 61620 100648
rect 61764 86902 61792 155246
rect 61948 103494 61976 205566
rect 63236 151814 63264 272070
rect 63328 251297 63356 402970
rect 63420 391338 63448 564402
rect 64708 479534 64736 579634
rect 64788 571396 64840 571402
rect 64788 571338 64840 571344
rect 64696 479528 64748 479534
rect 64696 479470 64748 479476
rect 64696 476808 64748 476814
rect 64696 476750 64748 476756
rect 64144 418192 64196 418198
rect 64144 418134 64196 418140
rect 63408 391332 63460 391338
rect 63408 391274 63460 391280
rect 63408 328432 63460 328438
rect 63408 328374 63460 328380
rect 63420 327146 63448 328374
rect 63408 327140 63460 327146
rect 63408 327082 63460 327088
rect 63420 276010 63448 327082
rect 64156 318850 64184 418134
rect 64708 395350 64736 476750
rect 64800 458862 64828 571338
rect 66074 567624 66130 567633
rect 66074 567559 66130 567568
rect 65984 545148 66036 545154
rect 65984 545090 66036 545096
rect 65996 485110 66024 545090
rect 65984 485104 66036 485110
rect 65984 485046 66036 485052
rect 66088 475386 66116 567559
rect 66180 545986 66208 702442
rect 66534 580000 66590 580009
rect 66534 579935 66590 579944
rect 66548 579698 66576 579935
rect 66536 579692 66588 579698
rect 66536 579634 66588 579640
rect 66902 578640 66958 578649
rect 66902 578575 66958 578584
rect 66442 575920 66498 575929
rect 66442 575855 66498 575864
rect 66456 575550 66484 575855
rect 66444 575544 66496 575550
rect 66444 575486 66496 575492
rect 66626 573200 66682 573209
rect 66626 573135 66682 573144
rect 66640 570654 66668 573135
rect 66718 571840 66774 571849
rect 66718 571775 66774 571784
rect 66732 571402 66760 571775
rect 66720 571396 66772 571402
rect 66720 571338 66772 571344
rect 66628 570648 66680 570654
rect 66628 570590 66680 570596
rect 66810 564768 66866 564777
rect 66810 564703 66866 564712
rect 66824 564466 66852 564703
rect 66812 564460 66864 564466
rect 66812 564402 66864 564408
rect 66536 564392 66588 564398
rect 66536 564334 66588 564340
rect 66548 564233 66576 564334
rect 66534 564224 66590 564233
rect 66534 564159 66590 564168
rect 66810 562048 66866 562057
rect 66810 561983 66866 561992
rect 66824 561746 66852 561983
rect 66812 561740 66864 561746
rect 66812 561682 66864 561688
rect 66810 560688 66866 560697
rect 66810 560623 66866 560632
rect 66824 560318 66852 560623
rect 66812 560312 66864 560318
rect 66812 560254 66864 560260
rect 66810 559328 66866 559337
rect 66810 559263 66866 559272
rect 66824 558958 66852 559263
rect 66812 558952 66864 558958
rect 66812 558894 66864 558900
rect 66810 557968 66866 557977
rect 66810 557903 66866 557912
rect 66824 557598 66852 557903
rect 66812 557592 66864 557598
rect 66812 557534 66864 557540
rect 66718 555248 66774 555257
rect 66718 555183 66774 555192
rect 66732 554810 66760 555183
rect 66720 554804 66772 554810
rect 66720 554746 66772 554752
rect 66810 553616 66866 553625
rect 66810 553551 66866 553560
rect 66824 553450 66852 553551
rect 66812 553444 66864 553450
rect 66812 553386 66864 553392
rect 66810 549536 66866 549545
rect 66810 549471 66866 549480
rect 66824 549302 66852 549471
rect 66812 549296 66864 549302
rect 66812 549238 66864 549244
rect 66534 546816 66590 546825
rect 66534 546751 66590 546760
rect 66548 546514 66576 546751
rect 66536 546508 66588 546514
rect 66536 546450 66588 546456
rect 66258 546000 66314 546009
rect 66180 545958 66258 545986
rect 66180 545154 66208 545958
rect 66258 545935 66314 545944
rect 66168 545148 66220 545154
rect 66168 545090 66220 545096
rect 66350 544504 66406 544513
rect 66350 544439 66406 544448
rect 66364 544406 66392 544439
rect 66352 544400 66404 544406
rect 66352 544342 66404 544348
rect 66626 543144 66682 543153
rect 66626 543079 66682 543088
rect 66640 543046 66668 543079
rect 66168 543040 66220 543046
rect 66168 542982 66220 542988
rect 66628 543040 66680 543046
rect 66628 542982 66680 542988
rect 66076 475380 66128 475386
rect 66076 475322 66128 475328
rect 65984 474088 66036 474094
rect 65984 474030 66036 474036
rect 64788 458856 64840 458862
rect 64788 458798 64840 458804
rect 64788 456068 64840 456074
rect 64788 456010 64840 456016
rect 64800 411369 64828 456010
rect 65892 444780 65944 444786
rect 65892 444722 65944 444728
rect 65904 425746 65932 444722
rect 65892 425740 65944 425746
rect 65892 425682 65944 425688
rect 64786 411360 64842 411369
rect 64786 411295 64842 411304
rect 64788 404388 64840 404394
rect 64788 404330 64840 404336
rect 64696 395344 64748 395350
rect 64696 395286 64748 395292
rect 64604 393372 64656 393378
rect 64604 393314 64656 393320
rect 63500 318844 63552 318850
rect 63500 318786 63552 318792
rect 64144 318844 64196 318850
rect 64144 318786 64196 318792
rect 63512 318102 63540 318786
rect 63500 318096 63552 318102
rect 63500 318038 63552 318044
rect 64144 285660 64196 285666
rect 64144 285602 64196 285608
rect 63408 276004 63460 276010
rect 63408 275946 63460 275952
rect 63420 274718 63448 275946
rect 63408 274712 63460 274718
rect 63408 274654 63460 274660
rect 63406 263528 63462 263537
rect 63406 263463 63462 263472
rect 63314 251288 63370 251297
rect 63314 251223 63370 251232
rect 63144 151786 63264 151814
rect 63144 149054 63172 151786
rect 63132 149048 63184 149054
rect 63132 148990 63184 148996
rect 63144 120193 63172 148990
rect 63314 135960 63370 135969
rect 63314 135895 63370 135904
rect 63224 124160 63276 124166
rect 63224 124102 63276 124108
rect 63236 122942 63264 124102
rect 63224 122936 63276 122942
rect 63224 122878 63276 122884
rect 63130 120184 63186 120193
rect 63130 120119 63186 120128
rect 61936 103488 61988 103494
rect 61936 103430 61988 103436
rect 61752 86896 61804 86902
rect 61752 86838 61804 86844
rect 63236 82142 63264 122878
rect 63328 92410 63356 135895
rect 63420 114458 63448 263463
rect 64156 240825 64184 285602
rect 64512 282260 64564 282266
rect 64512 282202 64564 282208
rect 64142 240816 64198 240825
rect 64142 240751 64198 240760
rect 64524 240038 64552 282202
rect 64616 244934 64644 393314
rect 64800 252793 64828 404330
rect 65890 401568 65946 401577
rect 65890 401503 65946 401512
rect 65904 334121 65932 401503
rect 65996 389162 66024 474030
rect 66180 446418 66208 542982
rect 66626 540016 66682 540025
rect 66626 539951 66682 539960
rect 66640 539646 66668 539951
rect 66628 539640 66680 539646
rect 66628 539582 66680 539588
rect 66168 446412 66220 446418
rect 66168 446354 66220 446360
rect 66352 434036 66404 434042
rect 66352 433978 66404 433984
rect 66074 433936 66130 433945
rect 66074 433871 66130 433880
rect 65984 389156 66036 389162
rect 65984 389098 66036 389104
rect 65996 388482 66024 389098
rect 65984 388476 66036 388482
rect 65984 388418 66036 388424
rect 65890 334112 65946 334121
rect 65890 334047 65946 334056
rect 65984 301300 66036 301306
rect 65984 301242 66036 301248
rect 65890 294128 65946 294137
rect 65890 294063 65946 294072
rect 65904 274650 65932 294063
rect 65892 274644 65944 274650
rect 65892 274586 65944 274592
rect 64786 252784 64842 252793
rect 64786 252719 64842 252728
rect 64878 249928 64934 249937
rect 64708 249886 64878 249914
rect 64604 244928 64656 244934
rect 64604 244870 64656 244876
rect 64512 240032 64564 240038
rect 64512 239974 64564 239980
rect 63420 114442 63540 114458
rect 63420 114436 63552 114442
rect 63420 114430 63500 114436
rect 63500 114378 63552 114384
rect 64604 114436 64656 114442
rect 64604 114378 64656 114384
rect 64616 113257 64644 114378
rect 64602 113248 64658 113257
rect 64602 113183 64658 113192
rect 63408 99544 63460 99550
rect 63408 99486 63460 99492
rect 63316 92404 63368 92410
rect 63316 92346 63368 92352
rect 63224 82136 63276 82142
rect 63224 82078 63276 82084
rect 62028 80776 62080 80782
rect 62028 80718 62080 80724
rect 60740 45552 60792 45558
rect 60740 45494 60792 45500
rect 61936 8968 61988 8974
rect 61936 8910 61988 8916
rect 60832 3596 60884 3602
rect 60832 3538 60884 3544
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 58624 3188 58676 3194
rect 58624 3130 58676 3136
rect 59648 480 59676 3470
rect 60844 480 60872 3538
rect 61948 3482 61976 8910
rect 62040 3602 62068 80718
rect 63420 77246 63448 99486
rect 63408 77240 63460 77246
rect 63408 77182 63460 77188
rect 64616 40730 64644 113183
rect 64708 102134 64736 249886
rect 64878 249863 64934 249872
rect 64786 241632 64842 241641
rect 64786 241567 64842 241576
rect 64696 102128 64748 102134
rect 64696 102070 64748 102076
rect 64800 93838 64828 241567
rect 65996 240145 66024 301242
rect 66088 300898 66116 433871
rect 66364 433401 66392 433978
rect 66350 433392 66406 433401
rect 66350 433327 66406 433336
rect 66810 432576 66866 432585
rect 66810 432511 66866 432520
rect 66824 432002 66852 432511
rect 66812 431996 66864 432002
rect 66812 431938 66864 431944
rect 66810 431488 66866 431497
rect 66810 431423 66866 431432
rect 66824 430642 66852 431423
rect 66812 430636 66864 430642
rect 66812 430578 66864 430584
rect 66810 430400 66866 430409
rect 66810 430335 66866 430344
rect 66258 429312 66314 429321
rect 66258 429247 66260 429256
rect 66312 429247 66314 429256
rect 66260 429218 66312 429224
rect 66824 429214 66852 430335
rect 66812 429208 66864 429214
rect 66812 429150 66864 429156
rect 66166 428224 66222 428233
rect 66166 428159 66222 428168
rect 66076 300892 66128 300898
rect 66076 300834 66128 300840
rect 66088 279614 66116 300834
rect 66076 279608 66128 279614
rect 66076 279550 66128 279556
rect 66076 277364 66128 277370
rect 66076 277306 66128 277312
rect 65982 240136 66038 240145
rect 65982 240071 66038 240080
rect 66088 159390 66116 277306
rect 66180 271561 66208 428159
rect 66810 427408 66866 427417
rect 66810 427343 66866 427352
rect 66824 426494 66852 427343
rect 66812 426488 66864 426494
rect 66812 426430 66864 426436
rect 66536 425740 66588 425746
rect 66536 425682 66588 425688
rect 66548 425241 66576 425682
rect 66534 425232 66590 425241
rect 66534 425167 66590 425176
rect 66626 424144 66682 424153
rect 66626 424079 66682 424088
rect 66640 423706 66668 424079
rect 66628 423700 66680 423706
rect 66628 423642 66680 423648
rect 66812 423496 66864 423502
rect 66812 423438 66864 423444
rect 66824 423337 66852 423438
rect 66810 423328 66866 423337
rect 66810 423263 66866 423272
rect 66810 421152 66866 421161
rect 66810 421087 66866 421096
rect 66824 420986 66852 421087
rect 66812 420980 66864 420986
rect 66812 420922 66864 420928
rect 66810 420064 66866 420073
rect 66810 419999 66866 420008
rect 66824 419558 66852 419999
rect 66812 419552 66864 419558
rect 66812 419494 66864 419500
rect 66812 419416 66864 419422
rect 66812 419358 66864 419364
rect 66824 418266 66852 419358
rect 66812 418260 66864 418266
rect 66812 418202 66864 418208
rect 66824 417081 66852 418202
rect 66810 417072 66866 417081
rect 66810 417007 66866 417016
rect 66720 416764 66772 416770
rect 66720 416706 66772 416712
rect 66732 415993 66760 416706
rect 66718 415984 66774 415993
rect 66718 415919 66774 415928
rect 66718 414896 66774 414905
rect 66718 414831 66774 414840
rect 66732 414118 66760 414831
rect 66720 414112 66772 414118
rect 66720 414054 66772 414060
rect 66260 413296 66312 413302
rect 66260 413238 66312 413244
rect 66272 413001 66300 413238
rect 66258 412992 66314 413001
rect 66258 412927 66314 412936
rect 66810 410816 66866 410825
rect 66810 410751 66866 410760
rect 66824 409902 66852 410751
rect 66812 409896 66864 409902
rect 66812 409838 66864 409844
rect 66626 408912 66682 408921
rect 66626 408847 66682 408856
rect 66640 408542 66668 408847
rect 66628 408536 66680 408542
rect 66628 408478 66680 408484
rect 66810 407824 66866 407833
rect 66810 407759 66866 407768
rect 66824 407182 66852 407759
rect 66812 407176 66864 407182
rect 66812 407118 66864 407124
rect 66442 405648 66498 405657
rect 66442 405583 66498 405592
rect 66352 404320 66404 404326
rect 66352 404262 66404 404268
rect 66364 403102 66392 404262
rect 66352 403096 66404 403102
rect 66352 403038 66404 403044
rect 66364 402665 66392 403038
rect 66350 402656 66406 402665
rect 66350 402591 66406 402600
rect 66456 400926 66484 405583
rect 66810 404560 66866 404569
rect 66810 404495 66866 404504
rect 66824 404394 66852 404495
rect 66812 404388 66864 404394
rect 66812 404330 66864 404336
rect 66916 404326 66944 578575
rect 67546 577280 67602 577289
rect 67546 577215 67602 577224
rect 66994 570208 67050 570217
rect 66994 570143 67050 570152
rect 67008 419626 67036 570143
rect 67454 552256 67510 552265
rect 67454 552191 67510 552200
rect 67468 539918 67496 552191
rect 67456 539912 67508 539918
rect 67456 539854 67508 539860
rect 67088 436756 67140 436762
rect 67088 436698 67140 436704
rect 66996 419620 67048 419626
rect 66996 419562 67048 419568
rect 67100 419506 67128 436698
rect 67456 433288 67508 433294
rect 67454 433256 67456 433265
rect 67508 433256 67510 433265
rect 67454 433191 67510 433200
rect 67008 419478 67128 419506
rect 67008 418198 67036 419478
rect 66996 418192 67048 418198
rect 66994 418160 66996 418169
rect 67048 418160 67050 418169
rect 66994 418095 67050 418104
rect 67454 409728 67510 409737
rect 67454 409663 67510 409672
rect 66904 404320 66956 404326
rect 66904 404262 66956 404268
rect 66810 403744 66866 403753
rect 66810 403679 66866 403688
rect 66824 403034 66852 403679
rect 66812 403028 66864 403034
rect 66812 402970 66864 402976
rect 66444 400920 66496 400926
rect 66444 400862 66496 400868
rect 66810 400480 66866 400489
rect 66810 400415 66866 400424
rect 66824 400246 66852 400415
rect 66812 400240 66864 400246
rect 66812 400182 66864 400188
rect 66810 399664 66866 399673
rect 66810 399599 66866 399608
rect 66824 398886 66852 399599
rect 66812 398880 66864 398886
rect 66812 398822 66864 398828
rect 66810 398576 66866 398585
rect 66810 398511 66866 398520
rect 66824 396778 66852 398511
rect 66902 397488 66958 397497
rect 66902 397423 66958 397432
rect 66812 396772 66864 396778
rect 66812 396714 66864 396720
rect 66810 396400 66866 396409
rect 66810 396335 66866 396344
rect 66824 396166 66852 396335
rect 66812 396160 66864 396166
rect 66812 396102 66864 396108
rect 66812 395344 66864 395350
rect 66810 395312 66812 395321
rect 66864 395312 66866 395321
rect 66810 395247 66866 395256
rect 66810 394496 66866 394505
rect 66810 394431 66866 394440
rect 66824 393378 66852 394431
rect 66812 393372 66864 393378
rect 66812 393314 66864 393320
rect 66810 392320 66866 392329
rect 66810 392255 66866 392264
rect 66824 392018 66852 392255
rect 66812 392012 66864 392018
rect 66812 391954 66864 391960
rect 66810 391232 66866 391241
rect 66810 391167 66866 391176
rect 66824 387569 66852 391167
rect 66810 387560 66866 387569
rect 66810 387495 66866 387504
rect 66916 304978 66944 397423
rect 67468 342310 67496 409663
rect 67560 405657 67588 577215
rect 67652 566681 67680 703054
rect 67732 587172 67784 587178
rect 67732 587114 67784 587120
rect 67744 575385 67772 587114
rect 70228 582457 70256 703258
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 84108 703044 84160 703050
rect 84108 702986 84160 702992
rect 71688 700324 71740 700330
rect 71688 700266 71740 700272
rect 71700 587178 71728 700266
rect 71688 587172 71740 587178
rect 71688 587114 71740 587120
rect 71792 584905 71820 702986
rect 79968 702704 80020 702710
rect 79968 702646 80020 702652
rect 74540 656940 74592 656946
rect 74540 656882 74592 656888
rect 74552 596174 74580 656882
rect 74552 596146 74672 596174
rect 72422 585168 72478 585177
rect 72422 585103 72478 585112
rect 71778 584896 71834 584905
rect 71778 584831 71834 584840
rect 69478 582448 69534 582457
rect 70214 582448 70270 582457
rect 69478 582383 69534 582392
rect 69940 582412 69992 582418
rect 69492 580938 69520 582383
rect 70214 582383 70270 582392
rect 69940 582354 69992 582360
rect 69664 581120 69716 581126
rect 69664 581062 69716 581068
rect 69952 581074 69980 582354
rect 72436 581074 72464 585103
rect 73804 582480 73856 582486
rect 73804 582422 73856 582428
rect 73528 582412 73580 582418
rect 73528 582354 73580 582360
rect 73540 581074 73568 582354
rect 69032 580910 69520 580938
rect 69032 580802 69060 580910
rect 68664 580774 69060 580802
rect 68664 578921 68692 580774
rect 69676 580718 69704 581062
rect 69952 581046 70288 581074
rect 72128 581046 72464 581074
rect 73232 581046 73568 581074
rect 73816 581074 73844 582422
rect 74644 581074 74672 596146
rect 79980 588033 80008 702646
rect 84120 590714 84148 702986
rect 86224 702772 86276 702778
rect 86224 702714 86276 702720
rect 83464 590708 83516 590714
rect 83464 590650 83516 590656
rect 84108 590708 84160 590714
rect 84108 590650 84160 590656
rect 79966 588024 80022 588033
rect 79966 587959 80022 587968
rect 78128 585812 78180 585818
rect 78128 585754 78180 585760
rect 76288 583840 76340 583846
rect 76288 583782 76340 583788
rect 75366 581088 75422 581097
rect 73816 581046 74152 581074
rect 74644 581046 75366 581074
rect 76300 581074 76328 583782
rect 77208 583160 77260 583166
rect 77208 583102 77260 583108
rect 77220 581074 77248 583102
rect 78140 581097 78168 585754
rect 79324 585200 79376 585206
rect 79324 585142 79376 585148
rect 79046 582720 79102 582729
rect 79046 582655 79102 582664
rect 78126 581088 78182 581097
rect 75992 581046 76328 581074
rect 76912 581046 77248 581074
rect 77832 581046 78126 581074
rect 75366 581023 75422 581032
rect 79060 581074 79088 582655
rect 78752 581046 79088 581074
rect 79336 581074 79364 585142
rect 79980 583166 80008 587959
rect 82726 583808 82782 583817
rect 82726 583743 82782 583752
rect 79968 583160 80020 583166
rect 79968 583102 80020 583108
rect 81808 582616 81860 582622
rect 81808 582558 81860 582564
rect 80244 581120 80296 581126
rect 79336 581046 79672 581074
rect 81820 581074 81848 582558
rect 82740 581074 82768 583743
rect 83476 582622 83504 590650
rect 86236 586514 86264 702714
rect 89180 702434 89208 703520
rect 89720 703248 89772 703254
rect 89720 703190 89772 703196
rect 86144 586486 86264 586514
rect 88352 702406 89208 702434
rect 83464 582616 83516 582622
rect 83464 582558 83516 582564
rect 83002 581224 83058 581233
rect 83002 581159 83058 581168
rect 80296 581068 80592 581074
rect 80244 581062 80592 581068
rect 80256 581046 80592 581062
rect 81512 581046 81848 581074
rect 82432 581046 82768 581074
rect 83016 581074 83044 581159
rect 83016 581046 83352 581074
rect 78126 581023 78182 581032
rect 78140 580963 78168 581023
rect 70950 580816 71006 580825
rect 84198 580816 84254 580825
rect 71006 580774 71208 580802
rect 70950 580751 71006 580760
rect 86144 580802 86172 586486
rect 88352 585818 88380 702406
rect 89732 596174 89760 703190
rect 101496 702976 101548 702982
rect 101496 702918 101548 702924
rect 99288 702772 99340 702778
rect 99288 702714 99340 702720
rect 96620 702636 96672 702642
rect 96620 702578 96672 702584
rect 94780 605872 94832 605878
rect 94780 605814 94832 605820
rect 89732 596146 89852 596174
rect 88340 585812 88392 585818
rect 88340 585754 88392 585760
rect 87512 585200 87564 585206
rect 87512 585142 87564 585148
rect 86592 581120 86644 581126
rect 87524 581074 87552 585142
rect 89718 582720 89774 582729
rect 89718 582655 89774 582664
rect 88246 582584 88302 582593
rect 88246 582519 88302 582528
rect 88260 581074 88288 582519
rect 89732 581641 89760 582655
rect 89718 581632 89774 581641
rect 89718 581567 89774 581576
rect 86592 581062 86644 581068
rect 86604 580802 86632 581062
rect 87216 581046 87552 581074
rect 88136 581046 88288 581074
rect 89824 581058 89852 596146
rect 92480 583772 92532 583778
rect 92480 583714 92532 583720
rect 90272 582480 90324 582486
rect 90272 582422 90324 582428
rect 92110 582448 92166 582457
rect 90284 581074 90312 582422
rect 92110 582383 92166 582392
rect 92124 581074 92152 582383
rect 89812 581052 89864 581058
rect 89976 581046 90312 581074
rect 90560 581058 90896 581074
rect 90548 581052 90896 581058
rect 89812 580994 89864 581000
rect 90600 581046 90896 581052
rect 91816 581046 92152 581074
rect 92492 581074 92520 583714
rect 92492 581046 92736 581074
rect 93656 581058 93808 581074
rect 93656 581052 93820 581058
rect 93656 581046 93768 581052
rect 90548 580994 90600 581000
rect 93768 580994 93820 581000
rect 84254 580774 84456 580802
rect 85376 580774 85528 580802
rect 86144 580774 86632 580802
rect 88706 580816 88762 580825
rect 84198 580751 84254 580760
rect 85500 580718 85528 580774
rect 88762 580774 89056 580802
rect 88706 580751 88762 580760
rect 69664 580712 69716 580718
rect 69664 580654 69716 580660
rect 85488 580712 85540 580718
rect 85488 580654 85540 580660
rect 94576 580366 94728 580394
rect 68650 578912 68706 578921
rect 68650 578847 68706 578856
rect 67730 575376 67786 575385
rect 67730 575311 67786 575320
rect 67730 568848 67786 568857
rect 67730 568783 67786 568792
rect 67638 566672 67694 566681
rect 67638 566607 67694 566616
rect 67652 565894 67680 566607
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67638 556608 67694 556617
rect 67638 556543 67694 556552
rect 67652 445194 67680 556543
rect 67744 474026 67772 568783
rect 67822 550896 67878 550905
rect 67822 550831 67878 550840
rect 67732 474020 67784 474026
rect 67732 473962 67784 473968
rect 67732 469872 67784 469878
rect 67732 469814 67784 469820
rect 67640 445188 67692 445194
rect 67640 445130 67692 445136
rect 67744 414089 67772 469814
rect 67836 464370 67864 550831
rect 71780 539912 71832 539918
rect 69110 539880 69166 539889
rect 71780 539854 71832 539860
rect 93858 539880 93914 539889
rect 69110 539815 69166 539824
rect 68816 539158 68968 539186
rect 68940 533390 68968 539158
rect 68928 533384 68980 533390
rect 68928 533326 68980 533332
rect 67824 464364 67876 464370
rect 67824 464306 67876 464312
rect 68468 451920 68520 451926
rect 68468 451862 68520 451868
rect 68480 436257 68508 451862
rect 68466 436248 68522 436257
rect 68466 436183 68522 436192
rect 68480 434330 68508 436183
rect 69124 435266 69152 539815
rect 69400 539158 69736 539186
rect 70656 539158 70992 539186
rect 69400 536110 69428 539158
rect 70964 538286 70992 539158
rect 71240 539158 71576 539186
rect 70952 538280 71004 538286
rect 70952 538222 71004 538228
rect 70964 537606 70992 538222
rect 70952 537600 71004 537606
rect 70952 537542 71004 537548
rect 69388 536104 69440 536110
rect 69388 536046 69440 536052
rect 71240 528554 71268 539158
rect 70504 528526 71268 528554
rect 70504 444786 70532 528526
rect 70492 444780 70544 444786
rect 70492 444722 70544 444728
rect 71136 437436 71188 437442
rect 71136 437378 71188 437384
rect 71148 436150 71176 437378
rect 71136 436144 71188 436150
rect 71136 436086 71188 436092
rect 69112 435260 69164 435266
rect 69112 435202 69164 435208
rect 69940 435260 69992 435266
rect 69940 435202 69992 435208
rect 69124 434858 69152 435202
rect 69112 434852 69164 434858
rect 69112 434794 69164 434800
rect 69952 434330 69980 435202
rect 68480 434302 68816 434330
rect 69952 434302 70288 434330
rect 68652 434240 68704 434246
rect 71148 434194 71176 436086
rect 71792 434586 71820 539854
rect 87604 539844 87656 539850
rect 93858 539815 93860 539824
rect 87604 539786 87656 539792
rect 93912 539815 93914 539824
rect 93860 539786 93912 539792
rect 71884 539158 72496 539186
rect 73416 539158 73476 539186
rect 74336 539158 74488 539186
rect 71884 450566 71912 539158
rect 73448 536790 73476 539158
rect 73436 536784 73488 536790
rect 73436 536726 73488 536732
rect 74460 471306 74488 539158
rect 74644 539158 75256 539186
rect 76176 539158 76512 539186
rect 74448 471300 74500 471306
rect 74448 471242 74500 471248
rect 71872 450560 71924 450566
rect 71872 450502 71924 450508
rect 74644 436762 74672 539158
rect 75184 538892 75236 538898
rect 75184 538834 75236 538840
rect 74724 439544 74776 439550
rect 74724 439486 74776 439492
rect 74632 436756 74684 436762
rect 74632 436698 74684 436704
rect 71780 434580 71832 434586
rect 71780 434522 71832 434528
rect 73022 434580 73074 434586
rect 73022 434522 73074 434528
rect 71792 434246 71820 434522
rect 73034 434316 73062 434522
rect 74736 434353 74764 439486
rect 75196 437442 75224 538834
rect 76484 536761 76512 539158
rect 76760 539158 77096 539186
rect 78016 539158 78352 539186
rect 76564 536784 76616 536790
rect 76470 536752 76526 536761
rect 76564 536726 76616 536732
rect 76470 536687 76526 536696
rect 76484 535673 76512 536687
rect 76470 535664 76526 535673
rect 76470 535599 76526 535608
rect 75918 535528 75974 535537
rect 75918 535463 75974 535472
rect 75932 474094 75960 535463
rect 76576 519586 76604 536726
rect 76760 535537 76788 539158
rect 78324 536654 78352 539158
rect 78692 539158 78936 539186
rect 80040 539158 80192 539186
rect 78312 536648 78364 536654
rect 78312 536590 78364 536596
rect 77206 535664 77262 535673
rect 77206 535599 77262 535608
rect 76746 535528 76802 535537
rect 76746 535463 76802 535472
rect 76564 519580 76616 519586
rect 76564 519522 76616 519528
rect 75920 474088 75972 474094
rect 75920 474030 75972 474036
rect 77116 467152 77168 467158
rect 77116 467094 77168 467100
rect 77128 441614 77156 467094
rect 77220 459746 77248 535599
rect 78692 465730 78720 539158
rect 79324 537600 79376 537606
rect 79324 537542 79376 537548
rect 78680 465724 78732 465730
rect 78680 465666 78732 465672
rect 77208 459740 77260 459746
rect 77208 459682 77260 459688
rect 77944 459740 77996 459746
rect 77944 459682 77996 459688
rect 76944 441586 77156 441614
rect 75184 437436 75236 437442
rect 75184 437378 75236 437384
rect 75458 434480 75514 434489
rect 75458 434415 75514 434424
rect 74722 434344 74778 434353
rect 75472 434330 75500 434415
rect 76194 434344 76250 434353
rect 74778 434302 75072 434330
rect 75472 434302 75808 434330
rect 74722 434279 74778 434288
rect 76944 434330 76972 441586
rect 77392 436484 77444 436490
rect 77392 436426 77444 436432
rect 77404 436257 77432 436426
rect 77390 436248 77446 436257
rect 77390 436183 77446 436192
rect 77404 434330 77432 436183
rect 77482 435432 77538 435441
rect 77482 435367 77538 435376
rect 76250 434302 76972 434330
rect 77280 434302 77432 434330
rect 77496 434330 77524 435367
rect 77956 434761 77984 459682
rect 79336 457502 79364 537542
rect 80164 535838 80192 539158
rect 80256 539158 80960 539186
rect 81880 539158 82124 539186
rect 82800 539158 82860 539186
rect 80152 535832 80204 535838
rect 80152 535774 80204 535780
rect 80256 528554 80284 539158
rect 81348 535832 81400 535838
rect 81348 535774 81400 535780
rect 80072 528526 80284 528554
rect 79324 457496 79376 457502
rect 79324 457438 79376 457444
rect 80072 453257 80100 528526
rect 81360 520985 81388 535774
rect 82096 535498 82124 539158
rect 82176 536648 82228 536654
rect 82176 536590 82228 536596
rect 82084 535492 82136 535498
rect 82084 535434 82136 535440
rect 82084 530664 82136 530670
rect 82084 530606 82136 530612
rect 81346 520976 81402 520985
rect 81346 520911 81402 520920
rect 80058 453248 80114 453257
rect 80058 453183 80114 453192
rect 80336 446412 80388 446418
rect 80336 446354 80388 446360
rect 77942 434752 77998 434761
rect 77942 434687 77998 434696
rect 80242 434344 80298 434353
rect 77496 434302 77832 434330
rect 80040 434302 80242 434330
rect 76194 434279 76250 434288
rect 80348 434330 80376 446354
rect 81346 444952 81402 444961
rect 81346 444887 81402 444896
rect 80426 434888 80482 434897
rect 80426 434823 80482 434832
rect 80298 434302 80376 434330
rect 80440 434330 80468 434823
rect 81360 434602 81388 444887
rect 81624 443692 81676 443698
rect 81624 443634 81676 443640
rect 81314 434574 81388 434602
rect 80978 434344 81034 434353
rect 80440 434302 80592 434330
rect 80242 434279 80298 434288
rect 81314 434330 81342 434574
rect 81034 434316 81342 434330
rect 81636 434330 81664 443634
rect 82096 436490 82124 530606
rect 82188 482322 82216 536590
rect 82176 482316 82228 482322
rect 82176 482258 82228 482264
rect 82832 445058 82860 539158
rect 82924 539158 83720 539186
rect 84212 539158 84640 539186
rect 85560 539158 85620 539186
rect 86480 539158 86724 539186
rect 82924 487830 82952 539158
rect 83464 525088 83516 525094
rect 83464 525030 83516 525036
rect 82912 487824 82964 487830
rect 82912 487766 82964 487772
rect 83096 445188 83148 445194
rect 83096 445130 83148 445136
rect 82820 445052 82872 445058
rect 82820 444994 82872 445000
rect 83108 441614 83136 445130
rect 83476 443601 83504 525030
rect 84212 476814 84240 539158
rect 84200 476808 84252 476814
rect 84200 476750 84252 476756
rect 85592 468518 85620 539158
rect 86696 536110 86724 539158
rect 86972 539158 87400 539186
rect 86684 536104 86736 536110
rect 86684 536046 86736 536052
rect 86224 535492 86276 535498
rect 86224 535434 86276 535440
rect 85580 468512 85632 468518
rect 85580 468454 85632 468460
rect 85672 449200 85724 449206
rect 86236 449177 86264 535434
rect 86868 478168 86920 478174
rect 86868 478110 86920 478116
rect 85672 449142 85724 449148
rect 86222 449168 86278 449177
rect 83462 443592 83518 443601
rect 83462 443527 83518 443536
rect 85684 441614 85712 449142
rect 86222 449103 86278 449112
rect 83108 441586 83228 441614
rect 85684 441586 85896 441614
rect 82084 436484 82136 436490
rect 82084 436426 82136 436432
rect 83200 436121 83228 441586
rect 83740 438184 83792 438190
rect 83740 438126 83792 438132
rect 83186 436112 83242 436121
rect 83186 436047 83242 436056
rect 82910 434752 82966 434761
rect 82910 434687 82966 434696
rect 81898 434344 81954 434353
rect 81034 434302 81328 434316
rect 81636 434302 81898 434330
rect 80978 434279 81034 434288
rect 81954 434302 82064 434330
rect 81898 434279 81954 434288
rect 68652 434182 68704 434188
rect 68284 433696 68336 433702
rect 68284 433638 68336 433644
rect 67730 414080 67786 414089
rect 67730 414015 67732 414024
rect 67784 414015 67786 414024
rect 67732 413986 67784 413992
rect 67744 413955 67772 413986
rect 67546 405648 67602 405657
rect 67546 405583 67602 405592
rect 67640 390176 67692 390182
rect 67640 390118 67692 390124
rect 66996 342304 67048 342310
rect 66996 342246 67048 342252
rect 67456 342304 67508 342310
rect 67456 342246 67508 342252
rect 67008 330546 67036 342246
rect 66996 330540 67048 330546
rect 66996 330482 67048 330488
rect 67548 327752 67600 327758
rect 67548 327694 67600 327700
rect 67560 326369 67588 327694
rect 67546 326360 67602 326369
rect 67546 326295 67602 326304
rect 66904 304972 66956 304978
rect 66904 304914 66956 304920
rect 67548 284980 67600 284986
rect 67548 284922 67600 284928
rect 67560 281353 67588 284922
rect 67546 281344 67602 281353
rect 67546 281279 67602 281288
rect 67560 280226 67588 281279
rect 67548 280220 67600 280226
rect 67548 280162 67600 280168
rect 66626 279712 66682 279721
rect 66626 279647 66682 279656
rect 66640 279614 66668 279647
rect 66628 279608 66680 279614
rect 66628 279550 66680 279556
rect 66812 279472 66864 279478
rect 66812 279414 66864 279420
rect 66824 278905 66852 279414
rect 66810 278896 66866 278905
rect 66810 278831 66866 278840
rect 66810 278080 66866 278089
rect 66810 278015 66812 278024
rect 66864 278015 66866 278024
rect 66812 277986 66864 277992
rect 66810 276448 66866 276457
rect 66810 276383 66866 276392
rect 66824 276078 66852 276383
rect 66812 276072 66864 276078
rect 66812 276014 66864 276020
rect 66904 276004 66956 276010
rect 66904 275946 66956 275952
rect 66916 275641 66944 275946
rect 66902 275632 66958 275641
rect 66902 275567 66958 275576
rect 66536 274644 66588 274650
rect 66536 274586 66588 274592
rect 66548 274009 66576 274586
rect 66534 274000 66590 274009
rect 66534 273935 66590 273944
rect 66258 273184 66314 273193
rect 66258 273119 66314 273128
rect 66272 271969 66300 273119
rect 66810 272368 66866 272377
rect 66810 272303 66866 272312
rect 66824 272134 66852 272303
rect 66812 272128 66864 272134
rect 66812 272070 66864 272076
rect 66258 271960 66314 271969
rect 66258 271895 66314 271904
rect 66812 271856 66864 271862
rect 66812 271798 66864 271804
rect 66166 271552 66222 271561
rect 66166 271487 66222 271496
rect 66180 270745 66208 271487
rect 66824 270745 66852 271798
rect 66166 270736 66222 270745
rect 66166 270671 66222 270680
rect 66810 270736 66866 270745
rect 66810 270671 66866 270680
rect 66168 268388 66220 268394
rect 66168 268330 66220 268336
rect 66180 268297 66208 268330
rect 66166 268288 66222 268297
rect 66166 268223 66222 268232
rect 66076 159384 66128 159390
rect 66076 159326 66128 159332
rect 65982 129024 66038 129033
rect 65982 128959 66038 128968
rect 65522 123856 65578 123865
rect 65522 123791 65578 123800
rect 65536 121446 65564 123791
rect 65524 121440 65576 121446
rect 65524 121382 65576 121388
rect 64788 93832 64840 93838
rect 64788 93774 64840 93780
rect 65536 66910 65564 121382
rect 65616 96688 65668 96694
rect 65616 96630 65668 96636
rect 65628 86970 65656 96630
rect 65616 86964 65668 86970
rect 65616 86906 65668 86912
rect 65524 66904 65576 66910
rect 65524 66846 65576 66852
rect 64604 40724 64656 40730
rect 64604 40666 64656 40672
rect 65996 17270 66024 128959
rect 66088 126041 66116 159326
rect 66180 145625 66208 268223
rect 66260 267708 66312 267714
rect 66260 267650 66312 267656
rect 66272 266529 66300 267650
rect 66810 267472 66866 267481
rect 66810 267407 66866 267416
rect 66258 266520 66314 266529
rect 66258 266455 66314 266464
rect 66824 266422 66852 267407
rect 66812 266416 66864 266422
rect 66812 266358 66864 266364
rect 66812 265192 66864 265198
rect 66812 265134 66864 265140
rect 66824 265033 66852 265134
rect 66810 265024 66866 265033
rect 66810 264959 66866 264968
rect 66628 264240 66680 264246
rect 66628 264182 66680 264188
rect 66640 263401 66668 264182
rect 66626 263392 66682 263401
rect 66626 263327 66682 263336
rect 66904 262880 66956 262886
rect 66904 262822 66956 262828
rect 66916 262585 66944 262822
rect 66902 262576 66958 262585
rect 66902 262511 66958 262520
rect 66720 261520 66772 261526
rect 66720 261462 66772 261468
rect 66732 260953 66760 261462
rect 66718 260944 66774 260953
rect 66718 260879 66774 260888
rect 66444 260840 66496 260846
rect 66444 260782 66496 260788
rect 66456 260137 66484 260782
rect 66442 260128 66498 260137
rect 66442 260063 66498 260072
rect 66260 258188 66312 258194
rect 66260 258130 66312 258136
rect 66272 258058 66300 258130
rect 66352 258120 66404 258126
rect 66352 258062 66404 258068
rect 66260 258052 66312 258058
rect 66260 257994 66312 258000
rect 66364 256873 66392 258062
rect 66626 257680 66682 257689
rect 66626 257615 66682 257624
rect 66640 257378 66668 257615
rect 66628 257372 66680 257378
rect 66628 257314 66680 257320
rect 66350 256864 66406 256873
rect 66350 256799 66406 256808
rect 66812 256692 66864 256698
rect 66812 256634 66864 256640
rect 66824 256057 66852 256634
rect 66810 256048 66866 256057
rect 66810 255983 66866 255992
rect 66810 255232 66866 255241
rect 66810 255167 66866 255176
rect 66824 253978 66852 255167
rect 66812 253972 66864 253978
rect 66812 253914 66864 253920
rect 66994 253600 67050 253609
rect 66994 253535 67050 253544
rect 67008 253230 67036 253535
rect 66996 253224 67048 253230
rect 66996 253166 67048 253172
rect 67364 253224 67416 253230
rect 67364 253166 67416 253172
rect 66812 251252 66864 251258
rect 66812 251194 66864 251200
rect 66824 251161 66852 251194
rect 66810 251152 66866 251161
rect 66810 251087 66866 251096
rect 66720 250504 66772 250510
rect 66720 250446 66772 250452
rect 66732 249529 66760 250446
rect 66718 249520 66774 249529
rect 66718 249455 66774 249464
rect 66994 246256 67050 246265
rect 66994 246191 67050 246200
rect 67008 246158 67036 246191
rect 66996 246152 67048 246158
rect 66996 246094 67048 246100
rect 67272 246152 67324 246158
rect 67272 246094 67324 246100
rect 66904 244928 66956 244934
rect 66904 244870 66956 244876
rect 66916 244633 66944 244870
rect 66902 244624 66958 244633
rect 66902 244559 66958 244568
rect 66810 243808 66866 243817
rect 66810 243743 66866 243752
rect 66824 242962 66852 243743
rect 66812 242956 66864 242962
rect 66812 242898 66864 242904
rect 67284 213858 67312 246094
rect 67376 235958 67404 253166
rect 67468 247110 67496 247141
rect 67456 247104 67508 247110
rect 67454 247072 67456 247081
rect 67508 247072 67510 247081
rect 67454 247007 67510 247016
rect 67364 235952 67416 235958
rect 67364 235894 67416 235900
rect 66812 213852 66864 213858
rect 66812 213794 66864 213800
rect 67272 213852 67324 213858
rect 67272 213794 67324 213800
rect 66166 145616 66222 145625
rect 66166 145551 66222 145560
rect 66074 126032 66130 126041
rect 66074 125967 66130 125976
rect 66074 119232 66130 119241
rect 66074 119167 66130 119176
rect 66088 84862 66116 119167
rect 66180 117609 66208 145551
rect 66260 135244 66312 135250
rect 66260 135186 66312 135192
rect 66272 134473 66300 135186
rect 66258 134464 66314 134473
rect 66258 134399 66314 134408
rect 66260 133884 66312 133890
rect 66260 133826 66312 133832
rect 66272 133657 66300 133826
rect 66258 133648 66314 133657
rect 66258 133583 66314 133592
rect 66260 132456 66312 132462
rect 66260 132398 66312 132404
rect 66272 132025 66300 132398
rect 66352 132388 66404 132394
rect 66352 132330 66404 132336
rect 66258 132016 66314 132025
rect 66258 131951 66314 131960
rect 66364 131209 66392 132330
rect 66350 131200 66406 131209
rect 66350 131135 66406 131144
rect 66444 129056 66496 129062
rect 66444 128998 66496 129004
rect 66456 128217 66484 128998
rect 66720 128240 66772 128246
rect 66442 128208 66498 128217
rect 66720 128182 66772 128188
rect 66442 128143 66498 128152
rect 66732 126857 66760 128182
rect 66718 126848 66774 126857
rect 66718 126783 66774 126792
rect 66260 125588 66312 125594
rect 66260 125530 66312 125536
rect 66272 124409 66300 125530
rect 66258 124400 66314 124409
rect 66258 124335 66314 124344
rect 66720 122732 66772 122738
rect 66720 122674 66772 122680
rect 66732 120601 66760 122674
rect 66718 120592 66774 120601
rect 66718 120527 66774 120536
rect 66260 120216 66312 120222
rect 66260 120158 66312 120164
rect 66272 119241 66300 120158
rect 66258 119232 66314 119241
rect 66258 119167 66314 119176
rect 66166 117600 66222 117609
rect 66166 117535 66222 117544
rect 66628 114504 66680 114510
rect 66628 114446 66680 114452
rect 66640 113257 66668 114446
rect 66626 113248 66682 113257
rect 66626 113183 66682 113192
rect 66258 110256 66314 110265
rect 66258 110191 66314 110200
rect 66272 109070 66300 110191
rect 66260 109064 66312 109070
rect 66260 109006 66312 109012
rect 66720 107568 66772 107574
rect 66720 107510 66772 107516
rect 66732 106457 66760 107510
rect 66718 106448 66774 106457
rect 66718 106383 66774 106392
rect 66260 104848 66312 104854
rect 66258 104816 66260 104825
rect 66312 104816 66314 104825
rect 66258 104751 66314 104760
rect 66444 102128 66496 102134
rect 66444 102070 66496 102076
rect 66456 101017 66484 102070
rect 66824 101946 66852 213794
rect 66904 128308 66956 128314
rect 66904 128250 66956 128256
rect 66916 127673 66944 128250
rect 66902 127664 66958 127673
rect 66902 127599 66958 127608
rect 66904 126268 66956 126274
rect 66904 126210 66956 126216
rect 66916 125225 66944 126210
rect 66902 125216 66958 125225
rect 66902 125151 66958 125160
rect 66902 123040 66958 123049
rect 66902 122975 66958 122984
rect 66916 122942 66944 122975
rect 66904 122936 66956 122942
rect 66904 122878 66956 122884
rect 66904 122800 66956 122806
rect 66904 122742 66956 122748
rect 66916 122233 66944 122742
rect 66902 122224 66958 122233
rect 66902 122159 66958 122168
rect 66904 120080 66956 120086
rect 66902 120048 66904 120057
rect 66956 120048 66958 120057
rect 66902 119983 66958 119992
rect 66904 118584 66956 118590
rect 66904 118526 66956 118532
rect 66916 118425 66944 118526
rect 66902 118416 66958 118425
rect 66902 118351 66958 118360
rect 66904 117292 66956 117298
rect 66904 117234 66956 117240
rect 66916 117065 66944 117234
rect 66902 117056 66958 117065
rect 66902 116991 66958 117000
rect 66904 115932 66956 115938
rect 66904 115874 66956 115880
rect 66916 115433 66944 115874
rect 66902 115424 66958 115433
rect 66902 115359 66958 115368
rect 67192 114646 67220 114677
rect 67180 114640 67232 114646
rect 67178 114608 67180 114617
rect 67232 114608 67234 114617
rect 67178 114543 67234 114552
rect 66904 113144 66956 113150
rect 66904 113086 66956 113092
rect 66916 112441 66944 113086
rect 66902 112432 66958 112441
rect 66902 112367 66958 112376
rect 66904 111784 66956 111790
rect 66904 111726 66956 111732
rect 66916 110809 66944 111726
rect 66902 110800 66958 110809
rect 66902 110735 66958 110744
rect 66904 110424 66956 110430
rect 66904 110366 66956 110372
rect 66916 109449 66944 110366
rect 66902 109440 66958 109449
rect 66902 109375 66958 109384
rect 66996 108996 67048 109002
rect 66996 108938 67048 108944
rect 66904 108928 66956 108934
rect 66904 108870 66956 108876
rect 66916 108633 66944 108870
rect 66902 108624 66958 108633
rect 66902 108559 66958 108568
rect 67008 107817 67036 108938
rect 66994 107808 67050 107817
rect 66994 107743 67050 107752
rect 66904 107636 66956 107642
rect 66904 107578 66956 107584
rect 66916 107001 66944 107578
rect 66902 106992 66958 107001
rect 66902 106927 66958 106936
rect 66904 106276 66956 106282
rect 66904 106218 66956 106224
rect 66916 105641 66944 106218
rect 66902 105632 66958 105641
rect 66902 105567 66958 105576
rect 66904 103488 66956 103494
rect 66904 103430 66956 103436
rect 66916 103193 66944 103430
rect 66902 103184 66958 103193
rect 66902 103119 66958 103128
rect 66824 101918 66944 101946
rect 66810 101824 66866 101833
rect 66810 101759 66866 101768
rect 66824 101454 66852 101759
rect 66812 101448 66864 101454
rect 66812 101390 66864 101396
rect 66442 101008 66498 101017
rect 66442 100943 66498 100952
rect 66812 100700 66864 100706
rect 66812 100642 66864 100648
rect 66824 100201 66852 100642
rect 66810 100192 66866 100201
rect 66810 100127 66866 100136
rect 66810 99648 66866 99657
rect 66810 99583 66866 99592
rect 66824 99550 66852 99583
rect 66812 99544 66864 99550
rect 66812 99486 66864 99492
rect 66812 99340 66864 99346
rect 66812 99282 66864 99288
rect 66824 98841 66852 99282
rect 66810 98832 66866 98841
rect 66810 98767 66866 98776
rect 66812 97300 66864 97306
rect 66812 97242 66864 97248
rect 66260 96620 66312 96626
rect 66260 96562 66312 96568
rect 66272 96393 66300 96562
rect 66258 96384 66314 96393
rect 66258 96319 66314 96328
rect 66824 95849 66852 97242
rect 66916 97209 66944 101918
rect 66902 97200 66958 97209
rect 66902 97135 66958 97144
rect 66810 95840 66866 95849
rect 66810 95775 66866 95784
rect 66444 95192 66496 95198
rect 66444 95134 66496 95140
rect 66456 95033 66484 95134
rect 66442 95024 66498 95033
rect 66442 94959 66498 94968
rect 66812 93832 66864 93838
rect 66812 93774 66864 93780
rect 66824 93401 66852 93774
rect 66810 93392 66866 93401
rect 66810 93327 66866 93336
rect 66076 84856 66128 84862
rect 66076 84798 66128 84804
rect 67192 79354 67220 114543
rect 67376 104009 67404 235894
rect 67362 104000 67418 104009
rect 67362 103935 67418 103944
rect 67468 98025 67496 247007
rect 67560 129849 67588 280162
rect 67652 241369 67680 390118
rect 68296 277409 68324 433638
rect 68664 284986 68692 434182
rect 71024 434166 71176 434194
rect 71780 434240 71832 434246
rect 74736 434219 74764 434279
rect 80256 434219 80284 434279
rect 81912 434219 81940 434279
rect 82924 434194 82952 434687
rect 83200 434330 83228 436047
rect 83752 434489 83780 438126
rect 85762 437608 85818 437617
rect 85762 437543 85818 437552
rect 85120 436620 85172 436626
rect 85120 436562 85172 436568
rect 84474 434616 84530 434625
rect 84474 434551 84530 434560
rect 83738 434480 83794 434489
rect 83738 434415 83794 434424
rect 83752 434330 83780 434415
rect 84488 434330 84516 434551
rect 85132 434330 85160 436562
rect 85776 434330 85804 437543
rect 85868 434353 85896 441586
rect 86880 437617 86908 478110
rect 86972 456074 87000 539158
rect 86960 456068 87012 456074
rect 86960 456010 87012 456016
rect 86866 437608 86922 437617
rect 86866 437543 86922 437552
rect 87616 436626 87644 539786
rect 88320 539158 88472 539186
rect 88340 530188 88392 530194
rect 88340 530130 88392 530136
rect 88248 522300 88300 522306
rect 88248 522242 88300 522248
rect 87604 436620 87656 436626
rect 87604 436562 87656 436568
rect 88260 436121 88288 522242
rect 88352 441017 88380 530130
rect 88444 463049 88472 539158
rect 88904 539158 89240 539186
rect 90160 539158 90220 539186
rect 88904 530194 88932 539158
rect 90192 538286 90220 539158
rect 91204 539158 91264 539186
rect 91848 539158 92184 539186
rect 92492 539158 93104 539186
rect 94024 539158 94544 539186
rect 89720 538280 89772 538286
rect 89720 538222 89772 538228
rect 90180 538280 90232 538286
rect 90180 538222 90232 538228
rect 88892 530188 88944 530194
rect 88892 530130 88944 530136
rect 89732 467158 89760 538222
rect 91008 536104 91060 536110
rect 91008 536046 91060 536052
rect 90364 535492 90416 535498
rect 90364 535434 90416 535440
rect 89720 467152 89772 467158
rect 89720 467094 89772 467100
rect 88430 463040 88486 463049
rect 88430 462975 88486 462984
rect 90376 451926 90404 535434
rect 90454 468480 90510 468489
rect 90454 468415 90510 468424
rect 90364 451920 90416 451926
rect 90364 451862 90416 451868
rect 88338 441008 88394 441017
rect 88338 440943 88394 440952
rect 88708 440904 88760 440910
rect 88708 440846 88760 440852
rect 87326 436112 87382 436121
rect 87326 436047 87382 436056
rect 88246 436112 88302 436121
rect 88246 436047 88302 436056
rect 83200 434302 83536 434330
rect 83752 434302 84088 434330
rect 84488 434302 85160 434330
rect 85560 434302 85804 434330
rect 85854 434344 85910 434353
rect 87142 434344 87198 434353
rect 85910 434302 86296 434330
rect 87032 434302 87142 434330
rect 85854 434279 85910 434288
rect 87340 434330 87368 436047
rect 87198 434302 87368 434330
rect 88720 434330 88748 440846
rect 90088 438932 90140 438938
rect 90088 438874 90140 438880
rect 90100 434330 90128 438874
rect 90468 437442 90496 468415
rect 91020 438190 91048 536046
rect 91204 530670 91232 539158
rect 91848 535498 91876 539158
rect 91836 535492 91888 535498
rect 91836 535434 91888 535440
rect 91192 530664 91244 530670
rect 91192 530606 91244 530612
rect 92492 461650 92520 539158
rect 94516 534138 94544 539158
rect 94700 538257 94728 580366
rect 94792 579630 94820 605814
rect 95884 582480 95936 582486
rect 95884 582422 95936 582428
rect 94780 579624 94832 579630
rect 94780 579566 94832 579572
rect 95330 575376 95386 575385
rect 95330 575311 95386 575320
rect 95238 563680 95294 563689
rect 95238 563615 95294 563624
rect 94778 555520 94834 555529
rect 94778 555455 94834 555464
rect 94686 538248 94742 538257
rect 94686 538183 94742 538192
rect 94504 534132 94556 534138
rect 94504 534074 94556 534080
rect 92572 479528 92624 479534
rect 92572 479470 92624 479476
rect 92480 461644 92532 461650
rect 92480 461586 92532 461592
rect 92584 441614 92612 479470
rect 94516 452606 94544 534074
rect 94792 518129 94820 555455
rect 95148 540932 95200 540938
rect 95148 540874 95200 540880
rect 94778 518120 94834 518129
rect 94778 518055 94834 518064
rect 94504 452600 94556 452606
rect 94504 452542 94556 452548
rect 92584 441586 92704 441614
rect 91008 438184 91060 438190
rect 91008 438126 91060 438132
rect 90456 437436 90508 437442
rect 90456 437378 90508 437384
rect 91098 436248 91154 436257
rect 91098 436183 91154 436192
rect 91112 434602 91140 436183
rect 92676 434761 92704 441586
rect 95160 440298 95188 540874
rect 95252 454753 95280 563615
rect 95344 478174 95372 575311
rect 95896 567866 95924 582422
rect 95884 567860 95936 567866
rect 95884 567802 95936 567808
rect 95422 567216 95478 567225
rect 95422 567151 95478 567160
rect 95436 527785 95464 567151
rect 96632 552537 96660 702578
rect 96712 589960 96764 589966
rect 96712 589902 96764 589908
rect 96724 558793 96752 589902
rect 96804 579624 96856 579630
rect 96804 579566 96856 579572
rect 96816 569129 96844 579566
rect 97538 577552 97594 577561
rect 97538 577487 97594 577496
rect 97552 576910 97580 577487
rect 97540 576904 97592 576910
rect 97540 576846 97592 576852
rect 97908 576768 97960 576774
rect 97906 576736 97908 576745
rect 99196 576768 99248 576774
rect 97960 576736 97962 576745
rect 99196 576710 99248 576716
rect 97906 576671 97962 576680
rect 97632 575476 97684 575482
rect 97632 575418 97684 575424
rect 97644 575385 97672 575418
rect 97630 575376 97686 575385
rect 97630 575311 97686 575320
rect 97446 573472 97502 573481
rect 97446 573407 97502 573416
rect 97460 572762 97488 573407
rect 97448 572756 97500 572762
rect 97448 572698 97500 572704
rect 97078 571432 97134 571441
rect 97078 571367 97080 571376
rect 97132 571367 97134 571376
rect 97080 571338 97132 571344
rect 97908 570648 97960 570654
rect 97908 570590 97960 570596
rect 97920 570353 97948 570590
rect 97906 570344 97962 570353
rect 97906 570279 97962 570288
rect 97908 569220 97960 569226
rect 97908 569162 97960 569168
rect 97920 569129 97948 569162
rect 96802 569120 96858 569129
rect 96802 569055 96858 569064
rect 97906 569120 97962 569129
rect 97906 569055 97962 569064
rect 97906 565856 97962 565865
rect 97962 565814 98040 565842
rect 97906 565791 97962 565800
rect 96802 562320 96858 562329
rect 96802 562255 96858 562264
rect 96816 561746 96844 562255
rect 96804 561740 96856 561746
rect 96804 561682 96856 561688
rect 96894 560960 96950 560969
rect 96894 560895 96950 560904
rect 96802 559600 96858 559609
rect 96802 559535 96858 559544
rect 96816 558958 96844 559535
rect 96804 558952 96856 558958
rect 96804 558894 96856 558900
rect 96710 558784 96766 558793
rect 96710 558719 96766 558728
rect 96802 556880 96858 556889
rect 96802 556815 96858 556824
rect 95514 552528 95570 552537
rect 95514 552463 95570 552472
rect 96618 552528 96674 552537
rect 96618 552463 96674 552472
rect 95528 540938 95556 552463
rect 96710 543008 96766 543017
rect 96710 542943 96766 542952
rect 95516 540932 95568 540938
rect 95516 540874 95568 540880
rect 96618 538928 96674 538937
rect 96618 538863 96674 538872
rect 96632 537538 96660 538863
rect 96620 537532 96672 537538
rect 96620 537474 96672 537480
rect 95422 527776 95478 527785
rect 95422 527711 95478 527720
rect 95332 478168 95384 478174
rect 95332 478110 95384 478116
rect 96724 469878 96752 542943
rect 96816 530602 96844 556815
rect 96908 538898 96936 560895
rect 97170 558784 97226 558793
rect 97170 558719 97172 558728
rect 97224 558719 97226 558728
rect 97172 558690 97224 558696
rect 96986 552800 97042 552809
rect 96986 552735 97042 552744
rect 97000 552090 97028 552735
rect 96988 552084 97040 552090
rect 96988 552026 97040 552032
rect 97906 550760 97962 550769
rect 97906 550695 97962 550704
rect 97920 550662 97948 550695
rect 97908 550656 97960 550662
rect 97908 550598 97960 550604
rect 97078 549400 97134 549409
rect 97078 549335 97080 549344
rect 97132 549335 97134 549344
rect 97080 549306 97132 549312
rect 96986 545728 97042 545737
rect 96986 545663 97042 545672
rect 96896 538892 96948 538898
rect 96896 538834 96948 538840
rect 96804 530596 96856 530602
rect 96804 530538 96856 530544
rect 96712 469872 96764 469878
rect 96712 469814 96764 469820
rect 97000 461553 97028 545663
rect 97354 544368 97410 544377
rect 97354 544303 97410 544312
rect 97368 543794 97396 544303
rect 97356 543788 97408 543794
rect 97356 543730 97408 543736
rect 98012 522306 98040 565814
rect 98000 522300 98052 522306
rect 98000 522242 98052 522248
rect 98644 475380 98696 475386
rect 98644 475322 98696 475328
rect 96986 461544 97042 461553
rect 96986 461479 97042 461488
rect 95238 454744 95294 454753
rect 95238 454679 95294 454688
rect 96712 452600 96764 452606
rect 96712 452542 96764 452548
rect 96618 444272 96674 444281
rect 96618 444207 96674 444216
rect 96632 443057 96660 444207
rect 96618 443048 96674 443057
rect 96618 442983 96674 442992
rect 95240 442264 95292 442270
rect 95240 442206 95292 442212
rect 94136 440292 94188 440298
rect 94136 440234 94188 440240
rect 95148 440292 95200 440298
rect 95148 440234 95200 440240
rect 92662 434752 92718 434761
rect 92662 434687 92718 434696
rect 88720 434302 89056 434330
rect 89792 434302 90128 434330
rect 91066 434574 91140 434602
rect 91066 434316 91094 434574
rect 87142 434279 87198 434288
rect 85868 434219 85896 434279
rect 87156 434219 87184 434279
rect 71780 434182 71832 434188
rect 82800 434166 82952 434194
rect 92676 434058 92704 434687
rect 94148 434330 94176 440234
rect 94228 437436 94280 437442
rect 94228 437378 94280 437384
rect 94240 434353 94268 437378
rect 95252 437170 95280 442206
rect 95240 437164 95292 437170
rect 95240 437106 95292 437112
rect 95884 437164 95936 437170
rect 95884 437106 95936 437112
rect 95896 436150 95924 437106
rect 95884 436144 95936 436150
rect 95884 436086 95936 436092
rect 93840 434302 94176 434330
rect 94226 434344 94282 434353
rect 94282 434302 94576 434330
rect 94226 434279 94282 434288
rect 94240 434219 94268 434279
rect 95896 434194 95924 436086
rect 96632 434602 96660 442983
rect 96724 441614 96752 452542
rect 96724 441586 96936 441614
rect 96586 434574 96660 434602
rect 96586 434316 96614 434574
rect 96908 434330 96936 441586
rect 98656 439521 98684 475322
rect 99208 456074 99236 576710
rect 99300 572665 99328 702714
rect 101402 585168 101458 585177
rect 101402 585103 101458 585112
rect 100852 572756 100904 572762
rect 100852 572698 100904 572704
rect 99286 572656 99342 572665
rect 99286 572591 99342 572600
rect 99300 572014 99328 572591
rect 99288 572008 99340 572014
rect 99288 571950 99340 571956
rect 100024 571396 100076 571402
rect 100024 571338 100076 571344
rect 100036 547913 100064 571338
rect 100760 558748 100812 558754
rect 100760 558690 100812 558696
rect 100116 549364 100168 549370
rect 100116 549306 100168 549312
rect 100022 547904 100078 547913
rect 100022 547839 100078 547848
rect 100024 533384 100076 533390
rect 100024 533326 100076 533332
rect 99196 456068 99248 456074
rect 99196 456010 99248 456016
rect 98642 439512 98698 439521
rect 98642 439447 98698 439456
rect 100036 435033 100064 533326
rect 100128 507929 100156 549306
rect 100114 507920 100170 507929
rect 100114 507855 100170 507864
rect 100116 465724 100168 465730
rect 100116 465666 100168 465672
rect 100128 437442 100156 465666
rect 100772 443698 100800 558690
rect 100864 525094 100892 572698
rect 100852 525088 100904 525094
rect 100852 525030 100904 525036
rect 101416 446457 101444 585103
rect 101508 576774 101536 702918
rect 105464 700330 105492 703520
rect 119344 703180 119396 703186
rect 119344 703122 119396 703128
rect 116584 702840 116636 702846
rect 116584 702782 116636 702788
rect 106924 702636 106976 702642
rect 106924 702578 106976 702584
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 104162 582584 104218 582593
rect 104162 582519 104218 582528
rect 102782 581632 102838 581641
rect 102782 581567 102838 581576
rect 101496 576768 101548 576774
rect 101496 576710 101548 576716
rect 102232 519580 102284 519586
rect 102232 519522 102284 519528
rect 101402 446448 101458 446457
rect 101402 446383 101458 446392
rect 100760 443692 100812 443698
rect 100760 443634 100812 443640
rect 102140 442060 102192 442066
rect 102140 442002 102192 442008
rect 100116 437436 100168 437442
rect 100116 437378 100168 437384
rect 100022 435024 100078 435033
rect 100022 434959 100078 434968
rect 100036 434602 100064 434959
rect 101218 434888 101274 434897
rect 101218 434823 101274 434832
rect 100036 434574 100110 434602
rect 97170 434344 97226 434353
rect 96908 434302 97170 434330
rect 97226 434302 97336 434330
rect 100082 434316 100110 434574
rect 101232 434330 101260 434823
rect 102152 434330 102180 442002
rect 102244 441614 102272 519522
rect 102796 442066 102824 581567
rect 103428 570648 103480 570654
rect 103428 570590 103480 570596
rect 103440 569294 103468 570590
rect 103428 569288 103480 569294
rect 103428 569230 103480 569236
rect 103520 567860 103572 567866
rect 103520 567802 103572 567808
rect 103532 448526 103560 567802
rect 103520 448520 103572 448526
rect 103520 448462 103572 448468
rect 103704 448520 103756 448526
rect 103704 448462 103756 448468
rect 102784 442060 102836 442066
rect 102784 442002 102836 442008
rect 102796 441658 102824 442002
rect 102784 441652 102836 441658
rect 102244 441586 102640 441614
rect 102784 441594 102836 441600
rect 103716 441614 103744 448462
rect 103716 441586 103928 441614
rect 102612 434353 102640 441586
rect 103796 436212 103848 436218
rect 103796 436154 103848 436160
rect 102598 434344 102654 434353
rect 101232 434302 101568 434330
rect 102152 434302 102304 434330
rect 97170 434279 97226 434288
rect 103808 434330 103836 436154
rect 102654 434302 103040 434330
rect 103592 434302 103836 434330
rect 103900 434330 103928 441586
rect 104176 435305 104204 582519
rect 105544 581052 105596 581058
rect 105544 580994 105596 581000
rect 105556 439550 105584 580994
rect 106936 575482 106964 702578
rect 107660 583840 107712 583846
rect 107660 583782 107712 583788
rect 106924 575476 106976 575482
rect 106924 575418 106976 575424
rect 106924 572008 106976 572014
rect 106924 571950 106976 571956
rect 106936 458833 106964 571950
rect 107016 458856 107068 458862
rect 106922 458824 106978 458833
rect 107016 458798 107068 458804
rect 106922 458759 106978 458768
rect 107028 441614 107056 458798
rect 106660 441586 107056 441614
rect 105544 439544 105596 439550
rect 105544 439486 105596 439492
rect 106096 438184 106148 438190
rect 106096 438126 106148 438132
rect 106108 437510 106136 438126
rect 106660 437578 106688 441586
rect 106648 437572 106700 437578
rect 106648 437514 106700 437520
rect 106096 437504 106148 437510
rect 106096 437446 106148 437452
rect 104624 437436 104676 437442
rect 104624 437378 104676 437384
rect 104636 436218 104664 437378
rect 104624 436212 104676 436218
rect 104624 436154 104676 436160
rect 104162 435296 104218 435305
rect 104162 435231 104218 435240
rect 104162 434344 104218 434353
rect 103900 434302 104162 434330
rect 102598 434279 102654 434288
rect 106108 434330 106136 437446
rect 106660 434330 106688 437514
rect 106738 436384 106794 436393
rect 106738 436319 106794 436328
rect 104218 434302 104328 434330
rect 105800 434302 106136 434330
rect 106352 434302 106688 434330
rect 106752 434330 106780 436319
rect 107672 436121 107700 583782
rect 110420 582412 110472 582418
rect 110420 582354 110472 582360
rect 108304 543788 108356 543794
rect 108304 543730 108356 543736
rect 108316 441614 108344 543730
rect 109684 482316 109736 482322
rect 109684 482258 109736 482264
rect 109040 445052 109092 445058
rect 109040 444994 109092 445000
rect 108132 441586 108344 441614
rect 109052 441614 109080 444994
rect 109052 441586 109448 441614
rect 108132 440366 108160 441586
rect 108120 440360 108172 440366
rect 108120 440302 108172 440308
rect 107658 436112 107714 436121
rect 107658 436047 107714 436056
rect 108132 434330 108160 440302
rect 109130 436248 109186 436257
rect 109130 436183 109186 436192
rect 108210 436112 108266 436121
rect 108210 436047 108266 436056
rect 108224 434353 108252 436047
rect 106752 434302 107088 434330
rect 107824 434302 108160 434330
rect 108210 434344 108266 434353
rect 104162 434279 104218 434288
rect 109144 434330 109172 436183
rect 108266 434302 108560 434330
rect 109144 434302 109296 434330
rect 108210 434279 108266 434288
rect 97184 434219 97212 434279
rect 102612 434219 102640 434279
rect 104176 434219 104204 434279
rect 108224 434219 108252 434279
rect 95896 434166 96048 434194
rect 92552 434030 92704 434058
rect 71226 433936 71282 433945
rect 100574 433936 100630 433945
rect 71282 433894 71576 433922
rect 71226 433871 71282 433880
rect 109420 433922 109448 441586
rect 109696 434790 109724 482258
rect 110432 436121 110460 582354
rect 113364 579692 113416 579698
rect 113364 579634 113416 579640
rect 111800 552084 111852 552090
rect 111800 552026 111852 552032
rect 111064 487824 111116 487830
rect 111064 487766 111116 487772
rect 110418 436112 110474 436121
rect 110418 436047 110474 436056
rect 110970 436112 111026 436121
rect 110970 436047 111026 436056
rect 109684 434784 109736 434790
rect 109684 434726 109736 434732
rect 109590 433936 109646 433945
rect 100630 433894 100832 433922
rect 109420 433894 109590 433922
rect 100574 433871 100630 433880
rect 109646 433894 109848 433922
rect 109590 433871 109646 433880
rect 72608 433832 72660 433838
rect 70858 433800 70914 433809
rect 72312 433780 72608 433786
rect 87970 433800 88026 433809
rect 72312 433774 72660 433780
rect 72312 433758 72648 433774
rect 74000 433770 74336 433786
rect 73988 433764 74336 433770
rect 70858 433735 70914 433744
rect 70872 433702 70900 433735
rect 74040 433758 74336 433764
rect 98458 433800 98514 433809
rect 88026 433758 88320 433786
rect 87970 433735 88026 433744
rect 98514 433758 98808 433786
rect 98458 433735 98514 433744
rect 73988 433706 74040 433712
rect 69204 433696 69256 433702
rect 70860 433696 70912 433702
rect 69256 433644 69552 433650
rect 69204 433638 69552 433644
rect 70860 433638 70912 433644
rect 73434 433664 73490 433673
rect 69216 433622 69552 433638
rect 78402 433664 78458 433673
rect 73490 433622 73784 433650
rect 73434 433599 73490 433608
rect 79598 433664 79654 433673
rect 78458 433622 78568 433650
rect 79304 433622 79598 433650
rect 78402 433599 78458 433608
rect 79598 433599 79654 433608
rect 87326 433664 87382 433673
rect 89994 433664 90050 433673
rect 87382 433622 87584 433650
rect 87326 433599 87382 433608
rect 91466 433664 91522 433673
rect 90050 433622 90344 433650
rect 89994 433599 90050 433608
rect 93490 433664 93546 433673
rect 91522 433622 91816 433650
rect 93288 433622 93490 433650
rect 91466 433599 91522 433608
rect 93490 433599 93546 433608
rect 95146 433664 95202 433673
rect 98366 433664 98422 433673
rect 95202 433622 95312 433650
rect 98072 433622 98366 433650
rect 95146 433599 95202 433608
rect 99838 433664 99894 433673
rect 99544 433622 99838 433650
rect 98366 433599 98422 433608
rect 105174 433664 105230 433673
rect 105064 433622 105174 433650
rect 99838 433599 99894 433608
rect 105174 433599 105230 433608
rect 110418 433664 110474 433673
rect 110984 433650 111012 436047
rect 111076 433838 111104 487766
rect 111812 434858 111840 552026
rect 112720 471300 112772 471306
rect 112720 471242 112772 471248
rect 111800 434852 111852 434858
rect 111800 434794 111852 434800
rect 112628 434852 112680 434858
rect 112628 434794 112680 434800
rect 112640 434714 112668 434794
rect 112456 434686 112668 434714
rect 112456 434058 112484 434686
rect 112456 434030 112608 434058
rect 111064 433832 111116 433838
rect 111064 433774 111116 433780
rect 111616 433696 111668 433702
rect 110474 433622 110584 433650
rect 110984 433644 111616 433650
rect 110984 433638 111668 433644
rect 111706 433664 111762 433673
rect 110984 433622 111656 433638
rect 110418 433599 110474 433608
rect 111762 433622 112056 433650
rect 111706 433599 111762 433608
rect 82082 391096 82138 391105
rect 81544 391054 82082 391082
rect 77404 390782 77832 390810
rect 72422 390416 72478 390425
rect 68802 390182 68830 390388
rect 69124 390374 69368 390402
rect 69768 390374 70104 390402
rect 70412 390374 70840 390402
rect 70964 390374 71576 390402
rect 71884 390374 72422 390402
rect 68790 390176 68842 390182
rect 68790 390118 68842 390124
rect 69020 387048 69072 387054
rect 69020 386990 69072 386996
rect 69032 301306 69060 386990
rect 69124 380186 69152 390374
rect 69768 387054 69796 390374
rect 69756 387048 69808 387054
rect 69756 386990 69808 386996
rect 70306 385112 70362 385121
rect 70306 385047 70362 385056
rect 69112 380180 69164 380186
rect 69112 380122 69164 380128
rect 69662 338056 69718 338065
rect 69662 337991 69718 338000
rect 69676 336870 69704 337991
rect 69664 336864 69716 336870
rect 69664 336806 69716 336812
rect 69110 314936 69166 314945
rect 69110 314871 69166 314880
rect 69020 301300 69072 301306
rect 69020 301242 69072 301248
rect 68652 284980 68704 284986
rect 68652 284922 68704 284928
rect 69018 284880 69074 284889
rect 69018 284815 69074 284824
rect 69032 283778 69060 284815
rect 68986 283750 69060 283778
rect 68986 283492 69014 283750
rect 69124 283150 69152 314871
rect 69676 283506 69704 336806
rect 70320 314945 70348 385047
rect 70306 314936 70362 314945
rect 70306 314871 70362 314880
rect 69756 302320 69808 302326
rect 69756 302262 69808 302268
rect 69216 283478 69704 283506
rect 69112 283144 69164 283150
rect 69112 283086 69164 283092
rect 68652 283076 68704 283082
rect 68652 283018 68704 283024
rect 68376 283008 68428 283014
rect 68376 282950 68428 282956
rect 68282 277400 68338 277409
rect 68282 277335 68284 277344
rect 68336 277335 68338 277344
rect 68284 277306 68336 277312
rect 68296 277275 68324 277306
rect 68284 261588 68336 261594
rect 68284 261530 68336 261536
rect 68190 258768 68246 258777
rect 68190 258703 68246 258712
rect 68204 258058 68232 258703
rect 68192 258052 68244 258058
rect 68192 257994 68244 258000
rect 67638 241360 67694 241369
rect 67638 241295 67694 241304
rect 67546 129840 67602 129849
rect 67546 129775 67602 129784
rect 67546 102640 67602 102649
rect 67546 102575 67602 102584
rect 67560 102241 67588 102575
rect 67546 102232 67602 102241
rect 67546 102167 67602 102176
rect 67454 98016 67510 98025
rect 67454 97951 67510 97960
rect 67180 79348 67232 79354
rect 67180 79290 67232 79296
rect 66076 68400 66128 68406
rect 66076 68342 66128 68348
rect 65984 17264 66036 17270
rect 65984 17206 66036 17212
rect 64788 15972 64840 15978
rect 64788 15914 64840 15920
rect 62028 3596 62080 3602
rect 62028 3538 62080 3544
rect 61948 3454 62068 3482
rect 64800 3466 64828 15914
rect 62040 480 62068 3454
rect 64328 3460 64380 3466
rect 64328 3402 64380 3408
rect 64788 3460 64840 3466
rect 64788 3402 64840 3408
rect 63222 3360 63278 3369
rect 63222 3295 63278 3304
rect 63236 480 63264 3295
rect 64340 480 64368 3402
rect 66088 3194 66116 68342
rect 67560 56574 67588 102167
rect 67652 92886 67680 241295
rect 68296 233986 68324 261530
rect 68388 241505 68416 282950
rect 68558 241768 68614 241777
rect 68558 241703 68560 241712
rect 68612 241703 68614 241712
rect 68560 241674 68612 241680
rect 68374 241496 68430 241505
rect 68374 241431 68430 241440
rect 68284 233980 68336 233986
rect 68284 233922 68336 233928
rect 68664 232665 68692 283018
rect 69216 283014 69244 283478
rect 69768 283014 69796 302262
rect 70412 288425 70440 390374
rect 70964 373994 70992 390374
rect 71884 389065 71912 390374
rect 77206 390416 77262 390425
rect 72422 390351 72478 390360
rect 72528 390374 72864 390402
rect 73264 390374 73600 390402
rect 74000 390374 74336 390402
rect 74644 390374 75072 390402
rect 75288 390374 75624 390402
rect 75932 390374 76360 390402
rect 76760 390374 77206 390402
rect 72528 389162 72556 390374
rect 72516 389156 72568 389162
rect 72516 389098 72568 389104
rect 71870 389056 71926 389065
rect 71870 388991 71926 389000
rect 72974 384432 73030 384441
rect 72974 384367 73030 384376
rect 71686 380896 71742 380905
rect 71686 380831 71742 380840
rect 70504 373966 70992 373994
rect 70504 328545 70532 373966
rect 70490 328536 70546 328545
rect 70490 328471 70546 328480
rect 71700 318073 71728 380831
rect 72988 325694 73016 384367
rect 73068 381540 73120 381546
rect 73068 381482 73120 381488
rect 72896 325666 73016 325694
rect 72422 319424 72478 319433
rect 72422 319359 72478 319368
rect 71686 318064 71742 318073
rect 71686 317999 71742 318008
rect 71688 313336 71740 313342
rect 71688 313278 71740 313284
rect 71044 298648 71096 298654
rect 71044 298590 71096 298596
rect 71056 289814 71084 298590
rect 70964 289786 71084 289814
rect 70398 288416 70454 288425
rect 70398 288351 70454 288360
rect 70964 287094 70992 289786
rect 71700 287706 71728 313278
rect 72436 291378 72464 319359
rect 72606 318880 72662 318889
rect 72606 318815 72662 318824
rect 72620 298654 72648 318815
rect 72896 316742 72924 325666
rect 72974 318880 73030 318889
rect 72974 318815 72976 318824
rect 73028 318815 73030 318824
rect 72976 318786 73028 318792
rect 72884 316736 72936 316742
rect 72884 316678 72936 316684
rect 72608 298648 72660 298654
rect 72608 298590 72660 298596
rect 72424 291372 72476 291378
rect 72424 291314 72476 291320
rect 72056 291236 72108 291242
rect 72056 291178 72108 291184
rect 71688 287700 71740 287706
rect 71688 287642 71740 287648
rect 70952 287088 71004 287094
rect 70952 287030 71004 287036
rect 70964 283234 70992 287030
rect 71180 283792 71236 283801
rect 71180 283727 71236 283736
rect 70656 283206 70992 283234
rect 71042 283248 71098 283257
rect 71194 283234 71222 283727
rect 71870 283520 71926 283529
rect 71760 283478 71870 283506
rect 72068 283506 72096 291178
rect 72436 283506 72464 291314
rect 73080 291242 73108 381482
rect 73264 300257 73292 390374
rect 74000 387802 74028 390374
rect 73988 387796 74040 387802
rect 73988 387738 74040 387744
rect 74264 387796 74316 387802
rect 74264 387738 74316 387744
rect 73802 343768 73858 343777
rect 73802 343703 73858 343712
rect 73816 343670 73844 343703
rect 73804 343664 73856 343670
rect 73804 343606 73856 343612
rect 73250 300248 73306 300257
rect 73250 300183 73306 300192
rect 73802 300248 73858 300257
rect 73802 300183 73858 300192
rect 73068 291236 73120 291242
rect 73068 291178 73120 291184
rect 73816 287745 73844 300183
rect 73802 287736 73858 287745
rect 73802 287671 73858 287680
rect 74080 286952 74132 286958
rect 74080 286894 74132 286900
rect 74092 285841 74120 286894
rect 74078 285832 74134 285841
rect 72516 285796 72568 285802
rect 74078 285767 74134 285776
rect 72516 285738 72568 285744
rect 71926 283478 72096 283506
rect 72312 283478 72464 283506
rect 72528 283506 72556 285738
rect 73526 283520 73582 283529
rect 72528 283478 72864 283506
rect 73416 283478 73526 283506
rect 71870 283455 71926 283464
rect 73526 283455 73582 283464
rect 71884 283395 71912 283455
rect 74092 283370 74120 285767
rect 74276 284209 74304 387738
rect 74644 336054 74672 390374
rect 75288 387802 75316 390374
rect 75276 387796 75328 387802
rect 75276 387738 75328 387744
rect 75826 386336 75882 386345
rect 75826 386271 75882 386280
rect 75182 379536 75238 379545
rect 75182 379471 75238 379480
rect 74632 336048 74684 336054
rect 74632 335990 74684 335996
rect 75196 313342 75224 379471
rect 75288 340950 75316 340981
rect 75276 340944 75328 340950
rect 75274 340912 75276 340921
rect 75328 340912 75330 340921
rect 75274 340847 75330 340856
rect 75184 313336 75236 313342
rect 75184 313278 75236 313284
rect 75184 294024 75236 294030
rect 75184 293966 75236 293972
rect 74540 287700 74592 287706
rect 74540 287642 74592 287648
rect 74262 284200 74318 284209
rect 74262 284135 74318 284144
rect 74552 283778 74580 287642
rect 74506 283750 74580 283778
rect 75046 283756 75098 283762
rect 74506 283492 74534 283750
rect 75046 283698 75098 283704
rect 75058 283492 75086 283698
rect 75196 283506 75224 293966
rect 75288 285870 75316 340847
rect 75840 322998 75868 386271
rect 75368 322992 75420 322998
rect 75368 322934 75420 322940
rect 75828 322992 75880 322998
rect 75828 322934 75880 322940
rect 75380 294030 75408 322934
rect 75828 313336 75880 313342
rect 75828 313278 75880 313284
rect 75840 312497 75868 313278
rect 75826 312488 75882 312497
rect 75826 312423 75882 312432
rect 75932 303634 75960 390374
rect 76760 389065 76788 390374
rect 77206 390351 77262 390360
rect 76010 389056 76066 389065
rect 76010 388991 76066 389000
rect 76746 389056 76802 389065
rect 76746 388991 76802 389000
rect 76024 376038 76052 388991
rect 76564 387660 76616 387666
rect 76564 387602 76616 387608
rect 76012 376032 76064 376038
rect 76012 375974 76064 375980
rect 75840 303606 75960 303634
rect 75840 302326 75868 303606
rect 75828 302320 75880 302326
rect 75828 302262 75880 302268
rect 75840 301481 75868 302262
rect 75826 301472 75882 301481
rect 75826 301407 75882 301416
rect 75368 294024 75420 294030
rect 75368 293966 75420 293972
rect 76196 290760 76248 290766
rect 76196 290702 76248 290708
rect 76208 289882 76236 290702
rect 76196 289876 76248 289882
rect 76196 289818 76248 289824
rect 75276 285864 75328 285870
rect 75276 285806 75328 285812
rect 75288 283762 75316 285806
rect 76208 283778 76236 289818
rect 76576 286958 76604 387602
rect 77300 387048 77352 387054
rect 77300 386990 77352 386996
rect 77312 338745 77340 386990
rect 77404 383042 77432 390782
rect 77482 390688 77538 390697
rect 77482 390623 77538 390632
rect 78968 390646 79120 390674
rect 77392 383036 77444 383042
rect 77392 382978 77444 382984
rect 77496 381546 77524 390623
rect 78048 390374 78384 390402
rect 78048 387054 78076 390374
rect 78968 389065 78996 390646
rect 79244 390374 79856 390402
rect 80592 390374 80928 390402
rect 78954 389056 79010 389065
rect 78954 388991 79010 389000
rect 78036 387048 78088 387054
rect 78036 386990 78088 386996
rect 78586 383752 78642 383761
rect 78586 383687 78642 383696
rect 77484 381540 77536 381546
rect 77484 381482 77536 381488
rect 77298 338736 77354 338745
rect 77298 338671 77354 338680
rect 78036 325712 78088 325718
rect 78036 325654 78088 325660
rect 76746 322960 76802 322969
rect 76746 322895 76802 322904
rect 76654 318744 76710 318753
rect 76654 318679 76710 318688
rect 76564 286952 76616 286958
rect 76564 286894 76616 286900
rect 76668 284374 76696 318679
rect 76760 290766 76788 322895
rect 77942 320784 77998 320793
rect 77942 320719 77998 320728
rect 77852 292664 77904 292670
rect 77852 292606 77904 292612
rect 77760 291848 77812 291854
rect 77760 291790 77812 291796
rect 77772 291310 77800 291790
rect 77760 291304 77812 291310
rect 77760 291246 77812 291252
rect 76748 290760 76800 290766
rect 76748 290702 76800 290708
rect 77392 286408 77444 286414
rect 77392 286350 77444 286356
rect 76656 284368 76708 284374
rect 76656 284310 76708 284316
rect 75276 283756 75328 283762
rect 75276 283698 75328 283704
rect 76162 283750 76236 283778
rect 76668 283778 76696 284310
rect 76668 283750 76742 283778
rect 75196 283478 75624 283506
rect 76162 283492 76190 283750
rect 76714 283492 76742 283750
rect 77404 283665 77432 286350
rect 77772 283778 77800 291246
rect 77864 285818 77892 292606
rect 77956 286414 77984 320719
rect 78048 292670 78076 325654
rect 78600 310486 78628 383687
rect 79244 373994 79272 390374
rect 80058 387968 80114 387977
rect 80058 387903 80114 387912
rect 79876 387796 79928 387802
rect 79876 387738 79928 387744
rect 78692 373966 79272 373994
rect 78128 310480 78180 310486
rect 78128 310422 78180 310428
rect 78588 310480 78640 310486
rect 78588 310422 78640 310428
rect 78140 309806 78168 310422
rect 78128 309800 78180 309806
rect 78128 309742 78180 309748
rect 78036 292664 78088 292670
rect 78036 292606 78088 292612
rect 78140 291854 78168 309742
rect 78692 303634 78720 373966
rect 79888 308446 79916 387738
rect 80072 387666 80100 387903
rect 80060 387660 80112 387666
rect 80060 387602 80112 387608
rect 80900 386306 80928 390374
rect 80992 390374 81328 390402
rect 80992 387705 81020 390374
rect 81544 388793 81572 391054
rect 82082 391031 82138 391040
rect 85486 391096 85542 391105
rect 89672 391096 89728 391105
rect 87984 391066 88288 391082
rect 85486 391031 85542 391040
rect 87972 391060 88288 391066
rect 82004 390374 82616 390402
rect 83016 390374 83352 390402
rect 83476 390374 84088 390402
rect 84304 390374 84824 390402
rect 81530 388784 81586 388793
rect 81530 388719 81586 388728
rect 81544 387802 81572 388719
rect 81532 387796 81584 387802
rect 81532 387738 81584 387744
rect 80978 387696 81034 387705
rect 80978 387631 81034 387640
rect 80888 386300 80940 386306
rect 80888 386242 80940 386248
rect 81348 386300 81400 386306
rect 81348 386242 81400 386248
rect 79966 385112 80022 385121
rect 79966 385047 80022 385056
rect 79876 308440 79928 308446
rect 79876 308382 79928 308388
rect 79874 304192 79930 304201
rect 79874 304127 79930 304136
rect 78600 303606 78720 303634
rect 78600 296002 78628 303606
rect 78588 295996 78640 296002
rect 78588 295938 78640 295944
rect 78680 295384 78732 295390
rect 78680 295326 78732 295332
rect 78128 291848 78180 291854
rect 78128 291790 78180 291796
rect 78692 287774 78720 295326
rect 79888 292641 79916 304127
rect 79980 295390 80008 385047
rect 81254 377360 81310 377369
rect 81254 377295 81310 377304
rect 81268 331362 81296 377295
rect 80704 331356 80756 331362
rect 80704 331298 80756 331304
rect 81256 331356 81308 331362
rect 81256 331298 81308 331304
rect 80244 327752 80296 327758
rect 80244 327694 80296 327700
rect 79968 295384 80020 295390
rect 79968 295326 80020 295332
rect 78770 292632 78826 292641
rect 78770 292567 78826 292576
rect 79874 292632 79930 292641
rect 79874 292567 79930 292576
rect 78680 287768 78732 287774
rect 78680 287710 78732 287716
rect 77944 286408 77996 286414
rect 77944 286350 77996 286356
rect 77864 285790 77984 285818
rect 77772 283750 77846 283778
rect 77390 283656 77446 283665
rect 77390 283591 77446 283600
rect 77404 283370 77432 283591
rect 77818 283492 77846 283750
rect 77956 283506 77984 285790
rect 78784 283506 78812 292567
rect 79968 288448 80020 288454
rect 79968 288390 80020 288396
rect 79140 287768 79192 287774
rect 79140 287710 79192 287716
rect 79152 283506 79180 287710
rect 79980 287054 80008 288390
rect 79980 287026 80100 287054
rect 80072 283778 80100 287026
rect 80026 283750 80100 283778
rect 77956 283478 78384 283506
rect 78784 283478 78936 283506
rect 79152 283478 79488 283506
rect 80026 283492 80054 283750
rect 80256 283506 80284 327694
rect 80716 292574 80744 331298
rect 81360 319569 81388 386242
rect 82004 373994 82032 390374
rect 83016 389230 83044 390374
rect 83004 389224 83056 389230
rect 83004 389166 83056 389172
rect 82726 387696 82782 387705
rect 82726 387631 82782 387640
rect 81544 373966 82032 373994
rect 81544 345014 81572 373966
rect 81452 344986 81572 345014
rect 81452 339522 81480 344986
rect 81440 339516 81492 339522
rect 81440 339458 81492 339464
rect 81452 338774 81480 339458
rect 81440 338768 81492 338774
rect 81440 338710 81492 338716
rect 82634 333296 82690 333305
rect 82634 333231 82690 333240
rect 81346 319560 81402 319569
rect 81346 319495 81402 319504
rect 80716 292546 80836 292574
rect 80808 287337 80836 292546
rect 81992 289876 82044 289882
rect 81992 289818 82044 289824
rect 80794 287328 80850 287337
rect 80794 287263 80850 287272
rect 80808 283506 80836 287263
rect 82004 283506 82032 289818
rect 82648 285977 82676 333231
rect 82740 289882 82768 387631
rect 83476 376038 83504 390374
rect 84304 388362 84332 390374
rect 85362 390130 85390 390388
rect 85362 390102 85436 390130
rect 84120 388334 84332 388362
rect 83464 376032 83516 376038
rect 83464 375974 83516 375980
rect 84120 356726 84148 388334
rect 85408 387870 85436 390102
rect 85396 387864 85448 387870
rect 85396 387806 85448 387812
rect 85394 380216 85450 380225
rect 85394 380151 85450 380160
rect 85302 378720 85358 378729
rect 85302 378655 85358 378664
rect 84108 356720 84160 356726
rect 84108 356662 84160 356668
rect 83554 339552 83610 339561
rect 83554 339487 83556 339496
rect 83608 339487 83610 339496
rect 83556 339458 83608 339464
rect 84106 329080 84162 329089
rect 84106 329015 84162 329024
rect 84120 325718 84148 329015
rect 84108 325712 84160 325718
rect 84108 325654 84160 325660
rect 83462 323640 83518 323649
rect 83462 323575 83518 323584
rect 82912 313336 82964 313342
rect 82912 313278 82964 313284
rect 82924 306374 82952 313278
rect 82924 306346 83412 306374
rect 82728 289876 82780 289882
rect 82728 289818 82780 289824
rect 83004 288516 83056 288522
rect 83004 288458 83056 288464
rect 82912 287020 82964 287026
rect 82912 286962 82964 286968
rect 82634 285968 82690 285977
rect 82634 285903 82690 285912
rect 82648 283506 82676 285903
rect 82924 283506 82952 286962
rect 80256 283478 80592 283506
rect 80808 283478 81144 283506
rect 81696 283478 82032 283506
rect 82248 283478 82676 283506
rect 82800 283478 82952 283506
rect 83016 283506 83044 288458
rect 83384 285954 83412 306346
rect 83476 288522 83504 323575
rect 85316 316062 85344 378655
rect 84200 316056 84252 316062
rect 84200 315998 84252 316004
rect 85304 316056 85356 316062
rect 85304 315998 85356 316004
rect 84108 305652 84160 305658
rect 84108 305594 84160 305600
rect 84120 289105 84148 305594
rect 84106 289096 84162 289105
rect 84106 289031 84162 289040
rect 83464 288516 83516 288522
rect 83464 288458 83516 288464
rect 83384 285926 83504 285954
rect 83476 283506 83504 285926
rect 84212 283506 84240 315998
rect 85408 292574 85436 380151
rect 85316 292546 85436 292574
rect 85316 287337 85344 292546
rect 85500 291417 85528 391031
rect 88024 391054 88288 391060
rect 87972 391002 88024 391008
rect 85592 390374 86112 390402
rect 85592 354006 85620 390374
rect 86834 390130 86862 390388
rect 87064 390374 87584 390402
rect 86834 390102 86908 390130
rect 86222 389056 86278 389065
rect 86222 388991 86278 389000
rect 86236 369073 86264 388991
rect 86880 387122 86908 390102
rect 86868 387116 86920 387122
rect 86868 387058 86920 387064
rect 86866 382392 86922 382401
rect 86866 382327 86922 382336
rect 86222 369064 86278 369073
rect 86222 368999 86278 369008
rect 86776 367804 86828 367810
rect 86776 367746 86828 367752
rect 85580 354000 85632 354006
rect 85580 353942 85632 353948
rect 85670 320920 85726 320929
rect 85670 320855 85726 320864
rect 85580 291848 85632 291854
rect 85580 291790 85632 291796
rect 85486 291408 85542 291417
rect 85486 291343 85542 291352
rect 85302 287328 85358 287337
rect 85302 287263 85358 287272
rect 85316 283506 85344 287263
rect 85500 287026 85528 291343
rect 85488 287020 85540 287026
rect 85488 286962 85540 286968
rect 85592 283778 85620 291790
rect 85684 287774 85712 320855
rect 86788 299130 86816 367746
rect 86880 301510 86908 382327
rect 87064 305658 87092 390374
rect 88260 390318 88288 391054
rect 89594 391048 89622 391068
rect 89594 391040 89672 391048
rect 92754 391096 92810 391105
rect 89728 391054 89944 391082
rect 89594 391031 89728 391040
rect 89594 391020 89714 391031
rect 89916 390998 89944 391054
rect 92810 391054 93440 391082
rect 99360 391066 99512 391082
rect 99360 391060 99524 391066
rect 99360 391054 99472 391060
rect 92754 391031 92810 391040
rect 89904 390992 89956 390998
rect 89904 390934 89956 390940
rect 92940 390992 92992 390998
rect 92940 390934 92992 390940
rect 88872 390374 89208 390402
rect 88248 390312 88300 390318
rect 88248 390254 88300 390260
rect 88984 390312 89036 390318
rect 88984 390254 89036 390260
rect 88246 373280 88302 373289
rect 88246 373215 88302 373224
rect 88260 334014 88288 373215
rect 88996 365022 89024 390254
rect 89180 389065 89208 390374
rect 89732 390374 90344 390402
rect 89166 389056 89222 389065
rect 89166 388991 89222 389000
rect 89626 387152 89682 387161
rect 89626 387087 89682 387096
rect 89534 385656 89590 385665
rect 89534 385591 89590 385600
rect 88984 365016 89036 365022
rect 88984 364958 89036 364964
rect 89444 359508 89496 359514
rect 89444 359450 89496 359456
rect 88248 334008 88300 334014
rect 88248 333950 88300 333956
rect 88156 321768 88208 321774
rect 88156 321710 88208 321716
rect 88168 320210 88196 321710
rect 88156 320204 88208 320210
rect 88156 320146 88208 320152
rect 88168 319433 88196 320146
rect 88154 319424 88210 319433
rect 88154 319359 88210 319368
rect 87052 305652 87104 305658
rect 87052 305594 87104 305600
rect 86868 301504 86920 301510
rect 86868 301446 86920 301452
rect 85764 299124 85816 299130
rect 85764 299066 85816 299072
rect 86776 299124 86828 299130
rect 86776 299066 86828 299072
rect 85672 287768 85724 287774
rect 85672 287710 85724 287716
rect 83016 283478 83352 283506
rect 83476 283478 83904 283506
rect 84212 283478 84792 283506
rect 85008 283478 85344 283506
rect 85546 283750 85620 283778
rect 85546 283492 85574 283750
rect 85776 283506 85804 299066
rect 86788 298178 86816 299066
rect 86776 298172 86828 298178
rect 86776 298114 86828 298120
rect 88260 292574 88288 333950
rect 88076 292546 88288 292574
rect 88076 291281 88104 292546
rect 88062 291272 88118 291281
rect 88062 291207 88118 291216
rect 86316 287768 86368 287774
rect 86316 287710 86368 287716
rect 86328 283506 86356 287710
rect 87510 285424 87566 285433
rect 87510 285359 87566 285368
rect 87524 283506 87552 285359
rect 88076 283506 88104 291207
rect 88616 288380 88668 288386
rect 88616 288322 88668 288328
rect 88628 283506 88656 288322
rect 89456 287473 89484 359450
rect 89548 289950 89576 385591
rect 89536 289944 89588 289950
rect 89536 289886 89588 289892
rect 89166 287464 89222 287473
rect 89166 287399 89222 287408
rect 89442 287464 89498 287473
rect 89442 287399 89498 287408
rect 89180 283506 89208 287399
rect 89548 283506 89576 289886
rect 89640 288561 89668 387087
rect 89732 333266 89760 390374
rect 91066 390130 91094 390388
rect 91204 390374 91632 390402
rect 91848 390374 92368 390402
rect 91066 390102 91140 390130
rect 91112 388482 91140 390102
rect 91100 388476 91152 388482
rect 91100 388418 91152 388424
rect 90364 387864 90416 387870
rect 90364 387806 90416 387812
rect 90376 366382 90404 387806
rect 91204 387036 91232 390374
rect 91112 387008 91232 387036
rect 91112 382401 91140 387008
rect 91848 383654 91876 390374
rect 92952 386414 92980 390934
rect 93214 389056 93270 389065
rect 93214 388991 93270 389000
rect 92952 386386 93164 386414
rect 91836 383648 91888 383654
rect 91836 383590 91888 383596
rect 91848 382498 91876 383590
rect 91192 382492 91244 382498
rect 91192 382434 91244 382440
rect 91836 382492 91888 382498
rect 91836 382434 91888 382440
rect 91098 382392 91154 382401
rect 91098 382327 91154 382336
rect 90364 366376 90416 366382
rect 90364 366318 90416 366324
rect 89720 333260 89772 333266
rect 89720 333202 89772 333208
rect 89720 329112 89772 329118
rect 89720 329054 89772 329060
rect 89732 327758 89760 329054
rect 89720 327752 89772 327758
rect 89720 327694 89772 327700
rect 91204 321774 91232 382434
rect 92388 376100 92440 376106
rect 92388 376042 92440 376048
rect 92400 335374 92428 376042
rect 93136 363662 93164 386386
rect 93228 380186 93256 388991
rect 93412 388346 93440 391054
rect 99472 391002 99524 391008
rect 106648 391060 106700 391066
rect 106648 391002 106700 391008
rect 98472 390646 98624 390674
rect 93826 390130 93854 390388
rect 93964 390374 94392 390402
rect 94792 390374 95128 390402
rect 95252 390374 95864 390402
rect 93826 390102 93900 390130
rect 93872 388929 93900 390102
rect 93858 388920 93914 388929
rect 93858 388855 93914 388864
rect 93400 388340 93452 388346
rect 93400 388282 93452 388288
rect 93860 387048 93912 387054
rect 93766 387016 93822 387025
rect 93860 386990 93912 386996
rect 93766 386951 93822 386960
rect 93216 380180 93268 380186
rect 93216 380122 93268 380128
rect 93674 364984 93730 364993
rect 93674 364919 93730 364928
rect 93124 363656 93176 363662
rect 93124 363598 93176 363604
rect 93688 346458 93716 364919
rect 93124 346452 93176 346458
rect 93124 346394 93176 346400
rect 93676 346452 93728 346458
rect 93676 346394 93728 346400
rect 92388 335368 92440 335374
rect 92388 335310 92440 335316
rect 92400 332761 92428 335310
rect 92386 332752 92442 332761
rect 92386 332687 92442 332696
rect 92386 322144 92442 322153
rect 92386 322079 92442 322088
rect 91192 321768 91244 321774
rect 91192 321710 91244 321716
rect 92400 312089 92428 322079
rect 91190 312080 91246 312089
rect 91190 312015 91246 312024
rect 92386 312080 92442 312089
rect 92386 312015 92442 312024
rect 91006 308408 91062 308417
rect 91006 308343 91062 308352
rect 89718 292632 89774 292641
rect 89718 292567 89774 292576
rect 91020 292574 91048 308343
rect 91204 306374 91232 312015
rect 91204 306346 91784 306374
rect 89626 288552 89682 288561
rect 89626 288487 89682 288496
rect 89640 288386 89668 288487
rect 89628 288380 89680 288386
rect 89628 288322 89680 288328
rect 85776 283478 86112 283506
rect 86328 283478 86664 283506
rect 87216 283478 87552 283506
rect 87768 283478 88104 283506
rect 88320 283478 88656 283506
rect 88872 283478 89208 283506
rect 89424 283478 89576 283506
rect 89732 283506 89760 292567
rect 90836 292546 91048 292574
rect 90836 289921 90864 292546
rect 90822 289912 90878 289921
rect 90822 289847 90878 289856
rect 90836 283506 90864 289847
rect 91468 287088 91520 287094
rect 91468 287030 91520 287036
rect 91376 283620 91428 283626
rect 91376 283562 91428 283568
rect 91388 283506 91416 283562
rect 89732 283478 89976 283506
rect 90528 283478 90864 283506
rect 91080 283478 91416 283506
rect 73968 283342 74120 283370
rect 77280 283342 77432 283370
rect 71098 283220 71222 283234
rect 71098 283206 71208 283220
rect 71042 283183 71098 283192
rect 69848 283144 69900 283150
rect 69900 283092 70104 283098
rect 69848 283086 70104 283092
rect 69860 283070 70104 283086
rect 80256 283082 80284 283478
rect 80244 283076 80296 283082
rect 80244 283018 80296 283024
rect 84764 283014 84792 283478
rect 91480 283234 91508 287030
rect 91756 283506 91784 306346
rect 93032 286340 93084 286346
rect 93032 286282 93084 286288
rect 93044 283506 93072 286282
rect 93136 283626 93164 346394
rect 93674 304192 93730 304201
rect 93674 304127 93730 304136
rect 93688 287162 93716 304127
rect 93780 294030 93808 386951
rect 93872 370530 93900 386990
rect 93964 373318 93992 390374
rect 94594 388920 94650 388929
rect 94594 388855 94650 388864
rect 93952 373312 94004 373318
rect 93952 373254 94004 373260
rect 93860 370524 93912 370530
rect 93860 370466 93912 370472
rect 94608 311166 94636 388855
rect 94792 387054 94820 390374
rect 94780 387048 94832 387054
rect 94780 386990 94832 386996
rect 95148 378276 95200 378282
rect 95148 378218 95200 378224
rect 95056 362228 95108 362234
rect 95056 362170 95108 362176
rect 94596 311160 94648 311166
rect 94596 311102 94648 311108
rect 95068 296714 95096 362170
rect 94976 296686 95096 296714
rect 93768 294024 93820 294030
rect 93768 293966 93820 293972
rect 93676 287156 93728 287162
rect 93676 287098 93728 287104
rect 93124 283620 93176 283626
rect 93124 283562 93176 283568
rect 93688 283506 93716 287098
rect 93780 286346 93808 293966
rect 93768 286340 93820 286346
rect 93768 286282 93820 286288
rect 94976 285569 95004 296686
rect 95160 292574 95188 378218
rect 95252 334626 95280 390374
rect 96586 390130 96614 390388
rect 96724 390374 97336 390402
rect 97552 390374 97888 390402
rect 96586 390102 96660 390130
rect 95884 388340 95936 388346
rect 95884 388282 95936 388288
rect 95240 334620 95292 334626
rect 95240 334562 95292 334568
rect 95896 293282 95924 388282
rect 96632 386374 96660 390102
rect 96620 386368 96672 386374
rect 96620 386310 96672 386316
rect 96724 382226 96752 390374
rect 96712 382220 96764 382226
rect 96712 382162 96764 382168
rect 96724 381614 96752 382162
rect 96712 381608 96764 381614
rect 96712 381550 96764 381556
rect 97552 376106 97580 390374
rect 98472 389337 98500 390646
rect 99196 389836 99248 389842
rect 99196 389778 99248 389784
rect 98458 389328 98514 389337
rect 98458 389263 98514 389272
rect 97908 386368 97960 386374
rect 97908 386310 97960 386316
rect 97814 385656 97870 385665
rect 97814 385591 97870 385600
rect 97540 376100 97592 376106
rect 97540 376042 97592 376048
rect 97828 338162 97856 385591
rect 97920 382974 97948 386310
rect 97908 382968 97960 382974
rect 97908 382910 97960 382916
rect 97998 381576 98054 381585
rect 97998 381511 98054 381520
rect 97908 377460 97960 377466
rect 97908 377402 97960 377408
rect 97816 338156 97868 338162
rect 97816 338098 97868 338104
rect 96528 323604 96580 323610
rect 96528 323546 96580 323552
rect 96436 305040 96488 305046
rect 96436 304982 96488 304988
rect 95884 293276 95936 293282
rect 95884 293218 95936 293224
rect 95068 292546 95188 292574
rect 95068 285705 95096 292546
rect 95240 288448 95292 288454
rect 95240 288390 95292 288396
rect 95252 287042 95280 288390
rect 95160 287014 95280 287042
rect 95054 285696 95110 285705
rect 95054 285631 95110 285640
rect 94134 285560 94190 285569
rect 94134 285495 94190 285504
rect 94962 285560 95018 285569
rect 94962 285495 95018 285504
rect 94148 284481 94176 285495
rect 94134 284472 94190 284481
rect 94134 284407 94190 284416
rect 94148 283506 94176 284407
rect 95068 283778 95096 285631
rect 94792 283750 95096 283778
rect 94792 283506 94820 283750
rect 95160 283506 95188 287014
rect 95608 285728 95660 285734
rect 95608 285670 95660 285676
rect 95620 283506 95648 285670
rect 91756 283478 92184 283506
rect 92736 283478 93072 283506
rect 93288 283478 93716 283506
rect 93840 283478 94176 283506
rect 94392 283478 94820 283506
rect 94944 283478 95188 283506
rect 95496 283478 95648 283506
rect 95698 283520 95754 283529
rect 96448 283506 96476 304982
rect 96540 288454 96568 323546
rect 97722 321056 97778 321065
rect 97722 320991 97778 321000
rect 96528 288448 96580 288454
rect 96528 288390 96580 288396
rect 97736 285569 97764 320991
rect 96710 285560 96766 285569
rect 96710 285495 96766 285504
rect 97722 285560 97778 285569
rect 97722 285495 97778 285504
rect 96724 284345 96752 285495
rect 96710 284336 96766 284345
rect 96710 284271 96766 284280
rect 96724 283506 96752 284271
rect 97828 283778 97856 338098
rect 97552 283750 97856 283778
rect 95754 283478 96476 283506
rect 96600 283478 96752 283506
rect 96802 283520 96858 283529
rect 95698 283455 95754 283464
rect 97552 283506 97580 283750
rect 97920 283506 97948 377402
rect 96858 283478 97580 283506
rect 97704 283490 97948 283506
rect 97704 283484 97960 283490
rect 97704 283478 97908 283484
rect 96802 283455 96858 283464
rect 97908 283426 97960 283432
rect 97920 283395 97948 283426
rect 91480 283206 91632 283234
rect 69204 283008 69256 283014
rect 69204 282950 69256 282956
rect 69756 283008 69808 283014
rect 69756 282950 69808 282956
rect 84752 283008 84804 283014
rect 84752 282950 84804 282956
rect 98012 282826 98040 381511
rect 98368 284980 98420 284986
rect 98368 284922 98420 284928
rect 98012 282798 98256 282826
rect 69018 282432 69074 282441
rect 69018 282367 69074 282376
rect 69032 282198 69060 282367
rect 69020 282192 69072 282198
rect 69020 282134 69072 282140
rect 98104 262177 98132 282798
rect 98380 281518 98408 284922
rect 98460 283484 98512 283490
rect 98460 283426 98512 283432
rect 98368 281512 98420 281518
rect 98368 281454 98420 281460
rect 98472 277394 98500 283426
rect 98624 282934 98960 282962
rect 98932 282878 98960 282934
rect 98920 282872 98972 282878
rect 98920 282814 98972 282820
rect 98472 277366 98776 277394
rect 98748 267073 98776 277366
rect 99208 273329 99236 389778
rect 99484 388385 99512 391002
rect 100666 390960 100722 390969
rect 100722 390932 100832 390946
rect 100722 390918 100846 390932
rect 100666 390895 100722 390904
rect 99760 390374 100096 390402
rect 99760 389065 99788 390374
rect 100818 390130 100846 390918
rect 105266 390416 105322 390425
rect 101384 390374 101720 390402
rect 100772 390102 100846 390130
rect 100772 389842 100800 390102
rect 100760 389836 100812 389842
rect 100760 389778 100812 389784
rect 101692 389162 101720 390374
rect 102106 390130 102134 390388
rect 102244 390374 102856 390402
rect 103592 390374 103744 390402
rect 102106 390102 102180 390130
rect 101680 389156 101732 389162
rect 101680 389098 101732 389104
rect 99746 389056 99802 389065
rect 99746 388991 99802 389000
rect 100114 389056 100170 389065
rect 100114 388991 100170 389000
rect 100024 388476 100076 388482
rect 100024 388418 100076 388424
rect 99470 388376 99526 388385
rect 99470 388311 99526 388320
rect 99288 329928 99340 329934
rect 99286 329896 99288 329905
rect 99340 329896 99342 329905
rect 99286 329831 99342 329840
rect 100036 299062 100064 388418
rect 100128 318170 100156 388991
rect 100666 388512 100722 388521
rect 100666 388447 100722 388456
rect 100680 328506 100708 388447
rect 102046 387152 102102 387161
rect 102046 387087 102102 387096
rect 101404 384396 101456 384402
rect 101404 384338 101456 384344
rect 100208 328500 100260 328506
rect 100208 328442 100260 328448
rect 100668 328500 100720 328506
rect 100668 328442 100720 328448
rect 100116 318164 100168 318170
rect 100116 318106 100168 318112
rect 100220 305046 100248 328442
rect 100668 306400 100720 306406
rect 100668 306342 100720 306348
rect 100208 305040 100260 305046
rect 100208 304982 100260 304988
rect 100116 301504 100168 301510
rect 100116 301446 100168 301452
rect 100024 299056 100076 299062
rect 100024 298998 100076 299004
rect 100022 285696 100078 285705
rect 100022 285631 100078 285640
rect 99472 283620 99524 283626
rect 99472 283562 99524 283568
rect 99380 282872 99432 282878
rect 99380 282814 99432 282820
rect 99392 280838 99420 282814
rect 99380 280832 99432 280838
rect 99380 280774 99432 280780
rect 99378 280256 99434 280265
rect 99378 280191 99434 280200
rect 99194 273320 99250 273329
rect 99194 273255 99250 273264
rect 99194 272096 99250 272105
rect 99194 272031 99250 272040
rect 98734 267064 98790 267073
rect 98734 266999 98790 267008
rect 98090 262168 98146 262177
rect 98090 262103 98146 262112
rect 98642 262168 98698 262177
rect 98642 262103 98698 262112
rect 98656 261089 98684 262103
rect 98642 261080 98698 261089
rect 98642 261015 98698 261024
rect 98090 259584 98146 259593
rect 98090 259519 98146 259528
rect 69020 242208 69072 242214
rect 69020 242150 69072 242156
rect 69032 241806 69060 242150
rect 69020 241800 69072 241806
rect 69020 241742 69072 241748
rect 69848 241800 69900 241806
rect 94780 241800 94832 241806
rect 69848 241742 69900 241748
rect 70122 241768 70178 241777
rect 69296 241732 69348 241738
rect 69296 241674 69348 241680
rect 68802 241369 68830 241604
rect 69124 241590 69184 241618
rect 68788 241360 68844 241369
rect 68788 241295 68844 241304
rect 69124 238746 69152 241590
rect 69112 238740 69164 238746
rect 69112 238682 69164 238688
rect 69124 237454 69152 238682
rect 69112 237448 69164 237454
rect 69112 237390 69164 237396
rect 68650 232656 68706 232665
rect 68650 232591 68706 232600
rect 68928 226364 68980 226370
rect 68928 226306 68980 226312
rect 68940 211138 68968 226306
rect 68468 211132 68520 211138
rect 68468 211074 68520 211080
rect 68928 211132 68980 211138
rect 68928 211074 68980 211080
rect 68284 193860 68336 193866
rect 68284 193802 68336 193808
rect 68296 136678 68324 193802
rect 68284 136672 68336 136678
rect 68284 136614 68336 136620
rect 67640 92880 67692 92886
rect 67640 92822 67692 92828
rect 67652 60042 67680 92822
rect 68480 92682 68508 211074
rect 68558 140856 68614 140865
rect 68558 140791 68614 140800
rect 68468 92676 68520 92682
rect 68468 92618 68520 92624
rect 68572 92449 68600 140791
rect 68652 134836 68704 134842
rect 68652 134778 68704 134784
rect 68664 113174 68692 134778
rect 69308 134722 69336 241674
rect 69400 241590 69736 241618
rect 69400 240145 69428 241590
rect 69386 240136 69442 240145
rect 69386 240071 69442 240080
rect 69860 238746 69888 241742
rect 71134 241768 71190 241777
rect 70178 241726 70288 241754
rect 70840 241726 71134 241754
rect 70122 241703 70178 241712
rect 72790 241768 72846 241777
rect 71134 241703 71190 241712
rect 72160 241726 72790 241754
rect 71056 241590 71392 241618
rect 71792 241604 71944 241618
rect 71792 241590 71958 241604
rect 70582 240816 70638 240825
rect 70582 240751 70638 240760
rect 70398 240136 70454 240145
rect 70398 240071 70454 240080
rect 70412 239873 70440 240071
rect 70398 239864 70454 239873
rect 70398 239799 70454 239808
rect 69848 238740 69900 238746
rect 69848 238682 69900 238688
rect 69664 237448 69716 237454
rect 69664 237390 69716 237396
rect 69676 220794 69704 237390
rect 70412 228410 70440 239799
rect 70400 228404 70452 228410
rect 70400 228346 70452 228352
rect 69664 220788 69716 220794
rect 69664 220730 69716 220736
rect 69676 134842 69704 220730
rect 70492 145580 70544 145586
rect 70492 145522 70544 145528
rect 69846 136912 69902 136921
rect 69846 136847 69902 136856
rect 69664 134836 69716 134842
rect 69664 134778 69716 134784
rect 69860 134722 69888 136847
rect 69940 136672 69992 136678
rect 69940 136614 69992 136620
rect 69000 134694 69336 134722
rect 69552 134694 69888 134722
rect 69952 134722 69980 136614
rect 69952 134694 70104 134722
rect 70504 134638 70532 145522
rect 70596 134994 70624 240751
rect 71056 240145 71084 241590
rect 71042 240136 71098 240145
rect 71042 240071 71098 240080
rect 71686 233880 71742 233889
rect 71686 233815 71742 233824
rect 71700 142154 71728 233815
rect 71792 226370 71820 241590
rect 71930 241466 71958 241590
rect 71918 241460 71970 241466
rect 71918 241402 71970 241408
rect 71964 232552 72016 232558
rect 71964 232494 72016 232500
rect 71780 226364 71832 226370
rect 71780 226306 71832 226312
rect 71780 220108 71832 220114
rect 71780 220050 71832 220056
rect 71424 142126 71728 142154
rect 70596 134966 70670 134994
rect 70642 134708 70670 134966
rect 71424 134722 71452 142126
rect 71688 140820 71740 140826
rect 71688 140762 71740 140768
rect 71700 134745 71728 140762
rect 71024 134694 71452 134722
rect 71686 134736 71742 134745
rect 71792 134722 71820 220050
rect 71976 140865 72004 232494
rect 71962 140856 72018 140865
rect 71962 140791 72018 140800
rect 72160 138145 72188 241726
rect 74262 241768 74318 241777
rect 74152 241726 74262 241754
rect 72790 241703 72846 241712
rect 74262 241703 74318 241712
rect 91558 241768 91614 241777
rect 91614 241726 92244 241754
rect 95882 241768 95938 241777
rect 94780 241742 94832 241748
rect 91558 241703 91614 241712
rect 72712 241590 73048 241618
rect 73264 241590 73600 241618
rect 72712 240009 72740 241590
rect 72422 240000 72478 240009
rect 72422 239935 72478 239944
rect 72698 240000 72754 240009
rect 72698 239935 72754 239944
rect 72436 230625 72464 239935
rect 73264 237386 73292 241590
rect 74276 238785 74304 241703
rect 74644 241590 74704 241618
rect 74920 241590 75256 241618
rect 75472 241590 75808 241618
rect 75932 241590 76360 241618
rect 76760 241604 76912 241618
rect 76760 241590 76926 241604
rect 74540 240168 74592 240174
rect 74540 240110 74592 240116
rect 74262 238776 74318 238785
rect 74262 238711 74318 238720
rect 74552 238678 74580 240110
rect 74644 240038 74672 241590
rect 74920 240174 74948 241590
rect 74908 240168 74960 240174
rect 74908 240110 74960 240116
rect 74632 240032 74684 240038
rect 74684 239980 74764 239986
rect 74632 239974 74764 239980
rect 74644 239958 74764 239974
rect 74630 238776 74686 238785
rect 74630 238711 74686 238720
rect 74540 238672 74592 238678
rect 74540 238614 74592 238620
rect 73252 237380 73304 237386
rect 73252 237322 73304 237328
rect 72792 233164 72844 233170
rect 72792 233106 72844 233112
rect 72804 232558 72832 233106
rect 72792 232552 72844 232558
rect 72792 232494 72844 232500
rect 72422 230616 72478 230625
rect 72422 230551 72478 230560
rect 72332 140072 72384 140078
rect 72332 140014 72384 140020
rect 72146 138136 72202 138145
rect 72146 138071 72202 138080
rect 72344 134722 72372 140014
rect 73160 137284 73212 137290
rect 73160 137226 73212 137232
rect 73172 134858 73200 137226
rect 73264 135969 73292 237322
rect 74552 234546 74580 238614
rect 74460 234518 74580 234546
rect 74460 216646 74488 234518
rect 74538 230616 74594 230625
rect 74538 230551 74594 230560
rect 73804 216640 73856 216646
rect 73804 216582 73856 216588
rect 74448 216640 74500 216646
rect 74448 216582 74500 216588
rect 73816 160750 73844 216582
rect 73804 160744 73856 160750
rect 73804 160686 73856 160692
rect 73344 148368 73396 148374
rect 73344 148310 73396 148316
rect 73250 135960 73306 135969
rect 73250 135895 73306 135904
rect 73172 134830 73246 134858
rect 71792 134694 72128 134722
rect 72344 134694 72680 134722
rect 73218 134708 73246 134830
rect 73356 134722 73384 148310
rect 74552 142866 74580 230551
rect 74540 142860 74592 142866
rect 74540 142802 74592 142808
rect 74644 138718 74672 238711
rect 74736 236774 74764 239958
rect 75472 238754 75500 241590
rect 74828 238726 75500 238754
rect 74724 236768 74776 236774
rect 74724 236710 74776 236716
rect 74828 233102 74856 238726
rect 75932 233170 75960 241590
rect 76104 236700 76156 236706
rect 76104 236642 76156 236648
rect 75920 233164 75972 233170
rect 75920 233106 75972 233112
rect 74816 233096 74868 233102
rect 74816 233038 74868 233044
rect 74828 229094 74856 233038
rect 74828 229066 75224 229094
rect 75196 155310 75224 229066
rect 75920 215960 75972 215966
rect 75920 215902 75972 215908
rect 75184 155304 75236 155310
rect 75184 155246 75236 155252
rect 74816 144288 74868 144294
rect 74816 144230 74868 144236
rect 74632 138712 74684 138718
rect 74632 138654 74684 138660
rect 73802 137320 73858 137329
rect 73802 137255 73858 137264
rect 73816 134722 73844 137255
rect 74724 136672 74776 136678
rect 74724 136614 74776 136620
rect 74736 134858 74764 136614
rect 74690 134830 74764 134858
rect 73356 134694 73600 134722
rect 73816 134694 74152 134722
rect 74690 134708 74718 134830
rect 74828 134722 74856 144230
rect 75932 138106 75960 215902
rect 76012 146124 76064 146130
rect 76012 146066 76064 146072
rect 75920 138100 75972 138106
rect 75920 138042 75972 138048
rect 75460 135176 75512 135182
rect 75460 135118 75512 135124
rect 75472 134722 75500 135118
rect 76024 134722 76052 146066
rect 76116 136678 76144 236642
rect 76656 233232 76708 233238
rect 76656 233174 76708 233180
rect 76562 225584 76618 225593
rect 76562 225519 76618 225528
rect 76576 140826 76604 225519
rect 76668 211818 76696 233174
rect 76760 224262 76788 241590
rect 76898 241505 76926 241590
rect 77450 241534 77478 241604
rect 78016 241590 78076 241618
rect 77438 241528 77490 241534
rect 76884 241496 76940 241505
rect 77438 241470 77490 241476
rect 76884 241431 76940 241440
rect 77450 241346 77478 241470
rect 77450 241318 77524 241346
rect 77300 240168 77352 240174
rect 77300 240110 77352 240116
rect 77312 235890 77340 240110
rect 77300 235884 77352 235890
rect 77300 235826 77352 235832
rect 77392 226296 77444 226302
rect 77392 226238 77444 226244
rect 76748 224256 76800 224262
rect 76748 224198 76800 224204
rect 76656 211812 76708 211818
rect 76656 211754 76708 211760
rect 76564 140820 76616 140826
rect 76564 140762 76616 140768
rect 76380 138100 76432 138106
rect 76380 138042 76432 138048
rect 76104 136672 76156 136678
rect 76104 136614 76156 136620
rect 76392 134722 76420 138042
rect 77404 134722 77432 226238
rect 77496 196654 77524 241318
rect 78048 240281 78076 241590
rect 78232 241590 78568 241618
rect 78692 241590 79120 241618
rect 79336 241590 79672 241618
rect 80164 241590 80224 241618
rect 80440 241590 80776 241618
rect 80992 241590 81328 241618
rect 81452 241590 81880 241618
rect 82004 241590 82432 241618
rect 82984 241590 83044 241618
rect 78034 240272 78090 240281
rect 78034 240207 78090 240216
rect 78232 240174 78260 241590
rect 78220 240168 78272 240174
rect 78220 240110 78272 240116
rect 78692 233238 78720 241590
rect 79336 238754 79364 241590
rect 80060 239488 80112 239494
rect 80060 239430 80112 239436
rect 78784 238726 79364 238754
rect 78784 234569 78812 238726
rect 80072 234598 80100 239430
rect 80164 238746 80192 241590
rect 80440 239494 80468 241590
rect 80428 239488 80480 239494
rect 80428 239430 80480 239436
rect 80992 238754 81020 241590
rect 80152 238740 80204 238746
rect 80152 238682 80204 238688
rect 80348 238726 81020 238754
rect 80164 237454 80192 238682
rect 80152 237448 80204 237454
rect 80152 237390 80204 237396
rect 80060 234592 80112 234598
rect 78770 234560 78826 234569
rect 80060 234534 80112 234540
rect 78770 234495 78826 234504
rect 78680 233232 78732 233238
rect 78680 233174 78732 233180
rect 77574 232656 77630 232665
rect 77574 232591 77630 232600
rect 77484 196648 77536 196654
rect 77484 196590 77536 196596
rect 74828 134694 75256 134722
rect 75472 134694 75808 134722
rect 76024 134694 76176 134722
rect 76392 134694 76728 134722
rect 77280 134694 77432 134722
rect 77588 134722 77616 232591
rect 78586 226944 78642 226953
rect 78586 226879 78642 226888
rect 78600 226302 78628 226879
rect 78588 226296 78640 226302
rect 78588 226238 78640 226244
rect 78784 140146 78812 234495
rect 80348 229838 80376 238726
rect 81452 237969 81480 241590
rect 82004 238754 82032 241590
rect 82082 240136 82138 240145
rect 82082 240071 82138 240080
rect 81544 238726 82032 238754
rect 81438 237960 81494 237969
rect 81438 237895 81494 237904
rect 80704 237448 80756 237454
rect 80704 237390 80756 237396
rect 80428 233980 80480 233986
rect 80428 233922 80480 233928
rect 80336 229832 80388 229838
rect 80336 229774 80388 229780
rect 79322 228304 79378 228313
rect 79322 228239 79378 228248
rect 78862 224224 78918 224233
rect 78862 224159 78918 224168
rect 78876 142154 78904 224159
rect 79336 146130 79364 228239
rect 80060 199436 80112 199442
rect 80060 199378 80112 199384
rect 79324 146124 79376 146130
rect 79324 146066 79376 146072
rect 78876 142126 79456 142154
rect 78772 140140 78824 140146
rect 78772 140082 78824 140088
rect 79324 138712 79376 138718
rect 79324 138654 79376 138660
rect 78496 137420 78548 137426
rect 78496 137362 78548 137368
rect 78508 134722 78536 137362
rect 79048 137284 79100 137290
rect 79048 137226 79100 137232
rect 79060 134722 79088 137226
rect 79336 134994 79364 138654
rect 77588 134694 77832 134722
rect 78200 134694 78536 134722
rect 78752 134694 79088 134722
rect 79290 134966 79364 134994
rect 79290 134708 79318 134966
rect 79428 134722 79456 142126
rect 80072 134722 80100 199378
rect 80440 137465 80468 233922
rect 80716 209098 80744 237390
rect 80980 233232 81032 233238
rect 80980 233174 81032 233180
rect 80992 233034 81020 233174
rect 80980 233028 81032 233034
rect 80980 232970 81032 232976
rect 81440 227996 81492 228002
rect 81440 227938 81492 227944
rect 80704 209092 80756 209098
rect 80704 209034 80756 209040
rect 81348 141500 81400 141506
rect 81348 141442 81400 141448
rect 81070 138680 81126 138689
rect 81070 138615 81126 138624
rect 80426 137456 80482 137465
rect 80426 137391 80428 137400
rect 80480 137391 80482 137400
rect 80428 137362 80480 137368
rect 80440 137331 80468 137362
rect 81084 134722 81112 138615
rect 81360 134994 81388 141442
rect 81452 138106 81480 227938
rect 81544 226137 81572 238726
rect 82096 227662 82124 240071
rect 83016 240038 83044 241590
rect 83200 241590 83536 241618
rect 83752 241590 84088 241618
rect 84640 241590 84700 241618
rect 83096 240168 83148 240174
rect 83096 240110 83148 240116
rect 83004 240032 83056 240038
rect 83004 239974 83056 239980
rect 82728 237448 82780 237454
rect 82728 237390 82780 237396
rect 82084 227656 82136 227662
rect 82084 227598 82136 227604
rect 81530 226128 81586 226137
rect 81530 226063 81586 226072
rect 82740 199578 82768 237390
rect 83108 206281 83136 240110
rect 83200 238746 83228 241590
rect 83752 240174 83780 241590
rect 84672 240854 84700 241590
rect 84764 241590 85192 241618
rect 85684 241590 85744 241618
rect 85960 241590 86296 241618
rect 86848 241590 86908 241618
rect 84660 240848 84712 240854
rect 84660 240790 84712 240796
rect 83740 240168 83792 240174
rect 83740 240110 83792 240116
rect 84016 240032 84068 240038
rect 84016 239974 84068 239980
rect 83188 238740 83240 238746
rect 83188 238682 83240 238688
rect 83200 237454 83228 238682
rect 83188 237448 83240 237454
rect 83188 237390 83240 237396
rect 84028 210361 84056 239974
rect 84764 238754 84792 241590
rect 85580 240168 85632 240174
rect 85580 240110 85632 240116
rect 85486 240000 85542 240009
rect 85486 239935 85542 239944
rect 84212 238726 84792 238754
rect 84108 235272 84160 235278
rect 84108 235214 84160 235220
rect 84014 210352 84070 210361
rect 84014 210287 84070 210296
rect 83094 206272 83150 206281
rect 83094 206207 83150 206216
rect 82912 203584 82964 203590
rect 82912 203526 82964 203532
rect 82728 199572 82780 199578
rect 82728 199514 82780 199520
rect 81532 180872 81584 180878
rect 81532 180814 81584 180820
rect 81440 138100 81492 138106
rect 81440 138042 81492 138048
rect 79428 134694 79856 134722
rect 80072 134694 80408 134722
rect 80776 134694 81112 134722
rect 81314 134966 81388 134994
rect 81314 134708 81342 134966
rect 81544 134722 81572 180814
rect 82924 151814 82952 203526
rect 84120 156738 84148 235214
rect 84212 207641 84240 238726
rect 84844 214600 84896 214606
rect 84844 214542 84896 214548
rect 84198 207632 84254 207641
rect 84198 207567 84254 207576
rect 84856 180878 84884 214542
rect 84844 180872 84896 180878
rect 84844 180814 84896 180820
rect 84108 156732 84160 156738
rect 84108 156674 84160 156680
rect 82924 151786 83780 151814
rect 82820 142180 82872 142186
rect 82820 142122 82872 142128
rect 82084 138100 82136 138106
rect 82084 138042 82136 138048
rect 82096 134722 82124 138042
rect 82832 134994 82860 142122
rect 83648 136672 83700 136678
rect 83648 136614 83700 136620
rect 82786 134966 82860 134994
rect 81544 134694 81880 134722
rect 82096 134694 82432 134722
rect 82786 134708 82814 134966
rect 83660 134722 83688 136614
rect 83352 134694 83688 134722
rect 83752 134722 83780 151786
rect 84568 147688 84620 147694
rect 84568 147630 84620 147636
rect 84108 145580 84160 145586
rect 84108 145522 84160 145528
rect 84120 136678 84148 145522
rect 84474 141400 84530 141409
rect 84474 141335 84530 141344
rect 84108 136672 84160 136678
rect 84108 136614 84160 136620
rect 84488 134994 84516 141335
rect 84442 134966 84516 134994
rect 83752 134694 83904 134722
rect 84442 134708 84470 134966
rect 84580 134722 84608 147630
rect 85500 142866 85528 239935
rect 85592 231305 85620 240110
rect 85684 233345 85712 241590
rect 85960 240174 85988 241590
rect 85948 240168 86000 240174
rect 85948 240110 86000 240116
rect 86880 240009 86908 241590
rect 87064 241590 87400 241618
rect 87524 241590 87952 241618
rect 88444 241590 88504 241618
rect 88720 241590 89056 241618
rect 89608 241590 89668 241618
rect 87064 240106 87092 241590
rect 87052 240100 87104 240106
rect 87052 240042 87104 240048
rect 86866 240000 86922 240009
rect 86866 239935 86922 239944
rect 87524 238754 87552 241590
rect 88156 240780 88208 240786
rect 88156 240722 88208 240728
rect 87064 238726 87552 238754
rect 87064 238134 87092 238726
rect 88064 238672 88116 238678
rect 88064 238614 88116 238620
rect 88076 238134 88104 238614
rect 87052 238128 87104 238134
rect 87052 238070 87104 238076
rect 88064 238128 88116 238134
rect 88064 238070 88116 238076
rect 86774 234152 86830 234161
rect 86774 234087 86830 234096
rect 86788 233345 86816 234087
rect 85670 233336 85726 233345
rect 85670 233271 85726 233280
rect 86774 233336 86830 233345
rect 86774 233271 86830 233280
rect 85578 231296 85634 231305
rect 85578 231231 85634 231240
rect 85578 231160 85634 231169
rect 85578 231095 85634 231104
rect 85592 228002 85620 231095
rect 85580 227996 85632 228002
rect 85580 227938 85632 227944
rect 86222 213208 86278 213217
rect 86222 213143 86278 213152
rect 85580 191208 85632 191214
rect 85580 191150 85632 191156
rect 85592 151814 85620 191150
rect 85592 151786 86080 151814
rect 85488 142860 85540 142866
rect 85488 142802 85540 142808
rect 85488 139460 85540 139466
rect 85488 139402 85540 139408
rect 85500 134722 85528 139402
rect 85948 136672 86000 136678
rect 85948 136614 86000 136620
rect 85960 134994 85988 136614
rect 84580 134694 85008 134722
rect 85376 134694 85528 134722
rect 85914 134966 85988 134994
rect 85914 134708 85942 134966
rect 86052 134722 86080 151786
rect 86236 142186 86264 213143
rect 86788 193866 86816 233271
rect 86868 222896 86920 222902
rect 86868 222838 86920 222844
rect 86776 193860 86828 193866
rect 86776 193802 86828 193808
rect 86224 142180 86276 142186
rect 86224 142122 86276 142128
rect 86880 137329 86908 222838
rect 88076 211818 88104 238070
rect 88168 237386 88196 240722
rect 88340 240168 88392 240174
rect 88340 240110 88392 240116
rect 88156 237380 88208 237386
rect 88156 237322 88208 237328
rect 88064 211812 88116 211818
rect 88064 211754 88116 211760
rect 88168 199442 88196 237322
rect 88352 235385 88380 240110
rect 88338 235376 88394 235385
rect 88338 235311 88394 235320
rect 88340 227792 88392 227798
rect 88340 227734 88392 227740
rect 88248 225684 88300 225690
rect 88248 225626 88300 225632
rect 88156 199436 88208 199442
rect 88156 199378 88208 199384
rect 88156 198008 88208 198014
rect 88156 197950 88208 197956
rect 88064 196648 88116 196654
rect 88064 196590 88116 196596
rect 88076 142154 88104 196590
rect 87800 142126 88104 142154
rect 86866 137320 86922 137329
rect 86866 137255 86868 137264
rect 86920 137255 86922 137264
rect 86868 137226 86920 137232
rect 86880 137195 86908 137226
rect 87326 136776 87382 136785
rect 87326 136711 87382 136720
rect 87340 134722 87368 136711
rect 87800 134722 87828 142126
rect 88168 141522 88196 197950
rect 88260 142186 88288 225626
rect 88352 151814 88380 227734
rect 88444 224942 88472 241590
rect 88720 240174 88748 241590
rect 88708 240168 88760 240174
rect 88708 240110 88760 240116
rect 89640 239426 89668 241590
rect 89732 241590 90160 241618
rect 90712 241590 91048 241618
rect 89628 239420 89680 239426
rect 89628 239362 89680 239368
rect 89732 237153 89760 241590
rect 90914 237416 90970 237425
rect 90914 237351 90970 237360
rect 89718 237144 89774 237153
rect 89718 237079 89774 237088
rect 89168 236768 89220 236774
rect 89168 236710 89220 236716
rect 88432 224936 88484 224942
rect 88432 224878 88484 224884
rect 88984 214668 89036 214674
rect 88984 214610 89036 214616
rect 88352 151786 88932 151814
rect 88248 142180 88300 142186
rect 88248 142122 88300 142128
rect 88076 141494 88196 141522
rect 88076 137358 88104 141494
rect 88156 141432 88208 141438
rect 88156 141374 88208 141380
rect 88168 140758 88196 141374
rect 88156 140752 88208 140758
rect 88156 140694 88208 140700
rect 88064 137352 88116 137358
rect 88064 137294 88116 137300
rect 88076 136678 88104 137294
rect 88064 136672 88116 136678
rect 88064 136614 88116 136620
rect 88168 134722 88196 140694
rect 88260 139398 88288 142122
rect 88798 140040 88854 140049
rect 88798 139975 88854 139984
rect 88248 139392 88300 139398
rect 88248 139334 88300 139340
rect 88812 134722 88840 139975
rect 88904 138122 88932 151786
rect 88996 139466 89024 214610
rect 89076 156664 89128 156670
rect 89076 156606 89128 156612
rect 89088 147694 89116 156606
rect 89180 151814 89208 236710
rect 89732 235278 89760 237079
rect 90824 236020 90876 236026
rect 90824 235962 90876 235968
rect 89720 235272 89772 235278
rect 89720 235214 89772 235220
rect 89720 224188 89772 224194
rect 89720 224130 89772 224136
rect 89180 151786 89300 151814
rect 89076 147688 89128 147694
rect 89076 147630 89128 147636
rect 88984 139460 89036 139466
rect 88984 139402 89036 139408
rect 88904 138094 89208 138122
rect 89076 137284 89128 137290
rect 89076 137226 89128 137232
rect 89088 134858 89116 137226
rect 86052 134694 86480 134722
rect 87032 134694 87368 134722
rect 87584 134694 87828 134722
rect 87952 134694 88196 134722
rect 88504 134694 88840 134722
rect 89042 134830 89116 134858
rect 89042 134708 89070 134830
rect 89180 134722 89208 138094
rect 89272 134842 89300 151786
rect 89732 138106 89760 224130
rect 90836 211857 90864 235962
rect 90822 211848 90878 211857
rect 90822 211783 90878 211792
rect 90928 206417 90956 237351
rect 90914 206408 90970 206417
rect 90914 206343 90970 206352
rect 91020 204950 91048 241590
rect 91204 241590 91264 241618
rect 91100 240168 91152 240174
rect 91100 240110 91152 240116
rect 91112 236026 91140 240110
rect 91204 237425 91232 241590
rect 92216 238754 92244 241726
rect 92308 241590 92368 241618
rect 92492 241590 92920 241618
rect 93044 241590 93472 241618
rect 94024 241590 94084 241618
rect 92308 240174 92336 241590
rect 92296 240168 92348 240174
rect 92296 240110 92348 240116
rect 92216 238726 92336 238754
rect 91190 237416 91246 237425
rect 91190 237351 91246 237360
rect 91100 236020 91152 236026
rect 91100 235962 91152 235968
rect 92204 227860 92256 227866
rect 92204 227802 92256 227808
rect 92216 209166 92244 227802
rect 92308 227769 92336 238726
rect 92388 229832 92440 229838
rect 92388 229774 92440 229780
rect 92294 227760 92350 227769
rect 92294 227695 92350 227704
rect 92294 227080 92350 227089
rect 92294 227015 92350 227024
rect 92204 209160 92256 209166
rect 92204 209102 92256 209108
rect 91008 204944 91060 204950
rect 91008 204886 91060 204892
rect 90364 199572 90416 199578
rect 90364 199514 90416 199520
rect 89812 199504 89864 199510
rect 89812 199446 89864 199452
rect 89720 138100 89772 138106
rect 89720 138042 89772 138048
rect 89260 134836 89312 134842
rect 89260 134778 89312 134784
rect 89824 134722 89852 199446
rect 90180 138100 90232 138106
rect 90180 138042 90232 138048
rect 90192 134722 90220 138042
rect 90376 134842 90404 199514
rect 91008 140072 91060 140078
rect 91008 140014 91060 140020
rect 91020 135930 91048 140014
rect 91008 135924 91060 135930
rect 91008 135866 91060 135872
rect 91284 135924 91336 135930
rect 91284 135866 91336 135872
rect 91192 135856 91244 135862
rect 91192 135798 91244 135804
rect 91204 135318 91232 135798
rect 91192 135312 91244 135318
rect 91192 135254 91244 135260
rect 90364 134836 90416 134842
rect 90364 134778 90416 134784
rect 91204 134722 91232 135254
rect 89180 134694 89608 134722
rect 89824 134694 89976 134722
rect 90192 134694 90528 134722
rect 91080 134694 91232 134722
rect 91296 134722 91324 135866
rect 92308 135318 92336 227015
rect 92296 135312 92348 135318
rect 92400 135289 92428 229774
rect 92492 220697 92520 241590
rect 93044 238754 93072 241590
rect 93860 240100 93912 240106
rect 93860 240042 93912 240048
rect 92584 238726 93072 238754
rect 92584 237386 92612 238726
rect 92572 237380 92624 237386
rect 92572 237322 92624 237328
rect 93124 236700 93176 236706
rect 93124 236642 93176 236648
rect 92662 235512 92718 235521
rect 92662 235447 92718 235456
rect 92478 220688 92534 220697
rect 92478 220623 92534 220632
rect 92478 148336 92534 148345
rect 92478 148271 92534 148280
rect 92296 135254 92348 135260
rect 92386 135280 92442 135289
rect 92308 134722 92336 135254
rect 92386 135215 92442 135224
rect 92492 134994 92520 148271
rect 92492 134966 92566 134994
rect 91296 134694 91632 134722
rect 92184 134694 92336 134722
rect 92538 134708 92566 134966
rect 92676 134722 92704 235447
rect 93136 227798 93164 236642
rect 93872 234546 93900 240042
rect 94056 235550 94084 241590
rect 94240 241590 94576 241618
rect 94240 240106 94268 241590
rect 94228 240100 94280 240106
rect 94228 240042 94280 240048
rect 94044 235544 94096 235550
rect 94044 235486 94096 235492
rect 94504 235544 94556 235550
rect 94504 235486 94556 235492
rect 93780 234518 93900 234546
rect 93124 227792 93176 227798
rect 93124 227734 93176 227740
rect 93780 207777 93808 234518
rect 93858 233880 93914 233889
rect 93858 233815 93914 233824
rect 93766 207768 93822 207777
rect 93766 207703 93822 207712
rect 92754 200696 92810 200705
rect 92754 200631 92810 200640
rect 92768 151814 92796 200631
rect 92768 151786 93256 151814
rect 93228 134722 93256 151786
rect 93872 134722 93900 233815
rect 94516 227798 94544 235486
rect 94504 227792 94556 227798
rect 94504 227734 94556 227740
rect 94686 227760 94742 227769
rect 94686 227695 94742 227704
rect 94596 138780 94648 138786
rect 94596 138722 94648 138728
rect 94608 134994 94636 138722
rect 94562 134966 94636 134994
rect 92676 134694 93104 134722
rect 93228 134694 93656 134722
rect 93872 134694 94208 134722
rect 94562 134708 94590 134966
rect 71686 134671 71742 134680
rect 70492 134632 70544 134638
rect 70492 134574 70544 134580
rect 71228 134632 71280 134638
rect 71280 134580 71576 134586
rect 71228 134574 71576 134580
rect 71240 134558 71576 134574
rect 94700 124166 94728 227695
rect 94792 224194 94820 241742
rect 95252 241726 95882 241754
rect 94962 241632 95018 241641
rect 95018 241604 95128 241618
rect 95018 241590 95142 241604
rect 94962 241567 95018 241576
rect 95114 241482 95142 241590
rect 95114 241454 95188 241482
rect 95160 227730 95188 241454
rect 95148 227724 95200 227730
rect 95148 227666 95200 227672
rect 94780 224188 94832 224194
rect 94780 224130 94832 224136
rect 94780 142860 94832 142866
rect 94780 142802 94832 142808
rect 94792 135250 94820 142802
rect 94962 137456 95018 137465
rect 94962 137391 95018 137400
rect 94780 135244 94832 135250
rect 94780 135186 94832 135192
rect 94872 134768 94924 134774
rect 94872 134710 94924 134716
rect 94884 134609 94912 134710
rect 94870 134600 94926 134609
rect 94870 134535 94926 134544
rect 94976 133210 95004 137391
rect 94964 133204 95016 133210
rect 94964 133146 95016 133152
rect 94688 124160 94740 124166
rect 94688 124102 94740 124108
rect 95148 124160 95200 124166
rect 95252 124137 95280 241726
rect 95882 241703 95938 241712
rect 95896 241590 96232 241618
rect 96724 241590 96784 241618
rect 97000 241590 97336 241618
rect 97828 241590 97888 241618
rect 95896 238754 95924 241590
rect 96620 240168 96672 240174
rect 96620 240110 96672 240116
rect 95344 238726 95924 238754
rect 95344 216753 95372 238726
rect 95976 227792 96028 227798
rect 95976 227734 96028 227740
rect 95882 217288 95938 217297
rect 95882 217223 95938 217232
rect 95896 216753 95924 217223
rect 95330 216744 95386 216753
rect 95330 216679 95386 216688
rect 95882 216744 95938 216753
rect 95882 216679 95938 216688
rect 95148 124102 95200 124108
rect 95238 124128 95294 124137
rect 95160 122754 95188 124102
rect 95238 124063 95294 124072
rect 95160 122726 95280 122754
rect 68664 113146 68968 113174
rect 68940 93514 68968 113146
rect 94780 104780 94832 104786
rect 94780 104722 94832 104728
rect 94688 93560 94740 93566
rect 68940 93486 69184 93514
rect 94392 93508 94688 93514
rect 94392 93502 94740 93508
rect 94392 93486 94728 93502
rect 68652 92880 68704 92886
rect 68704 92828 68816 92834
rect 68652 92822 68816 92828
rect 68664 92806 68816 92822
rect 69722 92721 69750 92820
rect 69570 92712 69626 92721
rect 69570 92647 69626 92656
rect 69708 92712 69764 92721
rect 70274 92698 70302 92820
rect 70274 92670 70348 92698
rect 70826 92687 70854 92820
rect 69708 92647 69764 92656
rect 69584 92562 69612 92647
rect 70320 92585 70348 92670
rect 70812 92678 70868 92687
rect 70812 92613 70868 92622
rect 70306 92576 70362 92585
rect 69584 92534 69888 92562
rect 68558 92440 68614 92449
rect 68558 92375 68614 92384
rect 69860 84153 69888 92534
rect 71194 92562 71222 92820
rect 71746 92682 71774 92820
rect 71734 92676 71786 92682
rect 71734 92618 71786 92624
rect 72298 92562 72326 92820
rect 72850 92750 72878 92820
rect 72838 92744 72890 92750
rect 72838 92686 72890 92692
rect 73402 92562 73430 92820
rect 70306 92511 70362 92520
rect 71148 92534 71222 92562
rect 72252 92534 72326 92562
rect 73356 92534 73430 92562
rect 73770 92562 73798 92820
rect 74322 92562 74350 92820
rect 74874 92562 74902 92820
rect 75426 92562 75454 92820
rect 75794 92562 75822 92820
rect 76346 92562 76374 92820
rect 76898 92562 76926 92820
rect 73770 92534 73844 92562
rect 74322 92534 74396 92562
rect 70320 84194 70348 92511
rect 71148 90953 71176 92534
rect 72252 91089 72280 92534
rect 73356 92410 73384 92534
rect 73344 92404 73396 92410
rect 73344 92346 73396 92352
rect 72238 91080 72294 91089
rect 72238 91015 72294 91024
rect 71134 90944 71190 90953
rect 71134 90879 71190 90888
rect 73816 88262 73844 92534
rect 74368 90778 74396 92534
rect 74828 92534 74902 92562
rect 75380 92534 75454 92562
rect 75748 92534 75822 92562
rect 76300 92534 76374 92562
rect 76852 92534 76926 92562
rect 77450 92562 77478 92820
rect 78002 92562 78030 92820
rect 78370 92562 78398 92820
rect 78922 92562 78950 92820
rect 77450 92534 77524 92562
rect 74356 90772 74408 90778
rect 74356 90714 74408 90720
rect 73804 88256 73856 88262
rect 74828 88233 74856 92534
rect 75276 90772 75328 90778
rect 75276 90714 75328 90720
rect 73804 88198 73856 88204
rect 74814 88224 74870 88233
rect 70228 84166 70348 84194
rect 69846 84144 69902 84153
rect 69846 84079 69902 84088
rect 68928 64184 68980 64190
rect 68928 64126 68980 64132
rect 67640 60036 67692 60042
rect 67640 59978 67692 59984
rect 67548 56568 67600 56574
rect 67548 56510 67600 56516
rect 67546 47560 67602 47569
rect 67546 47495 67602 47504
rect 67560 3534 67588 47495
rect 68940 3534 68968 64126
rect 70228 62830 70256 84166
rect 70308 68332 70360 68338
rect 70308 68274 70360 68280
rect 70216 62824 70268 62830
rect 70216 62766 70268 62772
rect 70214 11656 70270 11665
rect 70214 11591 70270 11600
rect 70228 3534 70256 11591
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 65524 3188 65576 3194
rect 65524 3130 65576 3136
rect 66076 3188 66128 3194
rect 66076 3130 66128 3136
rect 65536 480 65564 3130
rect 66732 480 66760 3470
rect 67928 480 67956 3470
rect 69124 480 69152 3470
rect 70320 480 70348 68274
rect 72424 61396 72476 61402
rect 72424 61338 72476 61344
rect 71688 57316 71740 57322
rect 71688 57258 71740 57264
rect 71700 6914 71728 57258
rect 72436 20670 72464 61338
rect 73816 49026 73844 88198
rect 74814 88159 74870 88168
rect 75184 86896 75236 86902
rect 75184 86838 75236 86844
rect 75196 53106 75224 86838
rect 75288 78674 75316 90714
rect 75380 86902 75408 92534
rect 75748 92449 75776 92534
rect 75734 92440 75790 92449
rect 75734 92375 75790 92384
rect 76300 89622 76328 92534
rect 76288 89616 76340 89622
rect 76288 89558 76340 89564
rect 76852 88330 76880 92534
rect 77496 90681 77524 92534
rect 77956 92534 78030 92562
rect 78324 92534 78398 92562
rect 78692 92534 78950 92562
rect 79474 92562 79502 92820
rect 80026 92562 80054 92820
rect 80578 92562 80606 92820
rect 80946 92562 80974 92820
rect 81498 92562 81526 92820
rect 79474 92534 79548 92562
rect 80026 92534 80100 92562
rect 80578 92534 80652 92562
rect 80946 92534 81020 92562
rect 77956 90817 77984 92534
rect 77942 90808 77998 90817
rect 77942 90743 77998 90752
rect 77482 90672 77538 90681
rect 77482 90607 77538 90616
rect 78324 89690 78352 92534
rect 78312 89684 78364 89690
rect 78312 89626 78364 89632
rect 76564 88324 76616 88330
rect 76564 88266 76616 88272
rect 76840 88324 76892 88330
rect 76840 88266 76892 88272
rect 75368 86896 75420 86902
rect 75368 86838 75420 86844
rect 75276 78668 75328 78674
rect 75276 78610 75328 78616
rect 75184 53100 75236 53106
rect 75184 53042 75236 53048
rect 75828 51740 75880 51746
rect 75828 51682 75880 51688
rect 73804 49020 73856 49026
rect 73804 48962 73856 48968
rect 74446 28248 74502 28257
rect 74446 28183 74502 28192
rect 72514 25528 72570 25537
rect 72514 25463 72570 25472
rect 72424 20664 72476 20670
rect 72424 20606 72476 20612
rect 71516 6886 71728 6914
rect 71516 480 71544 6886
rect 72528 3602 72556 25463
rect 72516 3596 72568 3602
rect 72516 3538 72568 3544
rect 74460 3534 74488 28183
rect 75840 3534 75868 51682
rect 76576 46238 76604 88266
rect 78692 84182 78720 92534
rect 79520 85513 79548 92534
rect 80072 88330 80100 92534
rect 80624 90817 80652 92534
rect 80610 90808 80666 90817
rect 80610 90743 80666 90752
rect 80992 89758 81020 92534
rect 81452 92534 81526 92562
rect 82050 92562 82078 92820
rect 82602 92562 82630 92820
rect 82970 92562 82998 92820
rect 83522 92562 83550 92820
rect 84074 92562 84102 92820
rect 84626 92562 84654 92820
rect 85178 92562 85206 92820
rect 85546 92562 85574 92820
rect 86098 92562 86126 92820
rect 82050 92534 82124 92562
rect 82602 92534 82676 92562
rect 82970 92534 83044 92562
rect 83522 92534 83596 92562
rect 84074 92534 84148 92562
rect 84626 92534 84700 92562
rect 85178 92534 85252 92562
rect 85546 92534 85620 92562
rect 81452 90953 81480 92534
rect 81438 90944 81494 90953
rect 81438 90879 81494 90888
rect 80980 89752 81032 89758
rect 82096 89729 82124 92534
rect 82648 89962 82676 92534
rect 82636 89956 82688 89962
rect 82636 89898 82688 89904
rect 80980 89694 81032 89700
rect 82082 89720 82138 89729
rect 82082 89655 82138 89664
rect 80060 88324 80112 88330
rect 80060 88266 80112 88272
rect 83016 88097 83044 92534
rect 83464 89752 83516 89758
rect 83464 89694 83516 89700
rect 83002 88088 83058 88097
rect 83002 88023 83058 88032
rect 79506 85504 79562 85513
rect 79506 85439 79562 85448
rect 78680 84176 78732 84182
rect 78680 84118 78732 84124
rect 78692 82890 78720 84118
rect 78680 82884 78732 82890
rect 78680 82826 78732 82832
rect 79324 82884 79376 82890
rect 79324 82826 79376 82832
rect 77206 73808 77262 73817
rect 77206 73743 77262 73752
rect 76564 46232 76616 46238
rect 76564 46174 76616 46180
rect 77220 3534 77248 73743
rect 79336 69698 79364 82826
rect 83476 82822 83504 89694
rect 83568 85377 83596 92534
rect 84120 89622 84148 92534
rect 84108 89616 84160 89622
rect 84108 89558 84160 89564
rect 84672 86873 84700 92534
rect 85224 89758 85252 92534
rect 85212 89752 85264 89758
rect 85212 89694 85264 89700
rect 84658 86864 84714 86873
rect 84658 86799 84714 86808
rect 83554 85368 83610 85377
rect 83554 85303 83610 85312
rect 85592 84114 85620 92534
rect 86052 92534 86126 92562
rect 86650 92562 86678 92820
rect 87202 92562 87230 92820
rect 87570 92698 87598 92820
rect 87570 92670 87644 92698
rect 86650 92534 86724 92562
rect 87202 92534 87276 92562
rect 86052 92478 86080 92534
rect 86040 92472 86092 92478
rect 86040 92414 86092 92420
rect 86696 92410 86724 92534
rect 86684 92404 86736 92410
rect 86684 92346 86736 92352
rect 86868 89956 86920 89962
rect 86868 89898 86920 89904
rect 86880 85542 86908 89898
rect 87248 88262 87276 92534
rect 87616 90574 87644 92670
rect 88122 92562 88150 92820
rect 88674 92562 88702 92820
rect 89226 92562 89254 92820
rect 89778 92562 89806 92820
rect 90146 92562 90174 92820
rect 90698 92562 90726 92820
rect 91250 92698 91278 92820
rect 91802 92750 91830 92820
rect 91790 92744 91842 92750
rect 91250 92670 91324 92698
rect 91790 92686 91842 92692
rect 88122 92534 88196 92562
rect 88674 92534 88748 92562
rect 89226 92534 89300 92562
rect 89778 92534 89852 92562
rect 90146 92534 90220 92562
rect 90698 92534 90772 92562
rect 87604 90568 87656 90574
rect 87604 90510 87656 90516
rect 87236 88256 87288 88262
rect 87236 88198 87288 88204
rect 88168 86902 88196 92534
rect 88248 90908 88300 90914
rect 88248 90850 88300 90856
rect 88260 90574 88288 90850
rect 88248 90568 88300 90574
rect 88248 90510 88300 90516
rect 88156 86896 88208 86902
rect 88156 86838 88208 86844
rect 86868 85536 86920 85542
rect 86868 85478 86920 85484
rect 85580 84108 85632 84114
rect 85580 84050 85632 84056
rect 86776 84108 86828 84114
rect 86776 84050 86828 84056
rect 83464 82816 83516 82822
rect 83464 82758 83516 82764
rect 84108 82816 84160 82822
rect 84108 82758 84160 82764
rect 79968 75200 80020 75206
rect 79968 75142 80020 75148
rect 79324 69692 79376 69698
rect 79324 69634 79376 69640
rect 78588 20052 78640 20058
rect 78588 19994 78640 20000
rect 77390 4856 77446 4865
rect 77390 4791 77446 4800
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 72608 3460 72660 3466
rect 72608 3402 72660 3408
rect 72620 480 72648 3402
rect 73816 480 73844 3470
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77404 480 77432 4791
rect 78600 480 78628 19994
rect 79980 6914 80008 75142
rect 83462 72448 83518 72457
rect 83462 72383 83518 72392
rect 82728 32428 82780 32434
rect 82728 32370 82780 32376
rect 79704 6886 80008 6914
rect 79704 480 79732 6886
rect 82740 3534 82768 32370
rect 83280 6180 83332 6186
rect 83280 6122 83332 6128
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 80888 3188 80940 3194
rect 80888 3130 80940 3136
rect 80900 480 80928 3130
rect 82096 480 82124 3470
rect 83292 480 83320 6122
rect 83476 3194 83504 72383
rect 84120 43450 84148 82758
rect 86788 58682 86816 84050
rect 86776 58676 86828 58682
rect 86776 58618 86828 58624
rect 84108 43444 84160 43450
rect 84108 43386 84160 43392
rect 85486 29608 85542 29617
rect 85486 29543 85542 29552
rect 85500 3534 85528 29543
rect 86880 15910 86908 85478
rect 87602 76528 87658 76537
rect 87602 76463 87658 76472
rect 86868 15904 86920 15910
rect 86868 15846 86920 15852
rect 87616 3534 87644 76463
rect 88168 54534 88196 86838
rect 88156 54528 88208 54534
rect 88156 54470 88208 54476
rect 88260 42090 88288 90510
rect 88720 88233 88748 92534
rect 89272 92478 89300 92534
rect 89260 92472 89312 92478
rect 89260 92414 89312 92420
rect 89824 92313 89852 92534
rect 89810 92304 89866 92313
rect 89810 92239 89866 92248
rect 90192 91050 90220 92534
rect 90180 91044 90232 91050
rect 90180 90986 90232 90992
rect 90744 90953 90772 92534
rect 91296 92449 91324 92670
rect 92354 92562 92382 92820
rect 92722 92698 92750 92820
rect 92722 92670 92796 92698
rect 92354 92534 92428 92562
rect 91282 92440 91338 92449
rect 91282 92375 91338 92384
rect 90730 90944 90786 90953
rect 90730 90879 90786 90888
rect 89536 89752 89588 89758
rect 89536 89694 89588 89700
rect 89548 89593 89576 89694
rect 92400 89690 92428 92534
rect 92570 91488 92626 91497
rect 92570 91423 92626 91432
rect 92584 90681 92612 91423
rect 92768 91089 92796 92670
rect 93274 92562 93302 92820
rect 93826 92698 93854 92820
rect 94792 92750 94820 104722
rect 95146 94344 95202 94353
rect 95146 94279 95202 94288
rect 95056 93152 95108 93158
rect 95056 93094 95108 93100
rect 94780 92744 94832 92750
rect 93826 92670 93900 92698
rect 94780 92686 94832 92692
rect 92952 92534 93302 92562
rect 92754 91080 92810 91089
rect 92754 91015 92810 91024
rect 92570 90672 92626 90681
rect 92570 90607 92626 90616
rect 92388 89684 92440 89690
rect 92388 89626 92440 89632
rect 89534 89584 89590 89593
rect 89590 89542 89668 89570
rect 89534 89519 89590 89528
rect 88706 88224 88762 88233
rect 88706 88159 88762 88168
rect 89534 88224 89590 88233
rect 89534 88159 89590 88168
rect 89548 87961 89576 88159
rect 89534 87952 89590 87961
rect 89534 87887 89590 87896
rect 89548 50386 89576 87887
rect 89536 50380 89588 50386
rect 89536 50322 89588 50328
rect 88248 42084 88300 42090
rect 88248 42026 88300 42032
rect 88984 26920 89036 26926
rect 88984 26862 89036 26868
rect 88248 18692 88300 18698
rect 88248 18634 88300 18640
rect 88260 6914 88288 18634
rect 87984 6886 88288 6914
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 86868 3528 86920 3534
rect 85488 3470 85540 3476
rect 85670 3496 85726 3505
rect 83464 3188 83516 3194
rect 83464 3130 83516 3136
rect 84488 480 84516 3470
rect 86868 3470 86920 3476
rect 87604 3528 87656 3534
rect 87604 3470 87656 3476
rect 85670 3431 85726 3440
rect 85684 480 85712 3431
rect 86880 480 86908 3470
rect 87984 480 88012 6886
rect 88996 3369 89024 26862
rect 89536 13184 89588 13190
rect 89536 13126 89588 13132
rect 88982 3360 89038 3369
rect 88982 3295 89038 3304
rect 89180 598 89392 626
rect 89180 480 89208 598
rect 89364 490 89392 598
rect 89548 490 89576 13126
rect 89640 11014 89668 89542
rect 92952 84194 92980 92534
rect 93872 92449 93900 92670
rect 93858 92440 93914 92449
rect 93858 92375 93914 92384
rect 95068 91497 95096 93094
rect 95054 91488 95110 91497
rect 95054 91423 95110 91432
rect 92492 84182 92980 84194
rect 92480 84176 92980 84182
rect 92532 84166 92980 84176
rect 93768 84176 93820 84182
rect 92480 84118 92532 84124
rect 93768 84118 93820 84124
rect 91006 71088 91062 71097
rect 91006 71023 91062 71032
rect 89628 11008 89680 11014
rect 89628 10950 89680 10956
rect 91020 3534 91048 71023
rect 93780 44878 93808 84118
rect 95056 61464 95108 61470
rect 95056 61406 95108 61412
rect 93768 44872 93820 44878
rect 93768 44814 93820 44820
rect 92386 30968 92442 30977
rect 92386 30903 92442 30912
rect 92400 3534 92428 30903
rect 92480 6248 92532 6254
rect 92480 6190 92532 6196
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89364 462 89576 490
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 92492 3466 92520 6190
rect 92756 3596 92808 3602
rect 92756 3538 92808 3544
rect 92480 3460 92532 3466
rect 92480 3402 92532 3408
rect 92768 480 92796 3538
rect 95068 3058 95096 61406
rect 93952 3052 94004 3058
rect 93952 2994 94004 3000
rect 95056 3052 95108 3058
rect 95056 2994 95108 3000
rect 93964 480 93992 2994
rect 95160 480 95188 94279
rect 95252 91050 95280 122726
rect 95896 93566 95924 216679
rect 95988 111897 96016 227734
rect 96632 207670 96660 240110
rect 96724 220289 96752 241590
rect 97000 240174 97028 241590
rect 96988 240168 97040 240174
rect 97828 240145 97856 241590
rect 96988 240110 97040 240116
rect 97814 240136 97870 240145
rect 97814 240071 97870 240080
rect 97828 233918 97856 240071
rect 98104 238754 98132 259519
rect 98552 242956 98604 242962
rect 98552 242898 98604 242904
rect 98564 242298 98592 242898
rect 98440 242270 98592 242298
rect 98012 238726 98132 238754
rect 97906 234696 97962 234705
rect 97906 234631 97962 234640
rect 97816 233912 97868 233918
rect 97816 233854 97868 233860
rect 97446 230344 97502 230353
rect 97446 230279 97502 230288
rect 96710 220280 96766 220289
rect 96710 220215 96766 220224
rect 96620 207664 96672 207670
rect 96620 207606 96672 207612
rect 97354 204912 97410 204921
rect 97354 204847 97410 204856
rect 96068 134836 96120 134842
rect 96068 134778 96120 134784
rect 96080 122330 96108 134778
rect 96712 133884 96764 133890
rect 96712 133826 96764 133832
rect 96724 133113 96752 133826
rect 96710 133104 96766 133113
rect 96710 133039 96766 133048
rect 96620 132456 96672 132462
rect 96620 132398 96672 132404
rect 96632 132297 96660 132398
rect 96618 132288 96674 132297
rect 96618 132223 96674 132232
rect 97368 131481 97396 204847
rect 97460 133929 97488 230279
rect 97446 133920 97502 133929
rect 97446 133855 97502 133864
rect 97354 131472 97410 131481
rect 97354 131407 97410 131416
rect 97262 130928 97318 130937
rect 97262 130863 97318 130872
rect 96712 129736 96764 129742
rect 96712 129678 96764 129684
rect 96724 129305 96752 129678
rect 97276 129674 97304 130863
rect 97264 129668 97316 129674
rect 97264 129610 97316 129616
rect 96710 129296 96766 129305
rect 96710 129231 96766 129240
rect 97172 128240 97224 128246
rect 97172 128182 97224 128188
rect 97184 127673 97212 128182
rect 97170 127664 97226 127673
rect 97170 127599 97226 127608
rect 96802 125488 96858 125497
rect 96802 125423 96858 125432
rect 96816 124914 96844 125423
rect 96804 124908 96856 124914
rect 96804 124850 96856 124856
rect 96620 124024 96672 124030
rect 96618 123992 96620 124001
rect 96672 123992 96674 124001
rect 96618 123927 96674 123936
rect 96068 122324 96120 122330
rect 96068 122266 96120 122272
rect 96620 117088 96672 117094
rect 96618 117056 96620 117065
rect 96672 117056 96674 117065
rect 96618 116991 96674 117000
rect 96618 114064 96674 114073
rect 96618 113999 96674 114008
rect 96632 113898 96660 113999
rect 96620 113892 96672 113898
rect 96620 113834 96672 113840
rect 95974 111888 96030 111897
rect 95974 111823 96030 111832
rect 95974 101416 96030 101425
rect 95974 101351 96030 101360
rect 95884 93560 95936 93566
rect 95884 93502 95936 93508
rect 95240 91044 95292 91050
rect 95240 90986 95292 90992
rect 95988 88097 96016 101351
rect 96160 91044 96212 91050
rect 96160 90986 96212 90992
rect 95974 88088 96030 88097
rect 95974 88023 96030 88032
rect 96172 80714 96200 90986
rect 96160 80708 96212 80714
rect 96160 80650 96212 80656
rect 96528 71052 96580 71058
rect 96528 70994 96580 71000
rect 96540 6914 96568 70994
rect 96632 10334 96660 113834
rect 96816 103514 96844 124850
rect 97172 104848 97224 104854
rect 97172 104790 97224 104796
rect 97184 104281 97212 104790
rect 97170 104272 97226 104281
rect 97170 104207 97226 104216
rect 96724 103486 96844 103514
rect 97172 103488 97224 103494
rect 96724 86970 96752 103486
rect 97172 103430 97224 103436
rect 97184 102921 97212 103430
rect 97170 102912 97226 102921
rect 97170 102847 97226 102856
rect 96712 86964 96764 86970
rect 96712 86906 96764 86912
rect 97276 61402 97304 129610
rect 97540 128308 97592 128314
rect 97540 128250 97592 128256
rect 97552 127129 97580 128250
rect 97538 127120 97594 127129
rect 97538 127055 97594 127064
rect 97816 126948 97868 126954
rect 97816 126890 97868 126896
rect 97828 126313 97856 126890
rect 97814 126304 97870 126313
rect 97814 126239 97870 126248
rect 97448 125588 97500 125594
rect 97448 125530 97500 125536
rect 97460 124681 97488 125530
rect 97446 124672 97502 124681
rect 97446 124607 97502 124616
rect 97816 124160 97868 124166
rect 97816 124102 97868 124108
rect 97828 123321 97856 124102
rect 97814 123312 97870 123321
rect 97814 123247 97870 123256
rect 97816 122800 97868 122806
rect 97816 122742 97868 122748
rect 97828 122505 97856 122742
rect 97814 122496 97870 122505
rect 97814 122431 97870 122440
rect 97816 121440 97868 121446
rect 97816 121382 97868 121388
rect 97828 120873 97856 121382
rect 97814 120864 97870 120873
rect 97814 120799 97870 120808
rect 97814 120320 97870 120329
rect 97814 120255 97870 120264
rect 97828 120222 97856 120255
rect 97816 120216 97868 120222
rect 97816 120158 97868 120164
rect 97816 118652 97868 118658
rect 97816 118594 97868 118600
rect 97828 117881 97856 118594
rect 97814 117872 97870 117881
rect 97814 117807 97870 117816
rect 97816 117292 97868 117298
rect 97816 117234 97868 117240
rect 97828 116521 97856 117234
rect 97814 116512 97870 116521
rect 97814 116447 97870 116456
rect 97724 115932 97776 115938
rect 97724 115874 97776 115880
rect 97736 114889 97764 115874
rect 97816 115864 97868 115870
rect 97816 115806 97868 115812
rect 97828 115705 97856 115806
rect 97814 115696 97870 115705
rect 97814 115631 97870 115640
rect 97722 114880 97778 114889
rect 97722 114815 97778 114824
rect 97816 113144 97868 113150
rect 97816 113086 97868 113092
rect 97828 112713 97856 113086
rect 97814 112704 97870 112713
rect 97814 112639 97870 112648
rect 97920 111874 97948 234631
rect 98012 232665 98040 238726
rect 98656 233889 98684 261015
rect 98642 233880 98698 233889
rect 98642 233815 98698 233824
rect 99102 233880 99158 233889
rect 99102 233815 99158 233824
rect 97998 232656 98054 232665
rect 97998 232591 98054 232600
rect 98644 220856 98696 220862
rect 98644 220798 98696 220804
rect 98000 122324 98052 122330
rect 98000 122266 98052 122272
rect 97736 111846 97948 111874
rect 97736 109562 97764 111846
rect 97908 111784 97960 111790
rect 97908 111726 97960 111732
rect 97920 111081 97948 111726
rect 97906 111072 97962 111081
rect 97906 111007 97962 111016
rect 97816 110424 97868 110430
rect 97816 110366 97868 110372
rect 97828 109721 97856 110366
rect 97908 110356 97960 110362
rect 97908 110298 97960 110304
rect 97920 110265 97948 110298
rect 97906 110256 97962 110265
rect 97906 110191 97962 110200
rect 97814 109712 97870 109721
rect 97814 109647 97870 109656
rect 97736 109534 97856 109562
rect 97724 108928 97776 108934
rect 97724 108870 97776 108876
rect 97736 108089 97764 108870
rect 97722 108080 97778 108089
rect 97722 108015 97778 108024
rect 97540 107364 97592 107370
rect 97540 107306 97592 107312
rect 97552 106729 97580 107306
rect 97538 106720 97594 106729
rect 97538 106655 97594 106664
rect 97632 106276 97684 106282
rect 97632 106218 97684 106224
rect 97644 105097 97672 106218
rect 97828 105890 97856 109534
rect 97908 108996 97960 109002
rect 97908 108938 97960 108944
rect 97920 108905 97948 108938
rect 97906 108896 97962 108905
rect 97906 108831 97962 108840
rect 97906 105904 97962 105913
rect 97828 105862 97906 105890
rect 97906 105839 97962 105848
rect 97920 105602 97948 105839
rect 97908 105596 97960 105602
rect 97908 105538 97960 105544
rect 97630 105088 97686 105097
rect 97630 105023 97686 105032
rect 97724 102808 97776 102814
rect 97724 102750 97776 102756
rect 97354 100056 97410 100065
rect 97354 99991 97410 100000
rect 97368 92857 97396 99991
rect 97736 99657 97764 102750
rect 97908 102128 97960 102134
rect 97906 102096 97908 102105
rect 97960 102096 97962 102105
rect 97816 102060 97868 102066
rect 97906 102031 97962 102040
rect 97816 102002 97868 102008
rect 97828 101289 97856 102002
rect 97814 101280 97870 101289
rect 97814 101215 97870 101224
rect 97908 100700 97960 100706
rect 97908 100642 97960 100648
rect 97920 100473 97948 100642
rect 97906 100464 97962 100473
rect 97906 100399 97962 100408
rect 97722 99648 97778 99657
rect 97722 99583 97778 99592
rect 97540 99340 97592 99346
rect 97540 99282 97592 99288
rect 97552 98297 97580 99282
rect 97538 98288 97594 98297
rect 97538 98223 97594 98232
rect 97908 97980 97960 97986
rect 97908 97922 97960 97928
rect 97540 97912 97592 97918
rect 97540 97854 97592 97860
rect 97552 96665 97580 97854
rect 97920 97481 97948 97922
rect 97906 97472 97962 97481
rect 97906 97407 97962 97416
rect 97538 96656 97594 96665
rect 97538 96591 97594 96600
rect 97908 96008 97960 96014
rect 97908 95950 97960 95956
rect 97920 95305 97948 95950
rect 97906 95296 97962 95305
rect 97906 95231 97962 95240
rect 97908 95192 97960 95198
rect 97908 95134 97960 95140
rect 97920 94489 97948 95134
rect 97906 94480 97962 94489
rect 97906 94415 97962 94424
rect 97908 93832 97960 93838
rect 97908 93774 97960 93780
rect 97920 93673 97948 93774
rect 97906 93664 97962 93673
rect 97906 93599 97962 93608
rect 97354 92848 97410 92857
rect 97354 92783 97410 92792
rect 98012 85542 98040 122266
rect 98656 117094 98684 220798
rect 99116 214713 99144 233815
rect 99102 214704 99158 214713
rect 99102 214639 99158 214648
rect 99208 206310 99236 272031
rect 99288 242956 99340 242962
rect 99288 242898 99340 242904
rect 99196 206304 99248 206310
rect 99196 206246 99248 206252
rect 99208 205698 99236 206246
rect 98736 205692 98788 205698
rect 98736 205634 98788 205640
rect 99196 205692 99248 205698
rect 99196 205634 99248 205640
rect 98748 124030 98776 205634
rect 98736 124024 98788 124030
rect 98736 123966 98788 123972
rect 98644 117088 98696 117094
rect 98644 117030 98696 117036
rect 98642 115152 98698 115161
rect 98642 115087 98698 115096
rect 98656 90953 98684 115087
rect 98734 111072 98790 111081
rect 98734 111007 98790 111016
rect 98748 92410 98776 111007
rect 99300 96014 99328 242898
rect 99392 204921 99420 280191
rect 99484 279478 99512 283562
rect 99472 279472 99524 279478
rect 99472 279414 99524 279420
rect 100036 276690 100064 285631
rect 100024 276684 100076 276690
rect 100024 276626 100076 276632
rect 100128 265674 100156 301446
rect 100574 287464 100630 287473
rect 100574 287399 100630 287408
rect 100588 283529 100616 287399
rect 100574 283520 100630 283529
rect 100574 283455 100630 283464
rect 100680 282441 100708 306342
rect 100666 282432 100722 282441
rect 100666 282367 100722 282376
rect 100758 281072 100814 281081
rect 100758 281007 100814 281016
rect 100772 278769 100800 281007
rect 100758 278760 100814 278769
rect 100758 278695 100814 278704
rect 100758 275360 100814 275369
rect 100758 275295 100760 275304
rect 100812 275295 100814 275304
rect 100760 275266 100812 275272
rect 100850 274544 100906 274553
rect 100850 274479 100906 274488
rect 100760 274032 100812 274038
rect 100760 273974 100812 273980
rect 100772 273737 100800 273974
rect 100864 273970 100892 274479
rect 100852 273964 100904 273970
rect 100852 273906 100904 273912
rect 100758 273728 100814 273737
rect 100758 273663 100814 273672
rect 101416 272105 101444 384338
rect 101956 374672 102008 374678
rect 101956 374614 102008 374620
rect 101968 331294 101996 374614
rect 101496 331288 101548 331294
rect 101496 331230 101548 331236
rect 101956 331288 102008 331294
rect 101956 331230 102008 331236
rect 101508 280265 101536 331230
rect 101588 288516 101640 288522
rect 101588 288458 101640 288464
rect 101494 280256 101550 280265
rect 101494 280191 101550 280200
rect 101600 279449 101628 288458
rect 101586 279440 101642 279449
rect 101586 279375 101642 279384
rect 101954 278624 102010 278633
rect 101954 278559 102010 278568
rect 101968 275913 101996 278559
rect 102060 278050 102088 387087
rect 102152 327049 102180 390102
rect 102244 335481 102272 390374
rect 103518 389192 103574 389201
rect 103518 389127 103574 389136
rect 102322 388512 102378 388521
rect 102322 388447 102378 388456
rect 102336 378282 102364 388447
rect 103532 378894 103560 389127
rect 103716 388482 103744 390374
rect 103808 390374 104144 390402
rect 104880 390374 105216 390402
rect 103808 389201 103836 390374
rect 104808 389836 104860 389842
rect 104808 389778 104860 389784
rect 103794 389192 103850 389201
rect 103794 389127 103850 389136
rect 103704 388476 103756 388482
rect 103704 388418 103756 388424
rect 103520 378888 103572 378894
rect 103520 378830 103572 378836
rect 102324 378276 102376 378282
rect 102324 378218 102376 378224
rect 104256 376100 104308 376106
rect 104256 376042 104308 376048
rect 104164 354000 104216 354006
rect 104164 353942 104216 353948
rect 102230 335472 102286 335481
rect 102230 335407 102286 335416
rect 102138 327040 102194 327049
rect 102138 326975 102194 326984
rect 102782 323640 102838 323649
rect 102782 323575 102838 323584
rect 102232 287156 102284 287162
rect 102232 287098 102284 287104
rect 102048 278044 102100 278050
rect 102048 277986 102100 277992
rect 102060 277817 102088 277986
rect 102046 277808 102102 277817
rect 102046 277743 102102 277752
rect 102140 276344 102192 276350
rect 102140 276286 102192 276292
rect 102046 276176 102102 276185
rect 102152 276162 102180 276286
rect 102102 276134 102180 276162
rect 102046 276111 102102 276120
rect 101954 275904 102010 275913
rect 101954 275839 102010 275848
rect 101402 272096 101458 272105
rect 101402 272031 101458 272040
rect 101678 271280 101734 271289
rect 101678 271215 101734 271224
rect 101692 271182 101720 271215
rect 101680 271176 101732 271182
rect 101680 271118 101732 271124
rect 100760 269952 100812 269958
rect 100760 269894 100812 269900
rect 100772 269657 100800 269894
rect 100758 269648 100814 269657
rect 100758 269583 100814 269592
rect 100850 268832 100906 268841
rect 100850 268767 100906 268776
rect 100760 268456 100812 268462
rect 100760 268398 100812 268404
rect 100772 268025 100800 268398
rect 100864 268394 100892 268767
rect 100852 268388 100904 268394
rect 100852 268330 100904 268336
rect 100758 268016 100814 268025
rect 100758 267951 100814 267960
rect 101402 267200 101458 267209
rect 101402 267135 101458 267144
rect 100116 265668 100168 265674
rect 100116 265610 100168 265616
rect 100022 265568 100078 265577
rect 100022 265503 100078 265512
rect 99470 252512 99526 252521
rect 99470 252447 99526 252456
rect 99484 234705 99512 252447
rect 99470 234696 99526 234705
rect 99470 234631 99526 234640
rect 100036 234025 100064 265503
rect 100852 264988 100904 264994
rect 100852 264930 100904 264936
rect 100758 264752 100814 264761
rect 100758 264687 100814 264696
rect 100772 264246 100800 264687
rect 100760 264240 100812 264246
rect 100760 264182 100812 264188
rect 100758 263936 100814 263945
rect 100758 263871 100814 263880
rect 100772 263634 100800 263871
rect 100760 263628 100812 263634
rect 100760 263570 100812 263576
rect 100758 263120 100814 263129
rect 100758 263055 100814 263064
rect 100772 262954 100800 263055
rect 100760 262948 100812 262954
rect 100760 262890 100812 262896
rect 100864 262313 100892 264930
rect 100850 262304 100906 262313
rect 100850 262239 100906 262248
rect 100760 261520 100812 261526
rect 100758 261488 100760 261497
rect 100812 261488 100814 261497
rect 100758 261423 100814 261432
rect 100850 260672 100906 260681
rect 100850 260607 100906 260616
rect 100864 259486 100892 260607
rect 100852 259480 100904 259486
rect 100852 259422 100904 259428
rect 100850 259040 100906 259049
rect 100850 258975 100906 258984
rect 100760 258800 100812 258806
rect 100760 258742 100812 258748
rect 100772 258233 100800 258742
rect 100864 258738 100892 258975
rect 100852 258732 100904 258738
rect 100852 258674 100904 258680
rect 100758 258224 100814 258233
rect 100864 258194 100892 258674
rect 100758 258159 100814 258168
rect 100852 258188 100904 258194
rect 100852 258130 100904 258136
rect 100760 258120 100812 258126
rect 100760 258062 100812 258068
rect 100392 252544 100444 252550
rect 100390 252512 100392 252521
rect 100444 252512 100446 252521
rect 100390 252447 100446 252456
rect 100022 234016 100078 234025
rect 100022 233951 100078 233960
rect 100668 233300 100720 233306
rect 100668 233242 100720 233248
rect 100574 229800 100630 229809
rect 100574 229735 100630 229744
rect 100588 218657 100616 229735
rect 100574 218648 100630 218657
rect 100574 218583 100630 218592
rect 100680 213246 100708 233242
rect 100772 227798 100800 258062
rect 100852 258052 100904 258058
rect 100852 257994 100904 258000
rect 100864 257417 100892 257994
rect 100850 257408 100906 257417
rect 100850 257343 100906 257352
rect 101034 257272 101090 257281
rect 101034 257207 101090 257216
rect 100942 256592 100998 256601
rect 100942 256527 100998 256536
rect 100852 256012 100904 256018
rect 100852 255954 100904 255960
rect 100864 255785 100892 255954
rect 100850 255776 100906 255785
rect 100850 255711 100906 255720
rect 100956 255338 100984 256527
rect 100944 255332 100996 255338
rect 100944 255274 100996 255280
rect 101048 254153 101076 257207
rect 101034 254144 101090 254153
rect 101034 254079 101090 254088
rect 100850 250880 100906 250889
rect 100850 250815 100906 250824
rect 100864 250510 100892 250815
rect 100852 250504 100904 250510
rect 100852 250446 100904 250452
rect 100850 250064 100906 250073
rect 100850 249999 100906 250008
rect 100864 249830 100892 249999
rect 100852 249824 100904 249830
rect 100852 249766 100904 249772
rect 100944 249756 100996 249762
rect 100944 249698 100996 249704
rect 100850 249248 100906 249257
rect 100850 249183 100906 249192
rect 100864 249082 100892 249183
rect 100852 249076 100904 249082
rect 100852 249018 100904 249024
rect 100956 248441 100984 249698
rect 100942 248432 100998 248441
rect 100852 248396 100904 248402
rect 100942 248367 100998 248376
rect 100852 248338 100904 248344
rect 100864 247625 100892 248338
rect 100850 247616 100906 247625
rect 100850 247551 100906 247560
rect 100852 246968 100904 246974
rect 100852 246910 100904 246916
rect 100864 246809 100892 246910
rect 100850 246800 100906 246809
rect 100850 246735 100906 246744
rect 100852 246356 100904 246362
rect 100852 246298 100904 246304
rect 100864 245993 100892 246298
rect 100850 245984 100906 245993
rect 100850 245919 100906 245928
rect 100944 245608 100996 245614
rect 100944 245550 100996 245556
rect 100850 245168 100906 245177
rect 100850 245103 100906 245112
rect 100864 244322 100892 245103
rect 100956 244361 100984 245550
rect 100942 244352 100998 244361
rect 100852 244316 100904 244322
rect 100942 244287 100998 244296
rect 100852 244258 100904 244264
rect 100852 242752 100904 242758
rect 100850 242720 100852 242729
rect 100904 242720 100906 242729
rect 100850 242655 100906 242664
rect 100850 241904 100906 241913
rect 100850 241839 100906 241848
rect 100864 233306 100892 241839
rect 101416 235521 101444 267135
rect 101494 254960 101550 254969
rect 101494 254895 101550 254904
rect 101402 235512 101458 235521
rect 101402 235447 101458 235456
rect 100852 233300 100904 233306
rect 100852 233242 100904 233248
rect 100760 227792 100812 227798
rect 100760 227734 100812 227740
rect 101508 225622 101536 254895
rect 102152 225690 102180 276134
rect 102244 237386 102272 287098
rect 102796 276350 102824 323575
rect 103426 318200 103482 318209
rect 103426 318135 103482 318144
rect 102784 276344 102836 276350
rect 102784 276286 102836 276292
rect 102322 273320 102378 273329
rect 102322 273255 102378 273264
rect 102232 237380 102284 237386
rect 102232 237322 102284 237328
rect 102244 236706 102272 237322
rect 102232 236700 102284 236706
rect 102232 236642 102284 236648
rect 102336 235550 102364 273255
rect 103440 271182 103468 318135
rect 103518 289096 103574 289105
rect 103518 289031 103574 289040
rect 103428 271176 103480 271182
rect 103428 271118 103480 271124
rect 102784 254584 102836 254590
rect 102784 254526 102836 254532
rect 102796 237153 102824 254526
rect 103428 243636 103480 243642
rect 103428 243578 103480 243584
rect 103440 242962 103468 243578
rect 103428 242956 103480 242962
rect 103428 242898 103480 242904
rect 103440 240106 103468 242898
rect 103428 240100 103480 240106
rect 103428 240042 103480 240048
rect 103532 238746 103560 289031
rect 104176 273222 104204 353942
rect 104268 304201 104296 376042
rect 104254 304192 104310 304201
rect 104254 304127 104310 304136
rect 104438 304192 104494 304201
rect 104438 304127 104494 304136
rect 104164 273216 104216 273222
rect 104164 273158 104216 273164
rect 104346 271144 104402 271153
rect 104346 271079 104402 271088
rect 103978 270464 104034 270473
rect 103978 270399 104034 270408
rect 103992 269142 104020 270399
rect 103980 269136 104032 269142
rect 103980 269078 104032 269084
rect 104164 262880 104216 262886
rect 104164 262822 104216 262828
rect 104176 240145 104204 262822
rect 104360 262177 104388 271079
rect 104452 269958 104480 304127
rect 104440 269952 104492 269958
rect 104440 269894 104492 269900
rect 104452 267034 104480 269894
rect 104440 267028 104492 267034
rect 104440 266970 104492 266976
rect 104346 262168 104402 262177
rect 104346 262103 104402 262112
rect 104820 261526 104848 389778
rect 105188 386374 105216 390374
rect 105322 390374 106044 390402
rect 105266 390351 105322 390360
rect 105176 386368 105228 386374
rect 105176 386310 105228 386316
rect 104900 384328 104952 384334
rect 104900 384270 104952 384276
rect 104912 383625 104940 384270
rect 106016 383654 106044 390374
rect 106338 390130 106366 390388
rect 106292 390102 106366 390130
rect 106016 383626 106228 383654
rect 104898 383616 104954 383625
rect 104898 383551 104954 383560
rect 104912 382401 104940 383551
rect 104898 382392 104954 382401
rect 104898 382327 104954 382336
rect 105544 376032 105596 376038
rect 105544 375974 105596 375980
rect 104992 293276 105044 293282
rect 104992 293218 105044 293224
rect 104900 269068 104952 269074
rect 104900 269010 104952 269016
rect 104912 268462 104940 269010
rect 104900 268456 104952 268462
rect 104900 268398 104952 268404
rect 104808 261520 104860 261526
rect 104808 261462 104860 261468
rect 104256 261112 104308 261118
rect 104256 261054 104308 261060
rect 104268 242758 104296 261054
rect 104348 256760 104400 256766
rect 104348 256702 104400 256708
rect 104360 246974 104388 256702
rect 104348 246968 104400 246974
rect 104348 246910 104400 246916
rect 104256 242752 104308 242758
rect 104256 242694 104308 242700
rect 104162 240136 104218 240145
rect 104162 240071 104218 240080
rect 103520 238740 103572 238746
rect 103520 238682 103572 238688
rect 102782 237144 102838 237153
rect 102782 237079 102838 237088
rect 102324 235544 102376 235550
rect 102324 235486 102376 235492
rect 102784 235272 102836 235278
rect 102784 235214 102836 235220
rect 102140 225684 102192 225690
rect 102140 225626 102192 225632
rect 101496 225616 101548 225622
rect 101496 225558 101548 225564
rect 100668 213240 100720 213246
rect 100668 213182 100720 213188
rect 99378 204912 99434 204921
rect 99378 204847 99434 204856
rect 102140 199436 102192 199442
rect 102140 199378 102192 199384
rect 100852 142180 100904 142186
rect 100852 142122 100904 142128
rect 99380 135244 99432 135250
rect 99380 135186 99432 135192
rect 99288 96008 99340 96014
rect 99288 95950 99340 95956
rect 98736 92404 98788 92410
rect 98736 92346 98788 92352
rect 98642 90944 98698 90953
rect 98642 90879 98698 90888
rect 98000 85536 98052 85542
rect 98000 85478 98052 85484
rect 99392 84114 99420 135186
rect 100758 134600 100814 134609
rect 100758 134535 100814 134544
rect 100024 116340 100076 116346
rect 100024 116282 100076 116288
rect 100036 89622 100064 116282
rect 100024 89616 100076 89622
rect 100024 89558 100076 89564
rect 99380 84108 99432 84114
rect 99380 84050 99432 84056
rect 100772 78674 100800 134535
rect 100864 128246 100892 142122
rect 100852 128240 100904 128246
rect 100852 128182 100904 128188
rect 101496 126268 101548 126274
rect 101496 126210 101548 126216
rect 101404 111036 101456 111042
rect 101404 110978 101456 110984
rect 100760 78668 100812 78674
rect 100760 78610 100812 78616
rect 101128 78668 101180 78674
rect 101128 78610 101180 78616
rect 101140 77994 101168 78610
rect 101128 77988 101180 77994
rect 101128 77930 101180 77936
rect 101416 71738 101444 110978
rect 101508 86902 101536 126210
rect 102152 112690 102180 199378
rect 102232 156732 102284 156738
rect 102232 156674 102284 156680
rect 102244 113174 102272 156674
rect 102796 140078 102824 235214
rect 103520 233300 103572 233306
rect 103520 233242 103572 233248
rect 103532 227662 103560 233242
rect 103520 227656 103572 227662
rect 103520 227598 103572 227604
rect 103426 225992 103482 226001
rect 103426 225927 103482 225936
rect 103440 204270 103468 225927
rect 102968 204264 103020 204270
rect 102968 204206 103020 204212
rect 103428 204264 103480 204270
rect 103428 204206 103480 204212
rect 102874 200016 102930 200025
rect 102874 199951 102930 199960
rect 102784 140072 102836 140078
rect 102784 140014 102836 140020
rect 102784 137352 102836 137358
rect 102784 137294 102836 137300
rect 102796 113830 102824 137294
rect 102888 128489 102916 199951
rect 102980 199510 103008 204206
rect 102968 199504 103020 199510
rect 102968 199446 103020 199452
rect 102874 128480 102930 128489
rect 102874 128415 102930 128424
rect 102784 113824 102836 113830
rect 102784 113766 102836 113772
rect 102244 113146 102456 113174
rect 102152 112662 102364 112690
rect 102140 112464 102192 112470
rect 102140 112406 102192 112412
rect 102152 107370 102180 112406
rect 102140 107364 102192 107370
rect 102140 107306 102192 107312
rect 102336 104786 102364 112662
rect 102324 104780 102376 104786
rect 102324 104722 102376 104728
rect 102046 104136 102102 104145
rect 102046 104071 102102 104080
rect 101496 86896 101548 86902
rect 101496 86838 101548 86844
rect 101404 71732 101456 71738
rect 101404 71674 101456 71680
rect 97264 61396 97316 61402
rect 97264 61338 97316 61344
rect 97908 17332 97960 17338
rect 97908 17274 97960 17280
rect 96620 10328 96672 10334
rect 96620 10270 96672 10276
rect 96264 6886 96568 6914
rect 96264 480 96292 6886
rect 97920 3534 97948 17274
rect 101034 7576 101090 7585
rect 101034 7511 101090 7520
rect 98642 3632 98698 3641
rect 98642 3567 98698 3576
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 97908 3528 97960 3534
rect 97908 3470 97960 3476
rect 97460 480 97488 3470
rect 98656 480 98684 3567
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 99852 480 99880 3470
rect 101048 480 101076 7511
rect 102060 3482 102088 104071
rect 102428 103514 102456 113146
rect 103428 106956 103480 106962
rect 103428 106898 103480 106904
rect 102244 103486 102456 103514
rect 102244 87961 102272 103486
rect 102230 87952 102286 87961
rect 102230 87887 102286 87896
rect 103440 6914 103468 106898
rect 103532 93158 103560 227598
rect 104176 217462 104204 240071
rect 104268 238066 104296 242694
rect 104256 238060 104308 238066
rect 104256 238002 104308 238008
rect 104806 228304 104862 228313
rect 104806 228239 104862 228248
rect 104164 217456 104216 217462
rect 104164 217398 104216 217404
rect 103612 209092 103664 209098
rect 103612 209034 103664 209040
rect 103520 93152 103572 93158
rect 103520 93094 103572 93100
rect 103624 85513 103652 209034
rect 104162 137320 104218 137329
rect 104162 137255 104218 137264
rect 104176 124817 104204 137255
rect 104162 124808 104218 124817
rect 104162 124743 104218 124752
rect 103610 85504 103666 85513
rect 103610 85439 103666 85448
rect 104820 6914 104848 228239
rect 104912 120222 104940 268398
rect 105004 238678 105032 293218
rect 105082 262168 105138 262177
rect 105082 262103 105138 262112
rect 104992 238672 105044 238678
rect 104992 238614 105044 238620
rect 104990 207632 105046 207641
rect 104990 207567 105046 207576
rect 104900 120216 104952 120222
rect 104900 120158 104952 120164
rect 104912 111042 104940 120158
rect 105004 116346 105032 207567
rect 105096 203590 105124 262103
rect 105556 243574 105584 375974
rect 106096 371272 106148 371278
rect 106096 371214 106148 371220
rect 106108 315314 106136 371214
rect 106200 322153 106228 383626
rect 106186 322144 106242 322153
rect 106186 322079 106242 322088
rect 106096 315308 106148 315314
rect 106096 315250 106148 315256
rect 105636 299056 105688 299062
rect 105636 298998 105688 299004
rect 105648 270473 105676 298998
rect 105634 270464 105690 270473
rect 105634 270399 105690 270408
rect 106094 256320 106150 256329
rect 106094 256255 106150 256264
rect 106108 255338 106136 256255
rect 106096 255332 106148 255338
rect 106096 255274 106148 255280
rect 106292 243642 106320 390102
rect 106660 389162 106688 391002
rect 112732 390726 112760 471242
rect 113270 441008 113326 441017
rect 113270 440943 113326 440952
rect 113180 433832 113232 433838
rect 113180 433774 113232 433780
rect 112812 433696 112864 433702
rect 112812 433638 112864 433644
rect 112824 433294 112852 433638
rect 112812 433288 112864 433294
rect 112812 433230 112864 433236
rect 113192 429321 113220 433774
rect 113284 431225 113312 440943
rect 113270 431216 113326 431225
rect 113270 431151 113326 431160
rect 113178 429312 113234 429321
rect 113178 429247 113234 429256
rect 113178 420064 113234 420073
rect 113178 419999 113234 420008
rect 112168 390720 112220 390726
rect 107750 390688 107806 390697
rect 107750 390623 107806 390632
rect 108762 390688 108818 390697
rect 108762 390623 108818 390632
rect 111706 390688 111762 390697
rect 111872 390668 112168 390674
rect 111872 390662 112220 390668
rect 112720 390720 112772 390726
rect 112720 390662 112772 390668
rect 111872 390660 112208 390662
rect 111706 390623 111762 390632
rect 111858 390646 112208 390660
rect 107764 390538 107792 390623
rect 107640 390510 107792 390538
rect 106738 390416 106794 390425
rect 106794 390374 107516 390402
rect 106738 390351 106794 390360
rect 106648 389156 106700 389162
rect 106648 389098 106700 389104
rect 106924 383036 106976 383042
rect 106924 382978 106976 382984
rect 106372 282940 106424 282946
rect 106372 282882 106424 282888
rect 106280 243636 106332 243642
rect 106280 243578 106332 243584
rect 105544 243568 105596 243574
rect 105544 243510 105596 243516
rect 105542 236600 105598 236609
rect 105542 236535 105598 236544
rect 105084 203584 105136 203590
rect 105084 203526 105136 203532
rect 104992 116340 105044 116346
rect 104992 116282 105044 116288
rect 104900 111036 104952 111042
rect 104900 110978 104952 110984
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 102060 3454 102272 3482
rect 102244 480 102272 3454
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 105556 3505 105584 236535
rect 106280 204944 106332 204950
rect 106280 204886 106332 204892
rect 105636 202088 105688 202094
rect 105636 202030 105688 202036
rect 105648 85377 105676 202030
rect 106292 92478 106320 204886
rect 106384 141506 106412 282882
rect 106830 269240 106886 269249
rect 106830 269175 106886 269184
rect 106844 269142 106872 269175
rect 106832 269136 106884 269142
rect 106832 269078 106884 269084
rect 106936 253978 106964 382978
rect 107488 381546 107516 390374
rect 107764 389065 107792 390510
rect 108376 390374 108712 390402
rect 107750 389056 107806 389065
rect 107750 388991 107806 389000
rect 108684 385014 108712 390374
rect 108672 385008 108724 385014
rect 108672 384950 108724 384956
rect 108776 383654 108804 390623
rect 109098 390130 109126 390388
rect 109848 390374 110184 390402
rect 110400 390374 110736 390402
rect 109052 390102 109126 390130
rect 108946 389056 109002 389065
rect 108946 388991 109002 389000
rect 108776 383626 108896 383654
rect 107476 381540 107528 381546
rect 107476 381482 107528 381488
rect 108868 326398 108896 383626
rect 108856 326392 108908 326398
rect 108856 326334 108908 326340
rect 108856 321632 108908 321638
rect 108856 321574 108908 321580
rect 107568 285728 107620 285734
rect 107568 285670 107620 285676
rect 107580 284209 107608 285670
rect 107014 284200 107070 284209
rect 107014 284135 107070 284144
rect 107566 284200 107622 284209
rect 107566 284135 107622 284144
rect 106924 253972 106976 253978
rect 106924 253914 106976 253920
rect 106646 249112 106702 249121
rect 106646 249047 106648 249056
rect 106700 249047 106702 249056
rect 106648 249018 106700 249024
rect 106464 239420 106516 239426
rect 106464 239362 106516 239368
rect 106372 141500 106424 141506
rect 106372 141442 106424 141448
rect 106476 126274 106504 239362
rect 106936 233238 106964 253914
rect 107028 235278 107056 284135
rect 107844 279472 107896 279478
rect 107844 279414 107896 279420
rect 107660 265668 107712 265674
rect 107660 265610 107712 265616
rect 107672 240009 107700 265610
rect 107752 252612 107804 252618
rect 107752 252554 107804 252560
rect 107764 250510 107792 252554
rect 107752 250504 107804 250510
rect 107752 250446 107804 250452
rect 107658 240000 107714 240009
rect 107658 239935 107714 239944
rect 107658 237960 107714 237969
rect 107658 237895 107714 237904
rect 107016 235272 107068 235278
rect 107016 235214 107068 235220
rect 106924 233232 106976 233238
rect 106924 233174 106976 233180
rect 107568 218748 107620 218754
rect 107568 218690 107620 218696
rect 106924 140820 106976 140826
rect 106924 140762 106976 140768
rect 106464 126268 106516 126274
rect 106464 126210 106516 126216
rect 106936 97918 106964 140762
rect 106924 97912 106976 97918
rect 106924 97854 106976 97860
rect 106280 92472 106332 92478
rect 106280 92414 106332 92420
rect 105634 85368 105690 85377
rect 105634 85303 105690 85312
rect 105726 8936 105782 8945
rect 105726 8871 105782 8880
rect 105542 3496 105598 3505
rect 105542 3431 105598 3440
rect 105740 480 105768 8871
rect 107580 3534 107608 218690
rect 107672 82822 107700 237895
rect 107764 104854 107792 250446
rect 107856 196654 107884 279414
rect 108304 279268 108356 279274
rect 108304 279210 108356 279216
rect 108316 261118 108344 279210
rect 108868 267734 108896 321574
rect 108960 280158 108988 388991
rect 108948 280152 109000 280158
rect 108948 280094 109000 280100
rect 108960 279274 108988 280094
rect 108948 279268 109000 279274
rect 108948 279210 109000 279216
rect 108868 267706 108988 267734
rect 108304 261112 108356 261118
rect 108304 261054 108356 261060
rect 108960 248402 108988 267706
rect 109052 252482 109080 390102
rect 110156 389162 110184 390374
rect 110144 389156 110196 389162
rect 110144 389098 110196 389104
rect 110708 387841 110736 390374
rect 110800 390374 111136 390402
rect 110694 387832 110750 387841
rect 110694 387767 110750 387776
rect 110800 373994 110828 390374
rect 110432 373966 110828 373994
rect 109682 325000 109738 325009
rect 109682 324935 109738 324944
rect 109316 308440 109368 308446
rect 109316 308382 109368 308388
rect 109328 307834 109356 308382
rect 109316 307828 109368 307834
rect 109316 307770 109368 307776
rect 109132 288448 109184 288454
rect 109132 288390 109184 288396
rect 109040 252476 109092 252482
rect 109040 252418 109092 252424
rect 108948 248396 109000 248402
rect 108948 248338 109000 248344
rect 108960 247722 108988 248338
rect 108948 247716 109000 247722
rect 108948 247658 109000 247664
rect 109040 246356 109092 246362
rect 109040 246298 109092 246304
rect 109052 246265 109080 246298
rect 109038 246256 109094 246265
rect 109038 246191 109094 246200
rect 108304 227044 108356 227050
rect 108304 226986 108356 226992
rect 107844 196648 107896 196654
rect 107844 196590 107896 196596
rect 107752 104848 107804 104854
rect 107752 104790 107804 104796
rect 107660 82816 107712 82822
rect 107660 82758 107712 82764
rect 108316 3670 108344 226986
rect 109038 207768 109094 207777
rect 109038 207703 109094 207712
rect 109052 91089 109080 207703
rect 109144 135930 109172 288390
rect 109224 261520 109276 261526
rect 109224 261462 109276 261468
rect 109132 135924 109184 135930
rect 109132 135866 109184 135872
rect 109236 113898 109264 261462
rect 109328 233170 109356 307770
rect 109696 277394 109724 324935
rect 109604 277366 109724 277394
rect 109604 269074 109632 277366
rect 109682 273184 109738 273193
rect 109682 273119 109738 273128
rect 109696 271930 109724 273119
rect 109684 271924 109736 271930
rect 109684 271866 109736 271872
rect 109592 269068 109644 269074
rect 109592 269010 109644 269016
rect 110432 257378 110460 373966
rect 111720 330449 111748 390623
rect 111858 390130 111886 390646
rect 112272 390374 112608 390402
rect 111858 390102 111932 390130
rect 111800 387048 111852 387054
rect 111800 386990 111852 386996
rect 111706 330440 111762 330449
rect 111706 330375 111762 330384
rect 111064 305652 111116 305658
rect 111064 305594 111116 305600
rect 110604 295384 110656 295390
rect 110604 295326 110656 295332
rect 110512 287700 110564 287706
rect 110512 287642 110564 287648
rect 110524 287094 110552 287642
rect 110512 287088 110564 287094
rect 110512 287030 110564 287036
rect 110420 257372 110472 257378
rect 110420 257314 110472 257320
rect 110432 256766 110460 257314
rect 110420 256760 110472 256766
rect 110420 256702 110472 256708
rect 109684 252476 109736 252482
rect 109684 252418 109736 252424
rect 109696 251258 109724 252418
rect 109684 251252 109736 251258
rect 109684 251194 109736 251200
rect 109696 245614 109724 251194
rect 109684 245608 109736 245614
rect 109684 245550 109736 245556
rect 109316 233164 109368 233170
rect 109316 233106 109368 233112
rect 110420 217456 110472 217462
rect 110420 217398 110472 217404
rect 109314 206272 109370 206281
rect 109314 206207 109370 206216
rect 109224 113892 109276 113898
rect 109224 113834 109276 113840
rect 109328 101425 109356 206207
rect 109314 101416 109370 101425
rect 109314 101351 109370 101360
rect 110432 95198 110460 217398
rect 110524 140758 110552 287030
rect 110616 216578 110644 295326
rect 111076 252618 111104 305594
rect 111064 252612 111116 252618
rect 111064 252554 111116 252560
rect 111812 249762 111840 386990
rect 111904 321638 111932 390102
rect 112272 387054 112300 390374
rect 112260 387048 112312 387054
rect 112260 386990 112312 386996
rect 113192 384402 113220 419999
rect 113376 416809 113404 579634
rect 114652 569288 114704 569294
rect 114652 569230 114704 569236
rect 114560 558952 114612 558958
rect 114560 558894 114612 558900
rect 114100 434784 114152 434790
rect 114100 434726 114152 434732
rect 113454 430128 113510 430137
rect 113454 430063 113510 430072
rect 113362 416800 113418 416809
rect 113362 416735 113418 416744
rect 113180 384396 113232 384402
rect 113180 384338 113232 384344
rect 113468 374678 113496 430063
rect 113822 429312 113878 429321
rect 113822 429247 113878 429256
rect 113456 374672 113508 374678
rect 113456 374614 113508 374620
rect 112444 356720 112496 356726
rect 112444 356662 112496 356668
rect 111892 321632 111944 321638
rect 111892 321574 111944 321580
rect 111892 318164 111944 318170
rect 111892 318106 111944 318112
rect 111904 317490 111932 318106
rect 111892 317484 111944 317490
rect 111892 317426 111944 317432
rect 111800 249756 111852 249762
rect 111800 249698 111852 249704
rect 111616 248464 111668 248470
rect 111616 248406 111668 248412
rect 111064 241596 111116 241602
rect 111064 241538 111116 241544
rect 111076 235958 111104 241538
rect 111064 235952 111116 235958
rect 111064 235894 111116 235900
rect 110604 216572 110656 216578
rect 110604 216514 110656 216520
rect 110616 215966 110644 216514
rect 110604 215960 110656 215966
rect 110604 215902 110656 215908
rect 110512 140752 110564 140758
rect 110512 140694 110564 140700
rect 111628 138718 111656 248406
rect 111800 243568 111852 243574
rect 111800 243510 111852 243516
rect 111812 234598 111840 243510
rect 111904 237318 111932 317426
rect 112076 289876 112128 289882
rect 112076 289818 112128 289824
rect 111892 237312 111944 237318
rect 111892 237254 111944 237260
rect 111800 234592 111852 234598
rect 111800 234534 111852 234540
rect 111706 186960 111762 186969
rect 111706 186895 111762 186904
rect 111616 138712 111668 138718
rect 111616 138654 111668 138660
rect 110420 95192 110472 95198
rect 110420 95134 110472 95140
rect 109038 91080 109094 91089
rect 109038 91015 109094 91024
rect 108948 73840 109000 73846
rect 108948 73782 109000 73788
rect 108304 3664 108356 3670
rect 108304 3606 108356 3612
rect 108960 3534 108988 73782
rect 111720 6914 111748 186895
rect 111812 88330 111840 234534
rect 111984 225616 112036 225622
rect 111984 225558 112036 225564
rect 111890 214704 111946 214713
rect 111890 214639 111946 214648
rect 111904 97986 111932 214639
rect 111996 108934 112024 225558
rect 112088 222902 112116 289818
rect 112258 271960 112314 271969
rect 112258 271895 112260 271904
rect 112312 271895 112314 271904
rect 112260 271866 112312 271872
rect 112456 250510 112484 356662
rect 113836 349178 113864 429247
rect 114112 426494 114140 434726
rect 114100 426488 114152 426494
rect 114100 426430 114152 426436
rect 114112 424969 114140 426430
rect 114098 424960 114154 424969
rect 114098 424895 114154 424904
rect 114572 422294 114600 558894
rect 114664 424153 114692 569230
rect 115940 550656 115992 550662
rect 115940 550598 115992 550604
rect 115202 435296 115258 435305
rect 115202 435231 115258 435240
rect 114742 432304 114798 432313
rect 114742 432239 114798 432248
rect 114756 432002 114784 432239
rect 114744 431996 114796 432002
rect 114744 431938 114796 431944
rect 114742 431216 114798 431225
rect 114742 431151 114798 431160
rect 114756 430642 114784 431151
rect 114744 430636 114796 430642
rect 114744 430578 114796 430584
rect 114650 424144 114706 424153
rect 114650 424079 114706 424088
rect 115216 422294 115244 435231
rect 115386 428224 115442 428233
rect 115386 428159 115442 428168
rect 115400 427854 115428 428159
rect 115388 427848 115440 427854
rect 115388 427790 115440 427796
rect 115846 426048 115902 426057
rect 115846 425983 115902 425992
rect 115860 425134 115888 425983
rect 115848 425128 115900 425134
rect 115848 425070 115900 425076
rect 115848 424380 115900 424386
rect 115848 424322 115900 424328
rect 115860 424153 115888 424322
rect 115846 424144 115902 424153
rect 115846 424079 115902 424088
rect 115846 423056 115902 423065
rect 115846 422991 115902 423000
rect 115860 422958 115888 422991
rect 115848 422952 115900 422958
rect 115848 422894 115900 422900
rect 114572 422266 114968 422294
rect 114742 418976 114798 418985
rect 114742 418911 114798 418920
rect 114650 417888 114706 417897
rect 114650 417823 114706 417832
rect 114558 406464 114614 406473
rect 114558 406399 114614 406408
rect 114572 398138 114600 406399
rect 114560 398132 114612 398138
rect 114560 398074 114612 398080
rect 114468 378820 114520 378826
rect 114468 378762 114520 378768
rect 113824 349172 113876 349178
rect 113824 349114 113876 349120
rect 113836 288522 113864 349114
rect 114480 320686 114508 378762
rect 113916 320680 113968 320686
rect 113916 320622 113968 320628
rect 114468 320680 114520 320686
rect 114468 320622 114520 320628
rect 113824 288516 113876 288522
rect 113824 288458 113876 288464
rect 113364 280832 113416 280838
rect 113364 280774 113416 280780
rect 113272 268388 113324 268394
rect 113272 268330 113324 268336
rect 113180 260772 113232 260778
rect 113180 260714 113232 260720
rect 113192 256018 113220 260714
rect 113180 256012 113232 256018
rect 113180 255954 113232 255960
rect 112444 250504 112496 250510
rect 112444 250446 112496 250452
rect 112352 249756 112404 249762
rect 112352 249698 112404 249704
rect 112364 249150 112392 249698
rect 112352 249144 112404 249150
rect 112352 249086 112404 249092
rect 112168 240848 112220 240854
rect 112168 240790 112220 240796
rect 112076 222896 112128 222902
rect 112076 222838 112128 222844
rect 112180 202094 112208 240790
rect 112168 202088 112220 202094
rect 112168 202030 112220 202036
rect 113192 109002 113220 255954
rect 113284 121446 113312 268330
rect 113376 138786 113404 280774
rect 113836 276758 113864 288458
rect 113824 276752 113876 276758
rect 113824 276694 113876 276700
rect 113928 268394 113956 320622
rect 114480 320210 114508 320622
rect 114468 320204 114520 320210
rect 114468 320146 114520 320152
rect 114468 311160 114520 311166
rect 114468 311102 114520 311108
rect 114480 310554 114508 311102
rect 114468 310548 114520 310554
rect 114468 310490 114520 310496
rect 113916 268388 113968 268394
rect 113916 268330 113968 268336
rect 114480 233918 114508 310490
rect 114664 307873 114692 417823
rect 114756 318209 114784 418911
rect 114940 406473 114968 422266
rect 115124 422266 115244 422294
rect 115124 415562 115152 422266
rect 115848 422000 115900 422006
rect 115846 421968 115848 421977
rect 115900 421968 115902 421977
rect 115846 421903 115902 421912
rect 115848 416832 115900 416838
rect 115846 416800 115848 416809
rect 115900 416800 115902 416809
rect 115846 416735 115902 416744
rect 115204 415744 115256 415750
rect 115202 415712 115204 415721
rect 115256 415712 115258 415721
rect 115202 415647 115258 415656
rect 115124 415534 115244 415562
rect 115216 414050 115244 415534
rect 115848 414928 115900 414934
rect 115846 414896 115848 414905
rect 115900 414896 115902 414905
rect 115846 414831 115902 414840
rect 115204 414044 115256 414050
rect 115204 413986 115256 413992
rect 115216 412729 115244 413986
rect 115848 413976 115900 413982
rect 115848 413918 115900 413924
rect 115860 413817 115888 413918
rect 115846 413808 115902 413817
rect 115846 413743 115902 413752
rect 115202 412720 115258 412729
rect 115202 412655 115258 412664
rect 115848 412072 115900 412078
rect 115848 412014 115900 412020
rect 115860 411641 115888 412014
rect 115846 411632 115902 411641
rect 115846 411567 115902 411576
rect 115848 410576 115900 410582
rect 115846 410544 115848 410553
rect 115900 410544 115902 410553
rect 115846 410479 115902 410488
rect 115846 409728 115902 409737
rect 115846 409663 115902 409672
rect 115860 408542 115888 409663
rect 115848 408536 115900 408542
rect 115848 408478 115900 408484
rect 115846 407552 115902 407561
rect 115846 407487 115902 407496
rect 115860 407182 115888 407487
rect 115848 407176 115900 407182
rect 115848 407118 115900 407124
rect 114926 406464 114982 406473
rect 114926 406399 114982 406408
rect 115572 405680 115624 405686
rect 115572 405622 115624 405628
rect 115846 405648 115902 405657
rect 115584 404569 115612 405622
rect 115846 405583 115902 405592
rect 115860 405006 115888 405583
rect 115848 405000 115900 405006
rect 115848 404942 115900 404948
rect 115570 404560 115626 404569
rect 115570 404495 115626 404504
rect 115846 403472 115902 403481
rect 115846 403407 115902 403416
rect 115860 403306 115888 403407
rect 115848 403300 115900 403306
rect 115848 403242 115900 403248
rect 115662 401296 115718 401305
rect 115662 401231 115718 401240
rect 115018 400480 115074 400489
rect 115018 400415 115020 400424
rect 115072 400415 115074 400424
rect 115020 400386 115072 400392
rect 115676 400246 115704 401231
rect 115664 400240 115716 400246
rect 115664 400182 115716 400188
rect 115202 399392 115258 399401
rect 115202 399327 115258 399336
rect 114928 398132 114980 398138
rect 114928 398074 114980 398080
rect 114940 389842 114968 398074
rect 114928 389836 114980 389842
rect 114928 389778 114980 389784
rect 115216 327214 115244 399327
rect 115846 398304 115902 398313
rect 115846 398239 115902 398248
rect 115860 398138 115888 398239
rect 115848 398132 115900 398138
rect 115848 398074 115900 398080
rect 115846 397216 115902 397225
rect 115846 397151 115902 397160
rect 115860 396778 115888 397151
rect 115848 396772 115900 396778
rect 115848 396714 115900 396720
rect 115846 396400 115902 396409
rect 115846 396335 115902 396344
rect 115860 396098 115888 396335
rect 115848 396092 115900 396098
rect 115848 396034 115900 396040
rect 115846 395312 115902 395321
rect 115846 395247 115902 395256
rect 115860 394738 115888 395247
rect 115848 394732 115900 394738
rect 115848 394674 115900 394680
rect 115570 394224 115626 394233
rect 115570 394159 115626 394168
rect 115584 393378 115612 394159
rect 115572 393372 115624 393378
rect 115572 393314 115624 393320
rect 115848 393168 115900 393174
rect 115846 393136 115848 393145
rect 115900 393136 115902 393145
rect 115846 393071 115902 393080
rect 115846 392048 115902 392057
rect 115846 391983 115848 391992
rect 115900 391983 115902 391992
rect 115848 391954 115900 391960
rect 115952 386306 115980 550598
rect 116596 536761 116624 702782
rect 118700 576904 118752 576910
rect 118700 576846 118752 576852
rect 116582 536752 116638 536761
rect 116582 536687 116638 536696
rect 118712 527882 118740 576846
rect 119356 536110 119384 703122
rect 132592 590708 132644 590714
rect 132592 590650 132644 590656
rect 125600 587172 125652 587178
rect 125600 587114 125652 587120
rect 121736 585812 121788 585818
rect 121736 585754 121788 585760
rect 121748 585206 121776 585754
rect 121460 585200 121512 585206
rect 121460 585142 121512 585148
rect 121736 585200 121788 585206
rect 121736 585142 121788 585148
rect 119344 536104 119396 536110
rect 119344 536046 119396 536052
rect 118700 527876 118752 527882
rect 118700 527818 118752 527824
rect 116124 468512 116176 468518
rect 116124 468454 116176 468460
rect 116032 436756 116084 436762
rect 116032 436698 116084 436704
rect 116044 436150 116072 436698
rect 116032 436144 116084 436150
rect 116032 436086 116084 436092
rect 115940 386300 115992 386306
rect 115940 386242 115992 386248
rect 115940 380180 115992 380186
rect 115940 380122 115992 380128
rect 115204 327208 115256 327214
rect 115204 327150 115256 327156
rect 114742 318200 114798 318209
rect 114742 318135 114798 318144
rect 114650 307864 114706 307873
rect 114650 307799 114706 307808
rect 114650 285968 114706 285977
rect 114650 285903 114706 285912
rect 114558 283520 114614 283529
rect 114558 283455 114614 283464
rect 114468 233912 114520 233918
rect 114468 233854 114520 233860
rect 114572 214674 114600 283455
rect 114664 248470 114692 285903
rect 115018 263664 115074 263673
rect 115018 263599 115074 263608
rect 115032 263566 115060 263599
rect 115020 263560 115072 263566
rect 115020 263502 115072 263508
rect 115032 262954 115060 263502
rect 115020 262948 115072 262954
rect 115020 262890 115072 262896
rect 115216 260778 115244 327150
rect 115846 285968 115902 285977
rect 115846 285903 115902 285912
rect 115860 285734 115888 285903
rect 115848 285728 115900 285734
rect 115848 285670 115900 285676
rect 115388 266416 115440 266422
rect 115388 266358 115440 266364
rect 115204 260772 115256 260778
rect 115204 260714 115256 260720
rect 114836 250504 114888 250510
rect 114836 250446 114888 250452
rect 114652 248464 114704 248470
rect 114652 248406 114704 248412
rect 114744 238060 114796 238066
rect 114744 238002 114796 238008
rect 114650 234560 114706 234569
rect 114650 234495 114706 234504
rect 114664 233306 114692 234495
rect 114652 233300 114704 233306
rect 114652 233242 114704 233248
rect 114560 214668 114612 214674
rect 114560 214610 114612 214616
rect 114558 206408 114614 206417
rect 114558 206343 114614 206352
rect 114468 164892 114520 164898
rect 114468 164834 114520 164840
rect 113364 138780 113416 138786
rect 113364 138722 113416 138728
rect 113272 121440 113324 121446
rect 113272 121382 113324 121388
rect 113180 108996 113232 109002
rect 113180 108938 113232 108944
rect 111984 108928 112036 108934
rect 111984 108870 112036 108876
rect 111892 97980 111944 97986
rect 111892 97922 111944 97928
rect 111800 88324 111852 88330
rect 111800 88266 111852 88272
rect 111812 87650 111840 88266
rect 111800 87644 111852 87650
rect 111800 87586 111852 87592
rect 111628 6886 111748 6914
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 110510 3496 110566 3505
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 110510 3431 110566 3440
rect 109314 3360 109370 3369
rect 109314 3295 109370 3304
rect 109328 480 109356 3295
rect 110524 480 110552 3431
rect 111628 480 111656 6886
rect 114480 3534 114508 164834
rect 114572 92313 114600 206343
rect 114652 193860 114704 193866
rect 114652 193802 114704 193808
rect 114558 92304 114614 92313
rect 114558 92239 114614 92248
rect 114664 86873 114692 193802
rect 114756 140826 114784 238002
rect 114848 229838 114876 250446
rect 114836 229832 114888 229838
rect 114836 229774 114888 229780
rect 115400 198014 115428 266358
rect 115952 240854 115980 380122
rect 116044 291854 116072 436086
rect 116136 402393 116164 468454
rect 117412 456068 117464 456074
rect 117412 456010 117464 456016
rect 117318 443048 117374 443057
rect 117318 442983 117374 442992
rect 116216 439544 116268 439550
rect 116216 439486 116268 439492
rect 116228 415750 116256 439486
rect 116216 415744 116268 415750
rect 116216 415686 116268 415692
rect 116122 402384 116178 402393
rect 116122 402319 116178 402328
rect 116136 371210 116164 402319
rect 116228 378826 116256 415686
rect 116216 378820 116268 378826
rect 116216 378762 116268 378768
rect 116124 371204 116176 371210
rect 116124 371146 116176 371152
rect 117332 367810 117360 442983
rect 117424 391270 117452 456010
rect 117502 439512 117558 439521
rect 117502 439447 117558 439456
rect 117516 410582 117544 439447
rect 117504 410576 117556 410582
rect 117504 410518 117556 410524
rect 118608 403300 118660 403306
rect 118608 403242 118660 403248
rect 118620 402286 118648 403242
rect 118608 402280 118660 402286
rect 118608 402222 118660 402228
rect 117504 400444 117556 400450
rect 117504 400386 117556 400392
rect 117412 391264 117464 391270
rect 117412 391206 117464 391212
rect 117516 383625 117544 400386
rect 118712 393174 118740 527818
rect 118792 485104 118844 485110
rect 118792 485046 118844 485052
rect 118804 427854 118832 485046
rect 120172 474020 120224 474026
rect 120172 473962 120224 473968
rect 118976 464364 119028 464370
rect 118976 464306 119028 464312
rect 118884 437572 118936 437578
rect 118884 437514 118936 437520
rect 118792 427848 118844 427854
rect 118792 427790 118844 427796
rect 118792 426420 118844 426426
rect 118792 426362 118844 426368
rect 118804 425134 118832 426362
rect 118792 425128 118844 425134
rect 118792 425070 118844 425076
rect 118700 393168 118752 393174
rect 118700 393110 118752 393116
rect 118712 392086 118740 393110
rect 118700 392080 118752 392086
rect 118700 392022 118752 392028
rect 117502 383616 117558 383625
rect 117502 383551 117558 383560
rect 117412 381608 117464 381614
rect 117412 381550 117464 381556
rect 117320 367804 117372 367810
rect 117320 367746 117372 367752
rect 116124 326392 116176 326398
rect 116124 326334 116176 326340
rect 116136 325786 116164 326334
rect 116124 325780 116176 325786
rect 116124 325722 116176 325728
rect 116032 291848 116084 291854
rect 116030 291816 116032 291825
rect 116084 291816 116086 291825
rect 116030 291751 116086 291760
rect 116030 287328 116086 287337
rect 116030 287263 116086 287272
rect 115940 240848 115992 240854
rect 115940 240790 115992 240796
rect 115940 233912 115992 233918
rect 115940 233854 115992 233860
rect 115952 224942 115980 233854
rect 115940 224936 115992 224942
rect 115940 224878 115992 224884
rect 115846 224224 115902 224233
rect 115846 224159 115902 224168
rect 115756 215280 115808 215286
rect 115756 215222 115808 215228
rect 115768 214674 115796 215222
rect 115756 214668 115808 214674
rect 115756 214610 115808 214616
rect 115388 198008 115440 198014
rect 115388 197950 115440 197956
rect 114744 140820 114796 140826
rect 114744 140762 114796 140768
rect 114650 86864 114706 86873
rect 114650 86799 114706 86808
rect 115754 86864 115810 86873
rect 115754 86799 115810 86808
rect 115768 86193 115796 86799
rect 115754 86184 115810 86193
rect 115754 86119 115810 86128
rect 115860 3534 115888 224159
rect 115952 88262 115980 224878
rect 116044 214606 116072 287263
rect 116136 284209 116164 325722
rect 117320 313336 117372 313342
rect 117320 313278 117372 313284
rect 116582 288552 116638 288561
rect 116582 288487 116638 288496
rect 116596 288454 116624 288487
rect 116584 288448 116636 288454
rect 116584 288390 116636 288396
rect 116122 284200 116178 284209
rect 116122 284135 116178 284144
rect 116032 214600 116084 214606
rect 116032 214542 116084 214548
rect 116596 156670 116624 288390
rect 116860 273216 116912 273222
rect 116860 273158 116912 273164
rect 116872 272542 116900 273158
rect 116860 272536 116912 272542
rect 116860 272478 116912 272484
rect 116872 271969 116900 272478
rect 116858 271960 116914 271969
rect 116858 271895 116914 271904
rect 116676 268932 116728 268938
rect 116676 268874 116728 268880
rect 116584 156664 116636 156670
rect 116584 156606 116636 156612
rect 116688 145586 116716 268874
rect 117228 241460 117280 241466
rect 117228 241402 117280 241408
rect 117240 240854 117268 241402
rect 117228 240848 117280 240854
rect 117228 240790 117280 240796
rect 117228 215212 117280 215218
rect 117228 215154 117280 215160
rect 117240 214606 117268 215154
rect 117228 214600 117280 214606
rect 117228 214542 117280 214548
rect 116768 211812 116820 211818
rect 116768 211754 116820 211760
rect 116780 195974 116808 211754
rect 116768 195968 116820 195974
rect 116768 195910 116820 195916
rect 116676 145580 116728 145586
rect 116676 145522 116728 145528
rect 116780 111081 116808 195910
rect 117332 138689 117360 313278
rect 117424 206961 117452 381550
rect 117964 366376 118016 366382
rect 117964 366318 118016 366324
rect 117780 313948 117832 313954
rect 117780 313890 117832 313896
rect 117792 313342 117820 313890
rect 117780 313336 117832 313342
rect 117780 313278 117832 313284
rect 117976 242962 118004 366318
rect 118056 301504 118108 301510
rect 118056 301446 118108 301452
rect 118068 258738 118096 301446
rect 118804 276049 118832 425070
rect 118896 362234 118924 437514
rect 118988 422006 119016 464306
rect 120078 437608 120134 437617
rect 120078 437543 120134 437552
rect 118976 422000 119028 422006
rect 118976 421942 119028 421948
rect 118988 421598 119016 421942
rect 118976 421592 119028 421598
rect 118976 421534 119028 421540
rect 119344 415404 119396 415410
rect 119344 415346 119396 415352
rect 119356 414934 119384 415346
rect 119344 414928 119396 414934
rect 119344 414870 119396 414876
rect 119068 363656 119120 363662
rect 119068 363598 119120 363604
rect 118884 362228 118936 362234
rect 118884 362170 118936 362176
rect 118882 320920 118938 320929
rect 118882 320855 118938 320864
rect 118896 320278 118924 320855
rect 118884 320272 118936 320278
rect 118884 320214 118936 320220
rect 118790 276040 118846 276049
rect 118790 275975 118846 275984
rect 118804 274689 118832 275975
rect 118790 274680 118846 274689
rect 118790 274615 118846 274624
rect 118896 268938 118924 320214
rect 118976 276684 119028 276690
rect 118976 276626 119028 276632
rect 118884 268932 118936 268938
rect 118884 268874 118936 268880
rect 118792 263560 118844 263566
rect 118792 263502 118844 263508
rect 118056 258732 118108 258738
rect 118056 258674 118108 258680
rect 117964 242956 118016 242962
rect 117964 242898 118016 242904
rect 117976 237969 118004 242898
rect 117962 237960 118018 237969
rect 117962 237895 118018 237904
rect 117686 235376 117742 235385
rect 117686 235311 117742 235320
rect 117700 234598 117728 235311
rect 117688 234592 117740 234598
rect 117688 234534 117740 234540
rect 117964 234592 118016 234598
rect 117964 234534 118016 234540
rect 117410 206952 117466 206961
rect 117410 206887 117466 206896
rect 117424 206417 117452 206887
rect 117410 206408 117466 206417
rect 117410 206343 117466 206352
rect 117318 138680 117374 138689
rect 117318 138615 117374 138624
rect 116766 111072 116822 111081
rect 116766 111007 116822 111016
rect 117976 90914 118004 234534
rect 118700 209160 118752 209166
rect 118700 209102 118752 209108
rect 118608 189780 118660 189786
rect 118608 189722 118660 189728
rect 117964 90908 118016 90914
rect 117964 90850 118016 90856
rect 115940 88256 115992 88262
rect 115940 88198 115992 88204
rect 116398 3632 116454 3641
rect 116398 3567 116454 3576
rect 114008 3528 114060 3534
rect 112810 3496 112866 3505
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 112810 3431 112866 3440
rect 112824 480 112852 3431
rect 114020 480 114048 3470
rect 115216 480 115244 3470
rect 116412 480 116440 3567
rect 118620 3534 118648 189722
rect 118712 89690 118740 209102
rect 118804 115870 118832 263502
rect 118988 242214 119016 276626
rect 118976 242208 119028 242214
rect 118976 242150 119028 242156
rect 119080 208321 119108 363598
rect 119356 325009 119384 414870
rect 119342 325000 119398 325009
rect 119342 324935 119398 324944
rect 119344 321972 119396 321978
rect 119344 321914 119396 321920
rect 119356 287706 119384 321914
rect 120092 320793 120120 437543
rect 120184 415410 120212 473962
rect 120356 450560 120408 450566
rect 120356 450502 120408 450508
rect 120264 433288 120316 433294
rect 120264 433230 120316 433236
rect 120172 415404 120224 415410
rect 120172 415346 120224 415352
rect 120276 377466 120304 433230
rect 120368 412078 120396 450502
rect 120356 412072 120408 412078
rect 120356 412014 120408 412020
rect 121472 389314 121500 585142
rect 122838 582448 122894 582457
rect 122838 582383 122894 582392
rect 121644 457496 121696 457502
rect 121644 457438 121696 457444
rect 121552 427848 121604 427854
rect 121552 427790 121604 427796
rect 121380 389286 121500 389314
rect 121380 388906 121408 389286
rect 121460 389156 121512 389162
rect 121460 389098 121512 389104
rect 121472 389065 121500 389098
rect 121458 389056 121514 389065
rect 121458 388991 121514 389000
rect 121380 388878 121500 388906
rect 121472 387802 121500 388878
rect 120724 387796 120776 387802
rect 120724 387738 120776 387744
rect 121460 387796 121512 387802
rect 121460 387738 121512 387744
rect 120736 387122 120764 387738
rect 120724 387116 120776 387122
rect 120724 387058 120776 387064
rect 120264 377460 120316 377466
rect 120264 377402 120316 377408
rect 120172 333260 120224 333266
rect 120172 333202 120224 333208
rect 120184 332654 120212 333202
rect 120172 332648 120224 332654
rect 120172 332590 120224 332596
rect 120078 320784 120134 320793
rect 120078 320719 120134 320728
rect 119344 287700 119396 287706
rect 119344 287642 119396 287648
rect 120184 282985 120212 332590
rect 120170 282976 120226 282985
rect 120170 282911 120226 282920
rect 119436 267028 119488 267034
rect 119436 266970 119488 266976
rect 119344 238060 119396 238066
rect 119344 238002 119396 238008
rect 119066 208312 119122 208321
rect 119066 208247 119122 208256
rect 119080 207641 119108 208247
rect 119066 207632 119122 207641
rect 119066 207567 119122 207576
rect 118792 115864 118844 115870
rect 118792 115806 118844 115812
rect 118700 89684 118752 89690
rect 118700 89626 118752 89632
rect 119356 3602 119384 238002
rect 119448 228614 119476 266970
rect 120080 263628 120132 263634
rect 120080 263570 120132 263576
rect 119436 228608 119488 228614
rect 119436 228550 119488 228556
rect 120092 117298 120120 263570
rect 120172 246356 120224 246362
rect 120172 246298 120224 246304
rect 120184 246265 120212 246298
rect 120170 246256 120226 246265
rect 120170 246191 120226 246200
rect 120080 117292 120132 117298
rect 120080 117234 120132 117240
rect 120184 102814 120212 246191
rect 120264 228608 120316 228614
rect 120264 228550 120316 228556
rect 120276 228342 120304 228550
rect 120264 228336 120316 228342
rect 120264 228278 120316 228284
rect 120276 121553 120304 228278
rect 120736 211041 120764 387058
rect 121460 365016 121512 365022
rect 121460 364958 121512 364964
rect 120908 302252 120960 302258
rect 120908 302194 120960 302200
rect 120816 294636 120868 294642
rect 120816 294578 120868 294584
rect 120828 252550 120856 294578
rect 120920 291854 120948 302194
rect 120908 291848 120960 291854
rect 120908 291790 120960 291796
rect 120908 289944 120960 289950
rect 120908 289886 120960 289892
rect 120920 281586 120948 289886
rect 120908 281580 120960 281586
rect 120908 281522 120960 281528
rect 120920 266422 120948 281522
rect 120908 266416 120960 266422
rect 120908 266358 120960 266364
rect 120816 252544 120868 252550
rect 120816 252486 120868 252492
rect 120354 211032 120410 211041
rect 120354 210967 120410 210976
rect 120722 211032 120778 211041
rect 120722 210967 120778 210976
rect 120368 210361 120396 210967
rect 120354 210352 120410 210361
rect 120354 210287 120410 210296
rect 121472 206281 121500 364958
rect 121564 275913 121592 427790
rect 121656 422958 121684 457438
rect 122852 426426 122880 582383
rect 122932 438932 122984 438938
rect 122932 438874 122984 438880
rect 122840 426420 122892 426426
rect 122840 426362 122892 426368
rect 121644 422952 121696 422958
rect 121644 422894 121696 422900
rect 121644 416832 121696 416838
rect 121644 416774 121696 416780
rect 121656 304201 121684 416774
rect 122840 392080 122892 392086
rect 122840 392022 122892 392028
rect 122852 306338 122880 392022
rect 122944 345014 122972 438874
rect 123024 437504 123076 437510
rect 123024 437446 123076 437452
rect 123036 376106 123064 437446
rect 123484 436212 123536 436218
rect 123484 436154 123536 436160
rect 123024 376100 123076 376106
rect 123024 376042 123076 376048
rect 122944 344986 123064 345014
rect 122932 334620 122984 334626
rect 122932 334562 122984 334568
rect 122944 325694 122972 334562
rect 123036 329118 123064 344986
rect 123496 343738 123524 436154
rect 124402 434752 124458 434761
rect 124402 434687 124458 434696
rect 124220 431996 124272 432002
rect 124220 431938 124272 431944
rect 124128 396772 124180 396778
rect 124128 396714 124180 396720
rect 124140 396681 124168 396714
rect 124126 396672 124182 396681
rect 124126 396607 124182 396616
rect 123484 343732 123536 343738
rect 123484 343674 123536 343680
rect 123024 329112 123076 329118
rect 123024 329054 123076 329060
rect 122944 325666 123064 325694
rect 122840 306332 122892 306338
rect 122840 306274 122892 306280
rect 122852 305658 122880 306274
rect 122840 305652 122892 305658
rect 122840 305594 122892 305600
rect 121642 304192 121698 304201
rect 121642 304127 121698 304136
rect 122102 292632 122158 292641
rect 122102 292567 122158 292576
rect 121642 291272 121698 291281
rect 121642 291207 121698 291216
rect 121550 275904 121606 275913
rect 121550 275839 121606 275848
rect 121564 274689 121592 275839
rect 121550 274680 121606 274689
rect 121550 274615 121606 274624
rect 121458 206272 121514 206281
rect 121458 206207 121514 206216
rect 121656 141409 121684 291207
rect 122116 244934 122144 292567
rect 122840 271924 122892 271930
rect 122840 271866 122892 271872
rect 122196 249076 122248 249082
rect 122196 249018 122248 249024
rect 122104 244928 122156 244934
rect 122104 244870 122156 244876
rect 122208 234598 122236 249018
rect 122196 234592 122248 234598
rect 122196 234534 122248 234540
rect 122104 233912 122156 233918
rect 122104 233854 122156 233860
rect 121642 141400 121698 141409
rect 121642 141335 121698 141344
rect 120262 121544 120318 121553
rect 120262 121479 120318 121488
rect 120172 102808 120224 102814
rect 120172 102750 120224 102756
rect 119988 89004 120040 89010
rect 119988 88946 120040 88952
rect 120000 6914 120028 88946
rect 119908 6886 120028 6914
rect 119344 3596 119396 3602
rect 119344 3538 119396 3544
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 117608 480 117636 3470
rect 118792 3460 118844 3466
rect 118792 3402 118844 3408
rect 118804 480 118832 3402
rect 119908 480 119936 6886
rect 122116 3534 122144 233854
rect 122748 229152 122800 229158
rect 122748 229094 122800 229100
rect 122760 201482 122788 229094
rect 122196 201476 122248 201482
rect 122196 201418 122248 201424
rect 122748 201476 122800 201482
rect 122748 201418 122800 201424
rect 122208 133890 122236 201418
rect 122196 133884 122248 133890
rect 122196 133826 122248 133832
rect 122852 125594 122880 271866
rect 123036 254590 123064 325666
rect 123496 321978 123524 343674
rect 123852 334620 123904 334626
rect 123852 334562 123904 334568
rect 123864 334082 123892 334562
rect 123852 334076 123904 334082
rect 123852 334018 123904 334024
rect 123484 321972 123536 321978
rect 123484 321914 123536 321920
rect 123484 307896 123536 307902
rect 123484 307838 123536 307844
rect 123116 307760 123168 307766
rect 123116 307702 123168 307708
rect 123128 306406 123156 307702
rect 123116 306400 123168 306406
rect 123116 306342 123168 306348
rect 123024 254584 123076 254590
rect 123024 254526 123076 254532
rect 122930 234560 122986 234569
rect 122930 234495 122986 234504
rect 122944 233889 122972 234495
rect 122930 233880 122986 233889
rect 122930 233815 122986 233824
rect 122840 125588 122892 125594
rect 122840 125530 122892 125536
rect 122944 118658 122972 233815
rect 123128 229158 123156 306342
rect 123116 229152 123168 229158
rect 123116 229094 123168 229100
rect 122932 118652 122984 118658
rect 122932 118594 122984 118600
rect 123496 4146 123524 307838
rect 124232 307766 124260 431938
rect 124312 373312 124364 373318
rect 124312 373254 124364 373260
rect 124220 307760 124272 307766
rect 124220 307702 124272 307708
rect 124324 249082 124352 373254
rect 124416 359514 124444 434687
rect 125612 402974 125640 587114
rect 126980 581120 127032 581126
rect 126980 581062 127032 581068
rect 125876 461644 125928 461650
rect 125876 461586 125928 461592
rect 125784 440292 125836 440298
rect 125784 440234 125836 440240
rect 125612 402946 125732 402974
rect 125704 398138 125732 402946
rect 125692 398132 125744 398138
rect 125692 398074 125744 398080
rect 124404 359508 124456 359514
rect 124404 359450 124456 359456
rect 124402 322144 124458 322153
rect 124402 322079 124458 322088
rect 125506 322144 125562 322153
rect 125506 322079 125562 322088
rect 124416 262886 124444 322079
rect 125520 321706 125548 322079
rect 125508 321700 125560 321706
rect 125508 321642 125560 321648
rect 125598 312080 125654 312089
rect 125598 312015 125654 312024
rect 124864 294024 124916 294030
rect 124864 293966 124916 293972
rect 124404 262880 124456 262886
rect 124404 262822 124456 262828
rect 124312 249076 124364 249082
rect 124312 249018 124364 249024
rect 124220 247716 124272 247722
rect 124220 247658 124272 247664
rect 124232 202162 124260 247658
rect 124310 244352 124366 244361
rect 124310 244287 124312 244296
rect 124364 244287 124366 244296
rect 124312 244258 124364 244264
rect 124324 212537 124352 244258
rect 124310 212528 124366 212537
rect 124310 212463 124366 212472
rect 124220 202156 124272 202162
rect 124220 202098 124272 202104
rect 123576 119400 123628 119406
rect 123576 119342 123628 119348
rect 123588 78062 123616 119342
rect 124232 102066 124260 202098
rect 124876 137290 124904 293966
rect 125508 293276 125560 293282
rect 125508 293218 125560 293224
rect 125520 258058 125548 293218
rect 125508 258052 125560 258058
rect 125508 257994 125560 258000
rect 125520 256766 125548 257994
rect 125508 256760 125560 256766
rect 125508 256702 125560 256708
rect 125508 217320 125560 217326
rect 125508 217262 125560 217268
rect 124864 137284 124916 137290
rect 124864 137226 124916 137232
rect 124220 102060 124272 102066
rect 124220 102002 124272 102008
rect 123576 78056 123628 78062
rect 123576 77998 123628 78004
rect 122288 4140 122340 4146
rect 122288 4082 122340 4088
rect 123484 4140 123536 4146
rect 123484 4082 123536 4088
rect 121092 3528 121144 3534
rect 121092 3470 121144 3476
rect 122104 3528 122156 3534
rect 122104 3470 122156 3476
rect 121104 480 121132 3470
rect 122300 480 122328 4082
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 123496 480 123524 3538
rect 125520 3534 125548 217262
rect 125612 140049 125640 312015
rect 125704 226302 125732 398074
rect 125796 313954 125824 440234
rect 125888 385014 125916 461586
rect 126992 405006 127020 581062
rect 128360 561740 128412 561746
rect 128360 561682 128412 561688
rect 128372 413982 128400 561682
rect 128452 441652 128504 441658
rect 128452 441594 128504 441600
rect 128360 413976 128412 413982
rect 128360 413918 128412 413924
rect 128372 413302 128400 413918
rect 128360 413296 128412 413302
rect 128360 413238 128412 413244
rect 127072 410576 127124 410582
rect 127072 410518 127124 410524
rect 126980 405000 127032 405006
rect 126980 404942 127032 404948
rect 125876 385008 125928 385014
rect 125876 384950 125928 384956
rect 126888 385008 126940 385014
rect 126888 384950 126940 384956
rect 126900 383761 126928 384950
rect 126886 383752 126942 383761
rect 126886 383687 126942 383696
rect 126980 382968 127032 382974
rect 126980 382910 127032 382916
rect 126244 370524 126296 370530
rect 126244 370466 126296 370472
rect 125784 313948 125836 313954
rect 125784 313890 125836 313896
rect 126256 305454 126284 370466
rect 126244 305448 126296 305454
rect 126244 305390 126296 305396
rect 126244 282940 126296 282946
rect 126244 282882 126296 282888
rect 125782 251832 125838 251841
rect 125782 251767 125838 251776
rect 125692 226296 125744 226302
rect 125692 226238 125744 226244
rect 125704 225622 125732 226238
rect 125692 225616 125744 225622
rect 125692 225558 125744 225564
rect 125690 218648 125746 218657
rect 125690 218583 125746 218592
rect 125598 140040 125654 140049
rect 125598 139975 125654 139984
rect 125704 112470 125732 218583
rect 125692 112464 125744 112470
rect 125692 112406 125744 112412
rect 125796 106282 125824 251767
rect 126256 241369 126284 282882
rect 126242 241360 126298 241369
rect 126242 241295 126298 241304
rect 126886 222048 126942 222057
rect 126886 221983 126942 221992
rect 126244 221468 126296 221474
rect 126244 221410 126296 221416
rect 125784 106276 125836 106282
rect 125784 106218 125836 106224
rect 125600 17264 125652 17270
rect 125600 17206 125652 17212
rect 125612 16574 125640 17206
rect 125612 16546 125916 16574
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 124692 480 124720 3470
rect 125888 480 125916 16546
rect 126256 3505 126284 221410
rect 126900 220862 126928 221983
rect 126888 220856 126940 220862
rect 126888 220798 126940 220804
rect 126992 205562 127020 382910
rect 127084 264246 127112 410518
rect 127440 405000 127492 405006
rect 127440 404942 127492 404948
rect 127452 403646 127480 404942
rect 127440 403640 127492 403646
rect 127440 403582 127492 403588
rect 128360 391264 128412 391270
rect 128360 391206 128412 391212
rect 127164 276752 127216 276758
rect 127164 276694 127216 276700
rect 127072 264240 127124 264246
rect 127072 264182 127124 264188
rect 127084 263673 127112 264182
rect 127070 263664 127126 263673
rect 127070 263599 127126 263608
rect 127072 256760 127124 256766
rect 127072 256702 127124 256708
rect 126980 205556 127032 205562
rect 126980 205498 127032 205504
rect 126992 204950 127020 205498
rect 126980 204944 127032 204950
rect 126980 204886 127032 204892
rect 127084 110362 127112 256702
rect 127176 129674 127204 276694
rect 127256 213240 127308 213246
rect 127256 213182 127308 213188
rect 127164 129668 127216 129674
rect 127164 129610 127216 129616
rect 127072 110356 127124 110362
rect 127072 110298 127124 110304
rect 127084 109750 127112 110298
rect 127072 109744 127124 109750
rect 127072 109686 127124 109692
rect 127268 95577 127296 213182
rect 128372 208185 128400 391206
rect 128464 309097 128492 441594
rect 132500 433356 132552 433362
rect 132500 433298 132552 433304
rect 129740 412072 129792 412078
rect 129740 412014 129792 412020
rect 129004 324964 129056 324970
rect 129004 324906 129056 324912
rect 128450 309088 128506 309097
rect 128450 309023 128506 309032
rect 128464 308417 128492 309023
rect 128450 308408 128506 308417
rect 128450 308343 128506 308352
rect 128544 305448 128596 305454
rect 128544 305390 128596 305396
rect 128452 281580 128504 281586
rect 128452 281522 128504 281528
rect 128464 278730 128492 281522
rect 128452 278724 128504 278730
rect 128452 278666 128504 278672
rect 128452 274032 128504 274038
rect 128452 273974 128504 273980
rect 128464 273902 128492 273974
rect 128452 273896 128504 273902
rect 128452 273838 128504 273844
rect 128358 208176 128414 208185
rect 128358 208111 128414 208120
rect 128372 207777 128400 208111
rect 128358 207768 128414 207777
rect 128358 207703 128414 207712
rect 128360 207664 128412 207670
rect 128360 207606 128412 207612
rect 127254 95568 127310 95577
rect 127254 95503 127310 95512
rect 128372 93838 128400 207606
rect 128464 124914 128492 273838
rect 128556 240038 128584 305390
rect 129016 273902 129044 324906
rect 129004 273896 129056 273902
rect 129004 273838 129056 273844
rect 129004 253224 129056 253230
rect 129004 253166 129056 253172
rect 128544 240032 128596 240038
rect 128544 239974 128596 239980
rect 128556 239426 128584 239974
rect 128544 239420 128596 239426
rect 128544 239362 128596 239368
rect 129016 227730 129044 253166
rect 129752 234569 129780 412014
rect 131120 396092 131172 396098
rect 131120 396034 131172 396040
rect 130568 274712 130620 274718
rect 130568 274654 130620 274660
rect 130384 271176 130436 271182
rect 130384 271118 130436 271124
rect 129738 234560 129794 234569
rect 129738 234495 129794 234504
rect 129738 232656 129794 232665
rect 129738 232591 129794 232600
rect 129004 227724 129056 227730
rect 129004 227666 129056 227672
rect 129016 226370 129044 227666
rect 128544 226364 128596 226370
rect 128544 226306 128596 226312
rect 129004 226364 129056 226370
rect 129004 226306 129056 226312
rect 128452 124908 128504 124914
rect 128452 124850 128504 124856
rect 128360 93832 128412 93838
rect 128360 93774 128412 93780
rect 128556 84182 128584 226306
rect 128636 212424 128688 212430
rect 128636 212366 128688 212372
rect 128648 211857 128676 212366
rect 128634 211848 128690 211857
rect 128634 211783 128690 211792
rect 129004 201544 129056 201550
rect 129004 201486 129056 201492
rect 129016 108361 129044 201486
rect 129752 113150 129780 232591
rect 130396 124166 130424 271118
rect 130476 257372 130528 257378
rect 130476 257314 130528 257320
rect 130488 223582 130516 257314
rect 130580 250510 130608 274654
rect 130568 250504 130620 250510
rect 130568 250446 130620 250452
rect 130476 223576 130528 223582
rect 130476 223518 130528 223524
rect 131028 223576 131080 223582
rect 131028 223518 131080 223524
rect 130384 124160 130436 124166
rect 130384 124102 130436 124108
rect 130568 124160 130620 124166
rect 130568 124102 130620 124108
rect 130580 123486 130608 124102
rect 130568 123480 130620 123486
rect 130568 123422 130620 123428
rect 129740 113144 129792 113150
rect 129740 113086 129792 113092
rect 129002 108352 129058 108361
rect 129002 108287 129058 108296
rect 130200 100700 130252 100706
rect 130200 100642 130252 100648
rect 130212 100026 130240 100642
rect 131040 100026 131068 223518
rect 131132 219201 131160 396034
rect 131764 291236 131816 291242
rect 131764 291178 131816 291184
rect 131212 278044 131264 278050
rect 131212 277986 131264 277992
rect 131118 219192 131174 219201
rect 131118 219127 131174 219136
rect 131132 218657 131160 219127
rect 131118 218648 131174 218657
rect 131118 218583 131174 218592
rect 131224 129742 131252 277986
rect 131776 269074 131804 291178
rect 131764 269068 131816 269074
rect 131764 269010 131816 269016
rect 131304 249144 131356 249150
rect 131304 249086 131356 249092
rect 131212 129736 131264 129742
rect 131212 129678 131264 129684
rect 131316 102134 131344 249086
rect 131764 224256 131816 224262
rect 131764 224198 131816 224204
rect 131776 132462 131804 224198
rect 131764 132456 131816 132462
rect 131764 132398 131816 132404
rect 131304 102128 131356 102134
rect 131304 102070 131356 102076
rect 131316 101454 131344 102070
rect 131304 101448 131356 101454
rect 131304 101390 131356 101396
rect 130200 100020 130252 100026
rect 130200 99962 130252 99968
rect 131028 100020 131080 100026
rect 131028 99962 131080 99968
rect 128544 84176 128596 84182
rect 128544 84118 128596 84124
rect 129004 61396 129056 61402
rect 129004 61338 129056 61344
rect 129016 7614 129044 61338
rect 132512 16574 132540 433298
rect 132604 405686 132632 590650
rect 133880 569220 133932 569226
rect 133880 569162 133932 569168
rect 132592 405680 132644 405686
rect 132592 405622 132644 405628
rect 133788 405680 133840 405686
rect 133788 405622 133840 405628
rect 133800 405006 133828 405622
rect 133788 405000 133840 405006
rect 133788 404942 133840 404948
rect 132590 396672 132646 396681
rect 132590 396607 132646 396616
rect 132604 258777 132632 396607
rect 133892 386374 133920 569162
rect 136652 538286 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 703322 154160 703520
rect 154120 703316 154172 703322
rect 154120 703258 154172 703264
rect 170324 703118 170352 703520
rect 170312 703112 170364 703118
rect 170312 703054 170364 703060
rect 202800 703050 202828 703520
rect 218992 703186 219020 703520
rect 235184 703254 235212 703520
rect 235172 703248 235224 703254
rect 235172 703190 235224 703196
rect 218980 703180 219032 703186
rect 218980 703122 219032 703128
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 267660 697610 267688 703520
rect 271144 703180 271196 703186
rect 271144 703122 271196 703128
rect 268384 703044 268436 703050
rect 268384 702986 268436 702992
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 136640 538280 136692 538286
rect 136640 538222 136692 538228
rect 136732 440360 136784 440366
rect 136732 440302 136784 440308
rect 134524 434784 134576 434790
rect 134524 434726 134576 434732
rect 133880 386368 133932 386374
rect 133880 386310 133932 386316
rect 134536 325694 134564 434726
rect 135260 430636 135312 430642
rect 135260 430578 135312 430584
rect 134536 325666 134656 325694
rect 134628 314770 134656 325666
rect 134616 314764 134668 314770
rect 134616 314706 134668 314712
rect 134524 299532 134576 299538
rect 134524 299474 134576 299480
rect 133788 265668 133840 265674
rect 133788 265610 133840 265616
rect 133800 264994 133828 265610
rect 133144 264988 133196 264994
rect 133144 264930 133196 264936
rect 133788 264988 133840 264994
rect 133788 264930 133840 264936
rect 132590 258768 132646 258777
rect 132590 258703 132646 258712
rect 132592 249824 132644 249830
rect 132592 249766 132644 249772
rect 132604 201550 132632 249766
rect 132592 201544 132644 201550
rect 132592 201486 132644 201492
rect 133156 115938 133184 264930
rect 134536 261526 134564 299474
rect 134628 280838 134656 314706
rect 134616 280832 134668 280838
rect 134616 280774 134668 280780
rect 135272 278769 135300 430578
rect 136640 386368 136692 386374
rect 136640 386310 136692 386316
rect 135258 278760 135314 278769
rect 135258 278695 135314 278704
rect 135272 277394 135300 278695
rect 135272 277366 135484 277394
rect 135260 273964 135312 273970
rect 135260 273906 135312 273912
rect 134524 261520 134576 261526
rect 134524 261462 134576 261468
rect 135168 260160 135220 260166
rect 135168 260102 135220 260108
rect 135180 259486 135208 260102
rect 133972 259480 134024 259486
rect 133972 259422 134024 259428
rect 135168 259480 135220 259486
rect 135168 259422 135220 259428
rect 133786 258768 133842 258777
rect 133786 258703 133788 258712
rect 133840 258703 133842 258712
rect 133788 258674 133840 258680
rect 133236 255332 133288 255338
rect 133236 255274 133288 255280
rect 133248 230450 133276 255274
rect 133788 250504 133840 250510
rect 133788 250446 133840 250452
rect 133800 249830 133828 250446
rect 133788 249824 133840 249830
rect 133788 249766 133840 249772
rect 133984 238754 134012 259422
rect 135168 251864 135220 251870
rect 135168 251806 135220 251812
rect 135180 251258 135208 251806
rect 134616 251252 134668 251258
rect 134616 251194 134668 251200
rect 135168 251252 135220 251258
rect 135168 251194 135220 251200
rect 133892 238726 134012 238754
rect 133236 230444 133288 230450
rect 133236 230386 133288 230392
rect 133144 115932 133196 115938
rect 133144 115874 133196 115880
rect 133248 110430 133276 230386
rect 133788 115932 133840 115938
rect 133788 115874 133840 115880
rect 133800 115258 133828 115874
rect 133788 115252 133840 115258
rect 133788 115194 133840 115200
rect 133892 113393 133920 238726
rect 134522 215928 134578 215937
rect 134522 215863 134578 215872
rect 133878 113384 133934 113393
rect 133878 113319 133934 113328
rect 133236 110424 133288 110430
rect 133236 110366 133288 110372
rect 132512 16546 133000 16574
rect 129004 7608 129056 7614
rect 129004 7550 129056 7556
rect 126242 3496 126298 3505
rect 126242 3431 126298 3440
rect 129372 2168 129424 2174
rect 129372 2110 129424 2116
rect 129384 480 129412 2110
rect 132972 480 133000 16546
rect 134536 3534 134564 215863
rect 134628 99346 134656 251194
rect 134708 235272 134760 235278
rect 134708 235214 134760 235220
rect 134720 128314 134748 235214
rect 134708 128308 134760 128314
rect 134708 128250 134760 128256
rect 135272 126954 135300 273906
rect 135350 244896 135406 244905
rect 135350 244831 135406 244840
rect 135260 126948 135312 126954
rect 135260 126890 135312 126896
rect 135364 103494 135392 244831
rect 135456 224262 135484 277366
rect 136548 276072 136600 276078
rect 136548 276014 136600 276020
rect 136560 273970 136588 276014
rect 136548 273964 136600 273970
rect 136548 273906 136600 273912
rect 135904 269816 135956 269822
rect 135904 269758 135956 269764
rect 135916 269142 135944 269758
rect 135904 269136 135956 269142
rect 135904 269078 135956 269084
rect 135444 224256 135496 224262
rect 135444 224198 135496 224204
rect 135916 122806 135944 269078
rect 136548 224936 136600 224942
rect 136548 224878 136600 224884
rect 136560 224262 136588 224878
rect 136548 224256 136600 224262
rect 136548 224198 136600 224204
rect 136652 208282 136680 386310
rect 136744 323610 136772 440302
rect 141424 426488 141476 426494
rect 141424 426430 141476 426436
rect 140780 413296 140832 413302
rect 140780 413238 140832 413244
rect 139400 381540 139452 381546
rect 139400 381482 139452 381488
rect 138020 378888 138072 378894
rect 138020 378830 138072 378836
rect 136732 323604 136784 323610
rect 136732 323546 136784 323552
rect 137100 315308 137152 315314
rect 137100 315250 137152 315256
rect 137112 314702 137140 315250
rect 136732 314696 136784 314702
rect 136732 314638 136784 314644
rect 137100 314696 137152 314702
rect 137100 314638 137152 314644
rect 136744 258806 136772 314638
rect 137284 306400 137336 306406
rect 137284 306342 137336 306348
rect 136732 258800 136784 258806
rect 136732 258742 136784 258748
rect 136640 208276 136692 208282
rect 136640 208218 136692 208224
rect 136652 207670 136680 208218
rect 136640 207664 136692 207670
rect 136640 207606 136692 207612
rect 136638 192536 136694 192545
rect 136638 192471 136694 192480
rect 135904 122800 135956 122806
rect 135904 122742 135956 122748
rect 135916 122126 135944 122742
rect 135904 122120 135956 122126
rect 135904 122062 135956 122068
rect 135352 103488 135404 103494
rect 135352 103430 135404 103436
rect 135364 102814 135392 103430
rect 135352 102808 135404 102814
rect 135352 102750 135404 102756
rect 134616 99340 134668 99346
rect 134616 99282 134668 99288
rect 135168 99340 135220 99346
rect 135168 99282 135220 99288
rect 135180 98666 135208 99282
rect 135168 98660 135220 98666
rect 135168 98602 135220 98608
rect 136454 4992 136510 5001
rect 136454 4927 136510 4936
rect 134524 3528 134576 3534
rect 134524 3470 134576 3476
rect 136468 480 136496 4927
rect 136652 2174 136680 192471
rect 136744 111790 136772 258742
rect 136732 111784 136784 111790
rect 136732 111726 136784 111732
rect 137296 89010 137324 306342
rect 138032 220289 138060 378830
rect 138664 233300 138716 233306
rect 138664 233242 138716 233248
rect 138018 220280 138074 220289
rect 138018 220215 138074 220224
rect 138676 202842 138704 233242
rect 139412 213858 139440 381482
rect 139492 298172 139544 298178
rect 139492 298114 139544 298120
rect 139504 213897 139532 298114
rect 140792 235385 140820 413238
rect 141436 345098 141464 426430
rect 142160 424380 142212 424386
rect 142160 424322 142212 424328
rect 141424 345092 141476 345098
rect 141424 345034 141476 345040
rect 141436 323649 141464 345034
rect 141422 323640 141478 323649
rect 141422 323575 141478 323584
rect 141424 300892 141476 300898
rect 141424 300834 141476 300840
rect 141436 274650 141464 300834
rect 142172 275330 142200 424322
rect 144184 422952 144236 422958
rect 144184 422894 144236 422900
rect 143540 414044 143592 414050
rect 143540 413986 143592 413992
rect 142804 402280 142856 402286
rect 142804 402222 142856 402228
rect 142816 339590 142844 402222
rect 142804 339584 142856 339590
rect 142804 339526 142856 339532
rect 142816 301510 142844 339526
rect 142804 301504 142856 301510
rect 142804 301446 142856 301452
rect 142988 278792 143040 278798
rect 142988 278734 143040 278740
rect 142160 275324 142212 275330
rect 142160 275266 142212 275272
rect 142896 275324 142948 275330
rect 142896 275266 142948 275272
rect 141424 274644 141476 274650
rect 141424 274586 141476 274592
rect 141516 267028 141568 267034
rect 141516 266970 141568 266976
rect 140778 235376 140834 235385
rect 140778 235311 140834 235320
rect 141422 225584 141478 225593
rect 141422 225519 141478 225528
rect 139490 213888 139546 213897
rect 139400 213852 139452 213858
rect 139490 213823 139546 213832
rect 139400 213794 139452 213800
rect 139412 213246 139440 213794
rect 139400 213240 139452 213246
rect 139504 213217 139532 213823
rect 139400 213182 139452 213188
rect 139490 213208 139546 213217
rect 139490 213143 139546 213152
rect 138664 202836 138716 202842
rect 138664 202778 138716 202784
rect 137284 89004 137336 89010
rect 137284 88946 137336 88952
rect 141436 3466 141464 225519
rect 141528 61470 141556 266970
rect 142804 256012 142856 256018
rect 142804 255954 142856 255960
rect 142160 244928 142212 244934
rect 142160 244870 142212 244876
rect 142172 191214 142200 244870
rect 142160 191208 142212 191214
rect 142160 191150 142212 191156
rect 141516 61464 141568 61470
rect 141516 61406 141568 61412
rect 142816 17338 142844 255954
rect 142908 241369 142936 275266
rect 143000 251841 143028 278734
rect 142986 251832 143042 251841
rect 142986 251767 143042 251776
rect 143552 248305 143580 413986
rect 144196 311914 144224 422894
rect 151084 421592 151136 421598
rect 151084 421534 151136 421540
rect 147680 408536 147732 408542
rect 147680 408478 147732 408484
rect 146300 405000 146352 405006
rect 146300 404942 146352 404948
rect 144920 403640 144972 403646
rect 144920 403582 144972 403588
rect 144184 311908 144236 311914
rect 144184 311850 144236 311856
rect 144196 276078 144224 311850
rect 144828 276684 144880 276690
rect 144828 276626 144880 276632
rect 144184 276072 144236 276078
rect 144184 276014 144236 276020
rect 143538 248296 143594 248305
rect 143538 248231 143594 248240
rect 143552 247625 143580 248231
rect 143538 247616 143594 247625
rect 143538 247551 143594 247560
rect 143448 244928 143500 244934
rect 143448 244870 143500 244876
rect 143460 244322 143488 244870
rect 143448 244316 143500 244322
rect 143448 244258 143500 244264
rect 142894 241360 142950 241369
rect 142894 241295 142950 241304
rect 142908 235278 142936 241295
rect 142896 235272 142948 235278
rect 142896 235214 142948 235220
rect 142804 17332 142856 17338
rect 142804 17274 142856 17280
rect 144840 3534 144868 276626
rect 144932 260166 144960 403582
rect 144920 260160 144972 260166
rect 144920 260102 144972 260108
rect 146312 233073 146340 404942
rect 147692 264738 147720 408478
rect 149060 407176 149112 407182
rect 149060 407118 149112 407124
rect 147772 392012 147824 392018
rect 147772 391954 147824 391960
rect 147600 264710 147720 264738
rect 147600 263634 147628 264710
rect 147588 263628 147640 263634
rect 147588 263570 147640 263576
rect 147600 262886 147628 263570
rect 147588 262880 147640 262886
rect 147588 262822 147640 262828
rect 146944 257372 146996 257378
rect 146944 257314 146996 257320
rect 146298 233064 146354 233073
rect 146298 232999 146354 233008
rect 146956 73846 146984 257314
rect 147784 250510 147812 391954
rect 148324 285796 148376 285802
rect 148324 285738 148376 285744
rect 148336 263566 148364 285738
rect 149072 266354 149100 407118
rect 151096 341018 151124 421534
rect 151820 400240 151872 400246
rect 151820 400182 151872 400188
rect 151084 341012 151136 341018
rect 151084 340954 151136 340960
rect 151096 324970 151124 340954
rect 151084 324964 151136 324970
rect 151084 324906 151136 324912
rect 151084 318912 151136 318918
rect 151084 318854 151136 318860
rect 151096 304298 151124 318854
rect 151084 304292 151136 304298
rect 151084 304234 151136 304240
rect 151082 302560 151138 302569
rect 151082 302495 151138 302504
rect 151096 278050 151124 302495
rect 151832 293282 151860 400182
rect 191104 394732 191156 394738
rect 191104 394674 191156 394680
rect 187700 393372 187752 393378
rect 187700 393314 187752 393320
rect 180154 313440 180210 313449
rect 180154 313375 180210 313384
rect 160744 311976 160796 311982
rect 160744 311918 160796 311924
rect 152462 307864 152518 307873
rect 152462 307799 152518 307808
rect 151820 293276 151872 293282
rect 151820 293218 151872 293224
rect 151176 284980 151228 284986
rect 151176 284922 151228 284928
rect 151084 278044 151136 278050
rect 151084 277986 151136 277992
rect 149060 266348 149112 266354
rect 149060 266290 149112 266296
rect 149072 265674 149100 266290
rect 149060 265668 149112 265674
rect 149060 265610 149112 265616
rect 148324 263560 148376 263566
rect 148324 263502 148376 263508
rect 148324 255332 148376 255338
rect 148324 255274 148376 255280
rect 147772 250504 147824 250510
rect 147772 250446 147824 250452
rect 147036 200796 147088 200802
rect 147036 200738 147088 200744
rect 146944 73840 146996 73846
rect 146944 73782 146996 73788
rect 147048 32434 147076 200738
rect 147036 32428 147088 32434
rect 147036 32370 147088 32376
rect 148336 15978 148364 255274
rect 151084 254040 151136 254046
rect 151084 253982 151136 253988
rect 151096 80782 151124 253982
rect 151188 184210 151216 284922
rect 151176 184204 151228 184210
rect 151176 184146 151228 184152
rect 151176 100020 151228 100026
rect 151176 99962 151228 99968
rect 151084 80776 151136 80782
rect 151084 80718 151136 80724
rect 151188 21418 151216 99962
rect 151176 21412 151228 21418
rect 151176 21354 151228 21360
rect 148324 15972 148376 15978
rect 148324 15914 148376 15920
rect 143540 3528 143592 3534
rect 143540 3470 143592 3476
rect 144828 3528 144880 3534
rect 144828 3470 144880 3476
rect 141424 3460 141476 3466
rect 141424 3402 141476 3408
rect 136640 2168 136692 2174
rect 136640 2110 136692 2116
rect 143552 480 143580 3470
rect 152476 3369 152504 307799
rect 160756 306338 160784 311918
rect 160836 310616 160888 310622
rect 160836 310558 160888 310564
rect 160744 306332 160796 306338
rect 160744 306274 160796 306280
rect 155408 305040 155460 305046
rect 155408 304982 155460 304988
rect 153108 293956 153160 293962
rect 153108 293898 153160 293904
rect 153120 293282 153148 293898
rect 153108 293276 153160 293282
rect 153108 293218 153160 293224
rect 155224 275324 155276 275330
rect 155224 275266 155276 275272
rect 155236 6254 155264 275266
rect 155316 263628 155368 263634
rect 155316 263570 155368 263576
rect 155328 71058 155356 263570
rect 155420 256018 155448 304982
rect 160848 304978 160876 310558
rect 180064 309868 180116 309874
rect 180064 309810 180116 309816
rect 178774 306640 178830 306649
rect 178774 306575 178830 306584
rect 176016 306468 176068 306474
rect 176016 306410 176068 306416
rect 160836 304972 160888 304978
rect 160836 304914 160888 304920
rect 160744 303680 160796 303686
rect 160744 303622 160796 303628
rect 159364 291916 159416 291922
rect 159364 291858 159416 291864
rect 156602 276720 156658 276729
rect 156602 276655 156658 276664
rect 155408 256012 155460 256018
rect 155408 255954 155460 255960
rect 156616 180130 156644 276655
rect 157982 257272 158038 257281
rect 157982 257207 158038 257216
rect 157996 191146 158024 257207
rect 157984 191140 158036 191146
rect 157984 191082 158036 191088
rect 156604 180124 156656 180130
rect 156604 180066 156656 180072
rect 155316 71052 155368 71058
rect 155316 70994 155368 71000
rect 155224 6248 155276 6254
rect 155224 6190 155276 6196
rect 159376 6186 159404 291858
rect 159456 265668 159508 265674
rect 159456 265610 159508 265616
rect 159468 119406 159496 265610
rect 159456 119400 159508 119406
rect 159456 119342 159508 119348
rect 160756 13122 160784 303622
rect 173164 302252 173216 302258
rect 173164 302194 173216 302200
rect 160836 300960 160888 300966
rect 160836 300902 160888 300908
rect 160848 37942 160876 300902
rect 166354 298888 166410 298897
rect 166354 298823 166410 298832
rect 166262 291816 166318 291825
rect 166262 291751 166318 291760
rect 162124 290488 162176 290494
rect 162124 290430 162176 290436
rect 160928 271924 160980 271930
rect 160928 271866 160980 271872
rect 160940 242865 160968 271866
rect 160926 242856 160982 242865
rect 160926 242791 160982 242800
rect 162136 68406 162164 290430
rect 165528 285796 165580 285802
rect 165528 285738 165580 285744
rect 162216 277432 162268 277438
rect 162216 277374 162268 277380
rect 162228 266354 162256 277374
rect 163596 271924 163648 271930
rect 163596 271866 163648 271872
rect 162216 266348 162268 266354
rect 162216 266290 162268 266296
rect 163504 251932 163556 251938
rect 163504 251874 163556 251880
rect 163516 200802 163544 251874
rect 163608 243574 163636 271866
rect 163596 243568 163648 243574
rect 163596 243510 163648 243516
rect 163504 200796 163556 200802
rect 163504 200738 163556 200744
rect 162124 68400 162176 68406
rect 162124 68342 162176 68348
rect 165540 57254 165568 285738
rect 165528 57248 165580 57254
rect 165528 57190 165580 57196
rect 166276 50454 166304 291751
rect 166368 182850 166396 298823
rect 170404 295384 170456 295390
rect 170404 295326 170456 295332
rect 169024 287700 169076 287706
rect 169024 287642 169076 287648
rect 168288 274712 168340 274718
rect 168288 274654 168340 274660
rect 166356 182844 166408 182850
rect 166356 182786 166408 182792
rect 168300 100026 168328 274654
rect 168288 100020 168340 100026
rect 168288 99962 168340 99968
rect 166264 50448 166316 50454
rect 166264 50390 166316 50396
rect 160836 37936 160888 37942
rect 160836 37878 160888 37884
rect 160744 13116 160796 13122
rect 160744 13058 160796 13064
rect 169036 8974 169064 287642
rect 169116 280220 169168 280226
rect 169116 280162 169168 280168
rect 169128 272542 169156 280162
rect 169116 272536 169168 272542
rect 169116 272478 169168 272484
rect 169128 112470 169156 272478
rect 170416 251870 170444 295326
rect 171784 271992 171836 271998
rect 171784 271934 171836 271940
rect 170496 252612 170548 252618
rect 170496 252554 170548 252560
rect 170404 251864 170456 251870
rect 170404 251806 170456 251812
rect 170404 249824 170456 249830
rect 170404 249766 170456 249772
rect 169116 112464 169168 112470
rect 169116 112406 169168 112412
rect 170416 14482 170444 249766
rect 170508 144226 170536 252554
rect 171796 217326 171824 271934
rect 173176 271182 173204 302194
rect 173256 284368 173308 284374
rect 173256 284310 173308 284316
rect 173164 271176 173216 271182
rect 173164 271118 173216 271124
rect 173164 256760 173216 256766
rect 173164 256702 173216 256708
rect 171784 217320 171836 217326
rect 171784 217262 171836 217268
rect 170496 144220 170548 144226
rect 170496 144162 170548 144168
rect 170496 137284 170548 137290
rect 170496 137226 170548 137232
rect 170508 19990 170536 137226
rect 173176 57322 173204 256702
rect 173268 253230 173296 284310
rect 175188 279472 175240 279478
rect 175188 279414 175240 279420
rect 175200 278798 175228 279414
rect 175188 278792 175240 278798
rect 175188 278734 175240 278740
rect 174544 262880 174596 262886
rect 174544 262822 174596 262828
rect 173348 258732 173400 258738
rect 173348 258674 173400 258680
rect 173256 253224 173308 253230
rect 173256 253166 173308 253172
rect 173360 237289 173388 258674
rect 173346 237280 173402 237289
rect 173346 237215 173402 237224
rect 174556 231810 174584 262822
rect 174544 231804 174596 231810
rect 174544 231746 174596 231752
rect 173256 123480 173308 123486
rect 173256 123422 173308 123428
rect 173164 57316 173216 57322
rect 173164 57258 173216 57264
rect 170496 19984 170548 19990
rect 170496 19926 170548 19932
rect 173268 14482 173296 123422
rect 175200 95946 175228 278734
rect 175924 258120 175976 258126
rect 175924 258062 175976 258068
rect 175188 95940 175240 95946
rect 175188 95882 175240 95888
rect 175936 20058 175964 258062
rect 176028 257378 176056 306410
rect 178682 301608 178738 301617
rect 178682 301543 178738 301552
rect 177396 266416 177448 266422
rect 177396 266358 177448 266364
rect 177304 258188 177356 258194
rect 177304 258130 177356 258136
rect 176016 257372 176068 257378
rect 176016 257314 176068 257320
rect 177316 51746 177344 258130
rect 177408 218754 177436 266358
rect 178696 246362 178724 301543
rect 178788 284986 178816 306575
rect 179418 295352 179474 295361
rect 179418 295287 179474 295296
rect 179432 288386 179460 295287
rect 179420 288380 179472 288386
rect 179420 288322 179472 288328
rect 178776 284980 178828 284986
rect 178776 284922 178828 284928
rect 178776 267776 178828 267782
rect 178776 267718 178828 267724
rect 178684 246356 178736 246362
rect 178684 246298 178736 246304
rect 178682 241632 178738 241641
rect 178682 241567 178738 241576
rect 177396 218748 177448 218754
rect 177396 218690 177448 218696
rect 178696 65550 178724 241567
rect 178788 164898 178816 267718
rect 178776 164892 178828 164898
rect 178776 164834 178828 164840
rect 178776 96008 178828 96014
rect 178776 95950 178828 95956
rect 178684 65544 178736 65550
rect 178684 65486 178736 65492
rect 177304 51740 177356 51746
rect 177304 51682 177356 51688
rect 175924 20052 175976 20058
rect 175924 19994 175976 20000
rect 170404 14476 170456 14482
rect 170404 14418 170456 14424
rect 173256 14476 173308 14482
rect 173256 14418 173308 14424
rect 178788 11762 178816 95950
rect 180076 68338 180104 309810
rect 180168 267034 180196 313375
rect 186964 313336 187016 313342
rect 186964 313278 187016 313284
rect 185674 309360 185730 309369
rect 185674 309295 185730 309304
rect 185582 305144 185638 305153
rect 182824 305108 182876 305114
rect 185582 305079 185638 305088
rect 182824 305050 182876 305056
rect 182836 276690 182864 305050
rect 184204 303748 184256 303754
rect 184204 303690 184256 303696
rect 182824 276684 182876 276690
rect 182824 276626 182876 276632
rect 181444 269136 181496 269142
rect 181444 269078 181496 269084
rect 180156 267028 180208 267034
rect 180156 266970 180208 266976
rect 180248 253972 180300 253978
rect 180248 253914 180300 253920
rect 180156 248464 180208 248470
rect 180156 248406 180208 248412
rect 180168 155242 180196 248406
rect 180260 238678 180288 253914
rect 180340 242208 180392 242214
rect 180340 242150 180392 242156
rect 180248 238672 180300 238678
rect 180248 238614 180300 238620
rect 180352 235958 180380 242150
rect 180340 235952 180392 235958
rect 180340 235894 180392 235900
rect 181456 189786 181484 269078
rect 182824 264988 182876 264994
rect 182824 264930 182876 264936
rect 181534 261080 181590 261089
rect 181534 261015 181590 261024
rect 181548 227730 181576 261015
rect 181536 227724 181588 227730
rect 181536 227666 181588 227672
rect 181444 189780 181496 189786
rect 181444 189722 181496 189728
rect 180156 155236 180208 155242
rect 180156 155178 180208 155184
rect 182836 106962 182864 264930
rect 182916 260160 182968 260166
rect 182916 260102 182968 260108
rect 182928 234598 182956 260102
rect 182916 234592 182968 234598
rect 182916 234534 182968 234540
rect 182824 106956 182876 106962
rect 182824 106898 182876 106904
rect 180156 105596 180208 105602
rect 180156 105538 180208 105544
rect 180064 68332 180116 68338
rect 180064 68274 180116 68280
rect 178776 11756 178828 11762
rect 178776 11698 178828 11704
rect 180168 8974 180196 105538
rect 184216 75206 184244 303690
rect 184296 302320 184348 302326
rect 184296 302262 184348 302268
rect 184308 257281 184336 302262
rect 185596 265674 185624 305079
rect 185688 284889 185716 309295
rect 186318 301472 186374 301481
rect 186318 301407 186374 301416
rect 186332 298926 186360 301407
rect 186320 298920 186372 298926
rect 186320 298862 186372 298868
rect 185674 284880 185730 284889
rect 185674 284815 185730 284824
rect 186976 280158 187004 313278
rect 187054 306776 187110 306785
rect 187054 306711 187110 306720
rect 187068 287706 187096 306711
rect 187056 287700 187108 287706
rect 187056 287642 187108 287648
rect 187148 282192 187200 282198
rect 187148 282134 187200 282140
rect 186964 280152 187016 280158
rect 186964 280094 187016 280100
rect 185584 265668 185636 265674
rect 185584 265610 185636 265616
rect 185584 262268 185636 262274
rect 185584 262210 185636 262216
rect 184294 257272 184350 257281
rect 184294 257207 184350 257216
rect 184386 247072 184442 247081
rect 184386 247007 184442 247016
rect 184296 245676 184348 245682
rect 184296 245618 184348 245624
rect 184308 167686 184336 245618
rect 184400 223514 184428 247007
rect 184388 223508 184440 223514
rect 184388 223450 184440 223456
rect 184296 167680 184348 167686
rect 184296 167622 184348 167628
rect 184296 102808 184348 102814
rect 184296 102750 184348 102756
rect 184204 75200 184256 75206
rect 184204 75142 184256 75148
rect 169024 8968 169076 8974
rect 169024 8910 169076 8916
rect 180156 8968 180208 8974
rect 180156 8910 180208 8916
rect 184308 7614 184336 102750
rect 185596 13190 185624 262210
rect 186964 251252 187016 251258
rect 186964 251194 187016 251200
rect 186976 18630 187004 251194
rect 187056 243024 187108 243030
rect 187056 242966 187108 242972
rect 187068 162178 187096 242966
rect 187160 240009 187188 282134
rect 187712 279478 187740 393314
rect 188342 317520 188398 317529
rect 188342 317455 188398 317464
rect 188356 309874 188384 317455
rect 188526 310856 188582 310865
rect 188526 310791 188582 310800
rect 188344 309868 188396 309874
rect 188344 309810 188396 309816
rect 188342 309496 188398 309505
rect 188342 309431 188398 309440
rect 187700 279472 187752 279478
rect 187700 279414 187752 279420
rect 188356 275330 188384 309431
rect 188540 306377 188568 310791
rect 189724 309188 189776 309194
rect 189724 309130 189776 309136
rect 188526 306368 188582 306377
rect 188526 306303 188582 306312
rect 188434 301336 188490 301345
rect 188434 301271 188490 301280
rect 188344 275324 188396 275330
rect 188344 275266 188396 275272
rect 188448 269822 188476 301271
rect 189736 281518 189764 309130
rect 189814 305008 189870 305017
rect 189814 304943 189870 304952
rect 189828 291922 189856 304943
rect 191116 299985 191144 394674
rect 232504 388476 232556 388482
rect 232504 388418 232556 388424
rect 191196 335368 191248 335374
rect 191196 335310 191248 335316
rect 191208 300937 191236 335310
rect 226984 329928 227036 329934
rect 226984 329870 227036 329876
rect 192484 324420 192536 324426
rect 192484 324362 192536 324368
rect 208676 324420 208728 324426
rect 208676 324362 208728 324368
rect 191378 308000 191434 308009
rect 191378 307935 191434 307944
rect 191286 302424 191342 302433
rect 191286 302359 191342 302368
rect 191194 300928 191250 300937
rect 191194 300863 191250 300872
rect 191102 299976 191158 299985
rect 191102 299911 191158 299920
rect 191116 294642 191144 299911
rect 191196 295996 191248 296002
rect 191196 295938 191248 295944
rect 191104 294636 191156 294642
rect 191104 294578 191156 294584
rect 191208 292233 191236 295938
rect 191194 292224 191250 292233
rect 191194 292159 191250 292168
rect 189816 291916 189868 291922
rect 189816 291858 189868 291864
rect 191104 291848 191156 291854
rect 191104 291790 191156 291796
rect 190828 288380 190880 288386
rect 190828 288322 190880 288328
rect 190840 287473 190868 288322
rect 190826 287464 190882 287473
rect 190826 287399 190882 287408
rect 190368 285728 190420 285734
rect 190368 285670 190420 285676
rect 190380 284345 190408 285670
rect 190366 284336 190422 284345
rect 190366 284271 190422 284280
rect 189724 281512 189776 281518
rect 189724 281454 189776 281460
rect 191116 276865 191144 291790
rect 191300 282849 191328 302359
rect 191392 291825 191420 307935
rect 191746 299024 191802 299033
rect 191746 298959 191802 298968
rect 191760 298926 191788 298959
rect 191748 298920 191800 298926
rect 191748 298862 191800 298868
rect 191470 297528 191526 297537
rect 191470 297463 191526 297472
rect 191484 296857 191512 297463
rect 191470 296848 191526 296857
rect 191470 296783 191526 296792
rect 191746 296168 191802 296177
rect 191746 296103 191802 296112
rect 191760 295390 191788 296103
rect 191748 295384 191800 295390
rect 191748 295326 191800 295332
rect 191654 294264 191710 294273
rect 191654 294199 191710 294208
rect 191668 294030 191696 294199
rect 191656 294024 191708 294030
rect 191656 293966 191708 293972
rect 191748 293956 191800 293962
rect 191748 293898 191800 293904
rect 191760 293185 191788 293898
rect 191746 293176 191802 293185
rect 191746 293111 191802 293120
rect 191472 292596 191524 292602
rect 191472 292538 191524 292544
rect 191378 291816 191434 291825
rect 191378 291751 191434 291760
rect 191286 282840 191342 282849
rect 191286 282775 191342 282784
rect 191484 281625 191512 292538
rect 191654 291272 191710 291281
rect 191654 291207 191710 291216
rect 191668 289105 191696 291207
rect 192496 290494 192524 324362
rect 201590 320240 201646 320249
rect 201590 320175 201646 320184
rect 193770 316296 193826 316305
rect 193770 316231 193826 316240
rect 193784 306374 193812 316231
rect 200302 311944 200358 311953
rect 200302 311879 200358 311888
rect 199658 306504 199714 306513
rect 199658 306439 199714 306448
rect 193508 306346 193812 306374
rect 192574 301744 192630 301753
rect 192574 301679 192630 301688
rect 192484 290488 192536 290494
rect 192484 290430 192536 290436
rect 191746 290320 191802 290329
rect 191746 290255 191802 290264
rect 191760 289882 191788 290255
rect 191748 289876 191800 289882
rect 191748 289818 191800 289824
rect 191746 289368 191802 289377
rect 191746 289303 191802 289312
rect 191654 289096 191710 289105
rect 191654 289031 191710 289040
rect 191760 288454 191788 289303
rect 191748 288448 191800 288454
rect 191748 288390 191800 288396
rect 192588 287065 192616 301679
rect 193508 300830 193536 306346
rect 197268 305108 197320 305114
rect 197268 305050 197320 305056
rect 195518 303920 195574 303929
rect 195518 303855 195574 303864
rect 195532 301580 195560 303855
rect 197280 301580 197308 305050
rect 197910 303648 197966 303657
rect 197910 303583 197966 303592
rect 197542 301744 197598 301753
rect 197542 301679 197598 301688
rect 197556 301481 197584 301679
rect 197924 301580 197952 303583
rect 199672 301580 199700 306439
rect 200316 303618 200344 311879
rect 200394 310720 200450 310729
rect 200394 310655 200450 310664
rect 200304 303612 200356 303618
rect 200304 303554 200356 303560
rect 200212 302320 200264 302326
rect 200212 302262 200264 302268
rect 200224 301580 200252 302262
rect 200408 301594 200436 310655
rect 201132 303612 201184 303618
rect 201132 303554 201184 303560
rect 201144 301594 201172 303554
rect 201604 301594 201632 320175
rect 203246 313304 203302 313313
rect 203246 313239 203302 313248
rect 203260 301594 203288 313239
rect 207754 308000 207810 308009
rect 207754 307935 207810 307944
rect 204258 306640 204314 306649
rect 204258 306575 204314 306584
rect 200408 301566 200790 301594
rect 201144 301566 201434 301594
rect 201604 301566 201986 301594
rect 203260 301566 203734 301594
rect 204272 301580 204300 306575
rect 206006 305144 206062 305153
rect 206006 305079 206062 305088
rect 205456 303748 205508 303754
rect 205456 303690 205508 303696
rect 205468 301580 205496 303690
rect 206020 301580 206048 305079
rect 207768 301580 207796 307935
rect 208398 306776 208454 306785
rect 208398 306711 208454 306720
rect 208412 301580 208440 306711
rect 208688 301594 208716 324362
rect 222198 316160 222254 316169
rect 222198 316095 222254 316104
rect 214562 314936 214618 314945
rect 214562 314871 214618 314880
rect 213182 313440 213238 313449
rect 213182 313375 213238 313384
rect 209778 309496 209834 309505
rect 209778 309431 209834 309440
rect 209792 301594 209820 309431
rect 211894 305008 211950 305017
rect 211894 304943 211950 304952
rect 211252 303748 211304 303754
rect 211252 303690 211304 303696
rect 208688 301566 208978 301594
rect 209792 301566 210174 301594
rect 211264 301580 211292 303690
rect 211908 301580 211936 304943
rect 213196 301594 213224 313375
rect 214576 305658 214604 314871
rect 218518 314800 218574 314809
rect 218518 314735 218574 314744
rect 218244 307896 218296 307902
rect 218244 307838 218296 307844
rect 215944 306468 215996 306474
rect 215944 306410 215996 306416
rect 214564 305652 214616 305658
rect 214564 305594 214616 305600
rect 214196 305040 214248 305046
rect 214196 304982 214248 304988
rect 213196 301566 213670 301594
rect 214208 301580 214236 304982
rect 215956 301580 215984 306410
rect 218256 301580 218284 307838
rect 218532 301594 218560 314735
rect 219622 310584 219678 310593
rect 219622 310519 219678 310528
rect 219636 301594 219664 310519
rect 220818 309224 220874 309233
rect 220818 309159 220874 309168
rect 220832 301594 220860 309159
rect 222212 301594 222240 316095
rect 226996 315353 227024 329870
rect 227718 317520 227774 317529
rect 227718 317455 227774 317464
rect 226982 315344 227038 315353
rect 226982 315279 227038 315288
rect 226982 305008 227038 305017
rect 226982 304943 227038 304952
rect 218532 301566 218914 301594
rect 219636 301566 220018 301594
rect 220832 301566 221214 301594
rect 222212 301566 222410 301594
rect 226996 301580 227024 304943
rect 227732 301594 227760 317455
rect 232516 305182 232544 388418
rect 260104 349172 260156 349178
rect 260104 349114 260156 349120
rect 240140 343664 240192 343670
rect 240140 343606 240192 343612
rect 238024 336048 238076 336054
rect 238024 335990 238076 335996
rect 233884 334076 233936 334082
rect 233884 334018 233936 334024
rect 233896 308446 233924 334018
rect 233884 308440 233936 308446
rect 233884 308382 233936 308388
rect 234618 307864 234674 307873
rect 234618 307799 234674 307808
rect 232504 305176 232556 305182
rect 232504 305118 232556 305124
rect 229374 303784 229430 303793
rect 229374 303719 229430 303728
rect 227732 301566 228206 301594
rect 229388 301580 229416 303719
rect 230478 303648 230534 303657
rect 230478 303583 230534 303592
rect 230492 301580 230520 303583
rect 234632 301580 234660 307799
rect 236368 306400 236420 306406
rect 236368 306342 236420 306348
rect 236380 301580 236408 306342
rect 238036 302297 238064 335990
rect 239864 305176 239916 305182
rect 239864 305118 239916 305124
rect 238666 303920 238722 303929
rect 238666 303855 238722 303864
rect 238022 302288 238078 302297
rect 238022 302223 238078 302232
rect 238036 301594 238064 302223
rect 238036 301566 238142 301594
rect 238680 301580 238708 303855
rect 194230 301472 194286 301481
rect 197542 301472 197598 301481
rect 194286 301430 194442 301458
rect 194230 301407 194286 301416
rect 197542 301407 197598 301416
rect 194506 301200 194562 301209
rect 212814 301200 212870 301209
rect 194562 301158 194994 301186
rect 194506 301135 194562 301144
rect 224958 301200 225014 301209
rect 212870 301158 213026 301186
rect 212814 301135 212870 301144
rect 225014 301158 225262 301186
rect 224958 301135 225014 301144
rect 210422 301064 210478 301073
rect 216310 301064 216366 301073
rect 210478 301022 210726 301050
rect 210422 300999 210478 301008
rect 220358 301064 220414 301073
rect 216366 301022 216522 301050
rect 216310 300999 216366 301008
rect 222750 301064 222806 301073
rect 220414 301022 220662 301050
rect 220358 300999 220414 301008
rect 224406 301064 224462 301073
rect 222806 301022 222962 301050
rect 222750 300999 222806 301008
rect 231398 301064 231454 301073
rect 224462 301022 224710 301050
rect 224406 300999 224462 301008
rect 232594 301064 232650 301073
rect 231454 301022 231702 301050
rect 231398 300999 231454 301008
rect 233790 301064 233846 301073
rect 232650 301022 232898 301050
rect 232594 300999 232650 301008
rect 235446 301064 235502 301073
rect 233846 301022 234002 301050
rect 233790 300999 233846 301008
rect 235502 301022 235750 301050
rect 235446 300999 235502 301008
rect 196348 300960 196400 300966
rect 196070 300928 196126 300937
rect 193600 300886 193890 300914
rect 193496 300824 193548 300830
rect 193496 300766 193548 300772
rect 193600 299538 193628 300886
rect 196126 300886 196190 300914
rect 198186 300928 198242 300937
rect 196400 300908 196742 300914
rect 196348 300902 196742 300908
rect 196360 300886 196742 300902
rect 196070 300863 196126 300872
rect 198830 300928 198886 300937
rect 198242 300886 198490 300914
rect 198186 300863 198242 300872
rect 202326 300928 202382 300937
rect 198886 300886 199042 300914
rect 198830 300863 198886 300872
rect 203062 300928 203118 300937
rect 202382 300886 202538 300914
rect 202326 300863 202382 300872
rect 204626 300928 204682 300937
rect 203118 300886 203182 300914
rect 203062 300863 203118 300872
rect 206282 300928 206338 300937
rect 204682 300886 204930 300914
rect 204626 300863 204682 300872
rect 207110 300928 207166 300937
rect 206338 300886 206678 300914
rect 206282 300863 206338 300872
rect 209318 300928 209374 300937
rect 207166 300886 207230 300914
rect 207110 300863 207166 300872
rect 212170 300928 212226 300937
rect 209374 300886 209530 300914
rect 209318 300863 209374 300872
rect 214286 300928 214342 300937
rect 212226 300886 212474 300914
rect 212170 300863 212226 300872
rect 215114 300928 215170 300937
rect 214342 300886 214774 300914
rect 214286 300863 214342 300872
rect 216678 300928 216734 300937
rect 215170 300886 215418 300914
rect 215114 300863 215170 300872
rect 217322 300928 217378 300937
rect 216734 300886 217166 300914
rect 216678 300863 216734 300872
rect 219530 300928 219586 300937
rect 217378 300886 217718 300914
rect 219466 300886 219530 300914
rect 217322 300863 217378 300872
rect 219530 300863 219586 300872
rect 221462 300928 221518 300937
rect 223210 300928 223266 300937
rect 221518 300886 221766 300914
rect 221462 300863 221518 300872
rect 224038 300928 224094 300937
rect 223266 300886 223514 300914
rect 223210 300863 223266 300872
rect 225602 300928 225658 300937
rect 224094 300886 224158 300914
rect 224038 300863 224094 300872
rect 226338 300928 226394 300937
rect 225658 300886 225906 300914
rect 225602 300863 225658 300872
rect 227258 300928 227314 300937
rect 226394 300886 226458 300914
rect 226338 300863 226394 300872
rect 228454 300928 228510 300937
rect 227314 300886 227654 300914
rect 227258 300863 227314 300872
rect 229742 300928 229798 300937
rect 228510 300886 228758 300914
rect 228454 300863 228510 300872
rect 231030 300928 231086 300937
rect 229798 300886 229954 300914
rect 229742 300863 229798 300872
rect 232318 300928 232374 300937
rect 231086 300886 231150 300914
rect 232254 300886 232318 300914
rect 231030 300863 231086 300872
rect 232318 300863 232374 300872
rect 233330 300928 233386 300937
rect 234894 300928 234950 300937
rect 233386 300886 233450 300914
rect 233330 300863 233386 300872
rect 236734 300928 236790 300937
rect 234950 300886 235198 300914
rect 234894 300863 234950 300872
rect 237838 300928 237894 300937
rect 236790 300886 236946 300914
rect 237498 300886 237838 300914
rect 236734 300863 236790 300872
rect 237838 300863 237894 300872
rect 238850 300928 238906 300937
rect 239876 300914 239904 305118
rect 240152 302190 240180 343606
rect 253296 340944 253348 340950
rect 253296 340886 253348 340892
rect 240416 339584 240468 339590
rect 240416 339526 240468 339532
rect 240140 302184 240192 302190
rect 240140 302126 240192 302132
rect 240428 301050 240456 339526
rect 251180 338768 251232 338774
rect 248418 338736 248474 338745
rect 251180 338710 251232 338716
rect 248418 338671 248474 338680
rect 242164 338156 242216 338162
rect 242164 338098 242216 338104
rect 240784 334008 240836 334014
rect 240784 333950 240836 333956
rect 240796 307766 240824 333950
rect 241520 331356 241572 331362
rect 241520 331298 241572 331304
rect 240784 307760 240836 307766
rect 240784 307702 240836 307708
rect 240968 302184 241020 302190
rect 240968 302126 241020 302132
rect 240980 301186 241008 302126
rect 241532 301594 241560 331298
rect 242176 305017 242204 338098
rect 246396 336864 246448 336870
rect 246396 336806 246448 336812
rect 246302 335472 246358 335481
rect 246302 335407 246358 335416
rect 244922 334112 244978 334121
rect 244922 334047 244978 334056
rect 242900 328500 242952 328506
rect 242900 328442 242952 328448
rect 242912 325694 242940 328442
rect 242912 325666 243032 325694
rect 242162 305008 242218 305017
rect 242162 304943 242218 304952
rect 241532 301566 241638 301594
rect 242176 301580 242204 304943
rect 242808 302932 242860 302938
rect 242808 302874 242860 302880
rect 242820 301594 242848 302874
rect 242742 301566 242848 301594
rect 243004 301594 243032 325666
rect 244936 308961 244964 334047
rect 245014 326360 245070 326369
rect 245014 326295 245070 326304
rect 244922 308952 244978 308961
rect 244922 308887 244978 308896
rect 245028 308446 245056 326295
rect 246210 308952 246266 308961
rect 246210 308887 246266 308896
rect 243912 308440 243964 308446
rect 243912 308382 243964 308388
rect 245016 308440 245068 308446
rect 245016 308382 245068 308388
rect 243004 301566 243386 301594
rect 243924 301580 243952 308382
rect 246224 307873 246252 308887
rect 246210 307864 246266 307873
rect 246210 307799 246266 307808
rect 244464 307760 244516 307766
rect 244464 307702 244516 307708
rect 244476 301580 244504 307702
rect 245658 306504 245714 306513
rect 245658 306439 245714 306448
rect 245108 303748 245160 303754
rect 245108 303690 245160 303696
rect 244830 301472 244886 301481
rect 245120 301458 245148 303690
rect 245672 301580 245700 306439
rect 246224 301580 246252 307799
rect 246316 304502 246344 335407
rect 246408 306406 246436 336806
rect 247684 332648 247736 332654
rect 247684 332590 247736 332596
rect 246488 327208 246540 327214
rect 246488 327150 246540 327156
rect 246396 306400 246448 306406
rect 246396 306342 246448 306348
rect 246304 304496 246356 304502
rect 246304 304438 246356 304444
rect 246500 301481 246528 327150
rect 247696 304201 247724 332590
rect 248432 307057 248460 338671
rect 249800 336796 249852 336802
rect 249800 336738 249852 336744
rect 249064 322992 249116 322998
rect 249064 322934 249116 322940
rect 248418 307048 248474 307057
rect 248418 306983 248474 306992
rect 248432 306490 248460 306983
rect 248340 306462 248460 306490
rect 247682 304192 247738 304201
rect 247682 304127 247738 304136
rect 248340 303686 248368 306462
rect 249076 306066 249104 322934
rect 249064 306060 249116 306066
rect 249064 306002 249116 306008
rect 249708 304496 249760 304502
rect 249708 304438 249760 304444
rect 247408 303680 247460 303686
rect 247408 303622 247460 303628
rect 248328 303680 248380 303686
rect 249720 303657 249748 304438
rect 248328 303622 248380 303628
rect 249706 303648 249762 303657
rect 246854 302560 246910 302569
rect 246854 302495 246910 302504
rect 246868 302297 246896 302495
rect 246854 302288 246910 302297
rect 246854 302223 246910 302232
rect 246868 301580 246896 302223
rect 247420 301580 247448 303622
rect 249706 303583 249762 303592
rect 248878 302832 248934 302841
rect 248878 302767 248934 302776
rect 247774 301608 247830 301617
rect 248892 301594 248920 302767
rect 249156 302252 249208 302258
rect 249156 302194 249208 302200
rect 247830 301580 247986 301594
rect 247830 301566 248000 301580
rect 248630 301566 248920 301594
rect 249168 301580 249196 302194
rect 249720 301580 249748 303583
rect 249812 302841 249840 336738
rect 250444 318912 250496 318918
rect 250444 318854 250496 318860
rect 250456 307766 250484 318854
rect 250536 318096 250588 318102
rect 250536 318038 250588 318044
rect 250444 307760 250496 307766
rect 250444 307702 250496 307708
rect 250548 307698 250576 318038
rect 250536 307692 250588 307698
rect 250536 307634 250588 307640
rect 250352 306400 250404 306406
rect 250352 306342 250404 306348
rect 249798 302832 249854 302841
rect 249798 302767 249854 302776
rect 250364 301753 250392 306342
rect 250902 303784 250958 303793
rect 250902 303719 250958 303728
rect 250350 301744 250406 301753
rect 250350 301679 250406 301688
rect 250364 301580 250392 301679
rect 250916 301594 250944 303719
rect 250640 301580 250944 301594
rect 251192 301594 251220 338710
rect 251824 318844 251876 318850
rect 251824 318786 251876 318792
rect 251836 302258 251864 318786
rect 252744 314764 252796 314770
rect 252744 314706 252796 314712
rect 252652 303680 252704 303686
rect 252652 303622 252704 303628
rect 252664 302433 252692 303622
rect 252650 302424 252706 302433
rect 252650 302359 252706 302368
rect 251824 302252 251876 302258
rect 251824 302194 251876 302200
rect 250640 301566 250930 301580
rect 251192 301566 251482 301594
rect 252664 301580 252692 302359
rect 247774 301543 247830 301552
rect 244886 301444 245148 301458
rect 246486 301472 246542 301481
rect 244886 301430 245134 301444
rect 244830 301407 244886 301416
rect 246486 301407 246542 301416
rect 240980 301172 241376 301186
rect 240994 301170 241376 301172
rect 240994 301164 241388 301170
rect 240994 301158 241336 301164
rect 241336 301106 241388 301112
rect 240784 301096 240836 301102
rect 240428 301044 240784 301050
rect 240428 301038 240836 301044
rect 247972 301050 248000 301566
rect 240428 301036 240824 301038
rect 247972 301036 248092 301050
rect 240442 301022 240824 301036
rect 247986 301022 248092 301036
rect 250640 301034 250668 301566
rect 251822 301336 251878 301345
rect 251878 301294 252126 301322
rect 251822 301271 251878 301280
rect 248064 300966 248092 301022
rect 250628 301028 250680 301034
rect 250628 300970 250680 300976
rect 248052 300960 248104 300966
rect 240046 300928 240102 300937
rect 238906 300886 239246 300914
rect 239876 300900 240046 300914
rect 239890 300886 240046 300900
rect 238850 300863 238906 300872
rect 248052 300902 248104 300908
rect 240046 300863 240102 300872
rect 193678 300248 193734 300257
rect 193678 300183 193734 300192
rect 193692 300150 193720 300183
rect 193680 300144 193732 300150
rect 193680 300086 193732 300092
rect 193588 299532 193640 299538
rect 193588 299474 193640 299480
rect 192574 287056 192630 287065
rect 192574 286991 192630 287000
rect 191746 286512 191802 286521
rect 191746 286447 191802 286456
rect 191760 285802 191788 286447
rect 191748 285796 191800 285802
rect 191748 285738 191800 285744
rect 191654 285560 191710 285569
rect 191654 285495 191710 285504
rect 191668 284345 191696 285495
rect 191746 284472 191802 284481
rect 191746 284407 191802 284416
rect 191760 284374 191788 284407
rect 191748 284368 191800 284374
rect 191654 284336 191710 284345
rect 191748 284310 191800 284316
rect 191654 284271 191710 284280
rect 191746 283520 191802 283529
rect 191746 283455 191802 283464
rect 191760 282946 191788 283455
rect 191748 282940 191800 282946
rect 191748 282882 191800 282888
rect 192482 282568 192538 282577
rect 192482 282503 192538 282512
rect 191470 281616 191526 281625
rect 191470 281551 191526 281560
rect 191562 280664 191618 280673
rect 191562 280599 191618 280608
rect 191576 280226 191604 280599
rect 191564 280220 191616 280226
rect 191564 280162 191616 280168
rect 191746 279712 191802 279721
rect 191746 279647 191802 279656
rect 191760 279546 191788 279647
rect 191748 279540 191800 279546
rect 191748 279482 191800 279488
rect 191654 278760 191710 278769
rect 191654 278695 191710 278704
rect 191748 278724 191800 278730
rect 191668 277438 191696 278695
rect 191748 278666 191800 278672
rect 191760 277817 191788 278666
rect 191746 277808 191802 277817
rect 191746 277743 191802 277752
rect 191656 277432 191708 277438
rect 191656 277374 191708 277380
rect 191102 276856 191158 276865
rect 191102 276791 191158 276800
rect 191654 275768 191710 275777
rect 191654 275703 191710 275712
rect 191668 274786 191696 275703
rect 191746 274816 191802 274825
rect 188988 274780 189040 274786
rect 188988 274722 189040 274728
rect 191656 274780 191708 274786
rect 191746 274751 191802 274760
rect 191656 274722 191708 274728
rect 188436 269816 188488 269822
rect 188436 269758 188488 269764
rect 188526 267880 188582 267889
rect 188526 267815 188582 267824
rect 188252 259480 188304 259486
rect 188252 259422 188304 259428
rect 188264 251938 188292 259422
rect 188344 252680 188396 252686
rect 188344 252622 188396 252628
rect 188252 251932 188304 251938
rect 188252 251874 188304 251880
rect 187240 249076 187292 249082
rect 187240 249018 187292 249024
rect 187146 240000 187202 240009
rect 187146 239935 187202 239944
rect 187252 237318 187280 249018
rect 187240 237312 187292 237318
rect 187240 237254 187292 237260
rect 187056 162172 187108 162178
rect 187056 162114 187108 162120
rect 187056 115252 187108 115258
rect 187056 115194 187108 115200
rect 186964 18624 187016 18630
rect 186964 18566 187016 18572
rect 185584 13184 185636 13190
rect 185584 13126 185636 13132
rect 184296 7608 184348 7614
rect 184296 7550 184348 7556
rect 159364 6180 159416 6186
rect 159364 6122 159416 6128
rect 187068 4826 187096 115194
rect 188356 86329 188384 252622
rect 188436 247104 188488 247110
rect 188436 247046 188488 247052
rect 188448 158030 188476 247046
rect 188540 236745 188568 267815
rect 188526 236736 188582 236745
rect 188526 236671 188582 236680
rect 189000 213217 189028 274722
rect 191760 274718 191788 274751
rect 191748 274712 191800 274718
rect 191748 274654 191800 274660
rect 191746 272912 191802 272921
rect 191746 272847 191802 272856
rect 191196 271992 191248 271998
rect 191194 271960 191196 271969
rect 191248 271960 191250 271969
rect 191760 271930 191788 272847
rect 191194 271895 191250 271904
rect 191748 271924 191800 271930
rect 191748 271866 191800 271872
rect 191102 271008 191158 271017
rect 191102 270943 191158 270952
rect 191010 264208 191066 264217
rect 191010 264143 191066 264152
rect 191024 263634 191052 264143
rect 191012 263628 191064 263634
rect 191012 263570 191064 263576
rect 191010 262304 191066 262313
rect 191010 262239 191012 262248
rect 191064 262239 191066 262248
rect 191012 262210 191064 262216
rect 190642 258360 190698 258369
rect 190642 258295 190698 258304
rect 190656 258194 190684 258295
rect 190644 258188 190696 258194
rect 190644 258130 190696 258136
rect 190552 258120 190604 258126
rect 190472 258068 190552 258074
rect 190472 258062 190604 258068
rect 190472 258058 190592 258062
rect 190460 258052 190592 258058
rect 190512 258046 190592 258052
rect 190460 257994 190512 258000
rect 189722 255776 189778 255785
rect 189722 255711 189778 255720
rect 188986 213208 189042 213217
rect 188986 213143 189042 213152
rect 188436 158024 188488 158030
rect 188436 157966 188488 157972
rect 188436 87644 188488 87650
rect 188436 87586 188488 87592
rect 188342 86320 188398 86329
rect 188342 86255 188398 86264
rect 187056 4820 187108 4826
rect 187056 4762 187108 4768
rect 188448 3466 188476 87586
rect 189736 64190 189764 255711
rect 191010 253600 191066 253609
rect 191010 253535 191066 253544
rect 191024 252686 191052 253535
rect 191012 252680 191064 252686
rect 191012 252622 191064 252628
rect 190642 249656 190698 249665
rect 190642 249591 190698 249600
rect 189814 248568 189870 248577
rect 189814 248503 189870 248512
rect 189828 231130 189856 248503
rect 190656 248470 190684 249591
rect 190644 248464 190696 248470
rect 190644 248406 190696 248412
rect 189906 245712 189962 245721
rect 189906 245647 189962 245656
rect 189920 232529 189948 245647
rect 191116 233918 191144 270943
rect 191746 270056 191802 270065
rect 191746 269991 191802 270000
rect 191760 269142 191788 269991
rect 191748 269136 191800 269142
rect 191654 269104 191710 269113
rect 191748 269078 191800 269084
rect 192496 269074 192524 282503
rect 252756 281330 252784 314706
rect 252836 309188 252888 309194
rect 252836 309130 252888 309136
rect 252848 286385 252876 309130
rect 253202 304192 253258 304201
rect 253202 304127 253258 304136
rect 252928 302252 252980 302258
rect 252928 302194 252980 302200
rect 252834 286376 252890 286385
rect 252834 286311 252890 286320
rect 252940 284209 252968 302194
rect 253216 301580 253244 304127
rect 253308 301617 253336 340886
rect 258262 332616 258318 332625
rect 258262 332551 258318 332560
rect 256790 328536 256846 328545
rect 256790 328471 256846 328480
rect 254032 325780 254084 325786
rect 254032 325722 254084 325728
rect 253938 312488 253994 312497
rect 253938 312423 253994 312432
rect 253294 301608 253350 301617
rect 253294 301543 253350 301552
rect 253478 301472 253534 301481
rect 253478 301407 253534 301416
rect 253202 300520 253258 300529
rect 253202 300455 253258 300464
rect 253216 299742 253244 300455
rect 253204 299736 253256 299742
rect 253204 299678 253256 299684
rect 253492 298761 253520 301407
rect 253478 298752 253534 298761
rect 253478 298687 253534 298696
rect 252926 284200 252982 284209
rect 252926 284135 252982 284144
rect 252834 281344 252890 281353
rect 252756 281302 252834 281330
rect 252834 281279 252890 281288
rect 193218 276856 193274 276865
rect 193218 276791 193274 276800
rect 193128 274644 193180 274650
rect 193128 274586 193180 274592
rect 193140 273873 193168 274586
rect 193126 273864 193182 273873
rect 193126 273799 193182 273808
rect 191654 269039 191710 269048
rect 192484 269068 192536 269074
rect 191668 267782 191696 269039
rect 192484 269010 192536 269016
rect 191656 267776 191708 267782
rect 191656 267718 191708 267724
rect 191470 267064 191526 267073
rect 191470 266999 191526 267008
rect 191484 266422 191512 266999
rect 191472 266416 191524 266422
rect 191472 266358 191524 266364
rect 191746 266112 191802 266121
rect 191746 266047 191802 266056
rect 191286 265160 191342 265169
rect 191286 265095 191342 265104
rect 191194 263256 191250 263265
rect 191194 263191 191250 263200
rect 191104 233912 191156 233918
rect 191104 233854 191156 233860
rect 189906 232520 189962 232529
rect 189906 232455 189962 232464
rect 189816 231124 189868 231130
rect 189816 231066 189868 231072
rect 191208 227050 191236 263191
rect 191300 238066 191328 265095
rect 191760 264994 191788 266047
rect 191748 264988 191800 264994
rect 191748 264930 191800 264936
rect 191378 261352 191434 261361
rect 191378 261287 191434 261296
rect 191288 238060 191340 238066
rect 191288 238002 191340 238008
rect 191392 236609 191420 261287
rect 191746 260400 191802 260409
rect 191746 260335 191802 260344
rect 191760 259486 191788 260335
rect 191748 259480 191800 259486
rect 191748 259422 191800 259428
rect 191746 257408 191802 257417
rect 191746 257343 191802 257352
rect 191760 256766 191788 257343
rect 191748 256760 191800 256766
rect 191748 256702 191800 256708
rect 191746 255504 191802 255513
rect 191746 255439 191802 255448
rect 191760 255338 191788 255439
rect 191748 255332 191800 255338
rect 191748 255274 191800 255280
rect 191562 254552 191618 254561
rect 191562 254487 191618 254496
rect 191576 254046 191604 254487
rect 191564 254040 191616 254046
rect 191564 253982 191616 253988
rect 191746 252648 191802 252657
rect 191746 252583 191748 252592
rect 191800 252583 191802 252592
rect 191748 252554 191800 252560
rect 191562 251696 191618 251705
rect 191562 251631 191618 251640
rect 191576 251258 191604 251631
rect 191564 251252 191616 251258
rect 191564 251194 191616 251200
rect 191746 250744 191802 250753
rect 191746 250679 191802 250688
rect 191760 249830 191788 250679
rect 191748 249824 191800 249830
rect 191748 249766 191800 249772
rect 191746 247752 191802 247761
rect 191746 247687 191802 247696
rect 191760 247110 191788 247687
rect 191748 247104 191800 247110
rect 191748 247046 191800 247052
rect 191562 245848 191618 245857
rect 191562 245783 191618 245792
rect 191576 245682 191604 245783
rect 191564 245676 191616 245682
rect 191564 245618 191616 245624
rect 191746 243944 191802 243953
rect 191746 243879 191802 243888
rect 191760 243030 191788 243879
rect 191748 243024 191800 243030
rect 191748 242966 191800 242972
rect 191838 239864 191894 239873
rect 191838 239799 191894 239808
rect 191378 236600 191434 236609
rect 191378 236535 191434 236544
rect 191852 229770 191880 239799
rect 192496 236609 192524 269010
rect 192576 250504 192628 250510
rect 192576 250446 192628 250452
rect 192588 238746 192616 250446
rect 193036 244316 193088 244322
rect 193036 244258 193088 244264
rect 193048 241398 193076 244258
rect 193036 241392 193088 241398
rect 193036 241334 193088 241340
rect 192576 238740 192628 238746
rect 192576 238682 192628 238688
rect 192482 236600 192538 236609
rect 192482 236535 192538 236544
rect 191840 229764 191892 229770
rect 191840 229706 191892 229712
rect 191196 227044 191248 227050
rect 191196 226986 191248 226992
rect 189724 64184 189776 64190
rect 189724 64126 189776 64132
rect 193140 51746 193168 273799
rect 193232 229770 193260 276791
rect 253952 273329 253980 312423
rect 254044 292505 254072 325722
rect 255412 325712 255464 325718
rect 255412 325654 255464 325660
rect 255320 311976 255372 311982
rect 255320 311918 255372 311924
rect 254124 307760 254176 307766
rect 254124 307702 254176 307708
rect 254030 292496 254086 292505
rect 254030 292431 254086 292440
rect 254136 284345 254164 307702
rect 254216 306060 254268 306066
rect 254216 306002 254268 306008
rect 254228 289377 254256 306002
rect 254214 289368 254270 289377
rect 254214 289303 254270 289312
rect 254122 284336 254178 284345
rect 254122 284271 254178 284280
rect 255332 280242 255360 311918
rect 255424 295866 255452 325654
rect 255504 317484 255556 317490
rect 255504 317426 255556 317432
rect 255412 295860 255464 295866
rect 255412 295802 255464 295808
rect 255410 295760 255466 295769
rect 255410 295695 255466 295704
rect 255424 295390 255452 295695
rect 255412 295384 255464 295390
rect 255412 295326 255464 295332
rect 255410 294808 255466 294817
rect 255410 294743 255466 294752
rect 255424 294030 255452 294743
rect 255412 294024 255464 294030
rect 255412 293966 255464 293972
rect 255412 293888 255464 293894
rect 255412 293830 255464 293836
rect 255424 293457 255452 293830
rect 255410 293448 255466 293457
rect 255410 293383 255466 293392
rect 255412 292120 255464 292126
rect 255410 292088 255412 292097
rect 255464 292088 255466 292097
rect 255410 292023 255466 292032
rect 255412 290896 255464 290902
rect 255412 290838 255464 290844
rect 255424 290737 255452 290838
rect 255410 290728 255466 290737
rect 255410 290663 255466 290672
rect 255410 289776 255466 289785
rect 255410 289711 255412 289720
rect 255464 289711 255466 289720
rect 255412 289682 255464 289688
rect 255410 288416 255466 288425
rect 255410 288351 255412 288360
rect 255464 288351 255466 288360
rect 255412 288322 255464 288328
rect 255516 288266 255544 317426
rect 256700 316736 256752 316742
rect 256700 316678 256752 316684
rect 255596 307692 255648 307698
rect 255596 307634 255648 307640
rect 255424 288238 255544 288266
rect 255424 285161 255452 288238
rect 255608 287065 255636 307634
rect 255686 300792 255742 300801
rect 255686 300727 255742 300736
rect 255700 299606 255728 300727
rect 255870 300248 255926 300257
rect 255870 300183 255926 300192
rect 255688 299600 255740 299606
rect 255688 299542 255740 299548
rect 255884 299538 255912 300183
rect 255872 299532 255924 299538
rect 255872 299474 255924 299480
rect 255780 299464 255832 299470
rect 255686 299432 255742 299441
rect 255780 299406 255832 299412
rect 255686 299367 255688 299376
rect 255740 299367 255742 299376
rect 255688 299338 255740 299344
rect 255792 298897 255820 299406
rect 255778 298888 255834 298897
rect 255778 298823 255834 298832
rect 255780 298104 255832 298110
rect 255686 298072 255742 298081
rect 255780 298046 255832 298052
rect 255686 298007 255742 298016
rect 255700 297430 255728 298007
rect 255688 297424 255740 297430
rect 255688 297366 255740 297372
rect 255792 297129 255820 298046
rect 255778 297120 255834 297129
rect 255778 297055 255834 297064
rect 255688 296676 255740 296682
rect 255688 296618 255740 296624
rect 255700 296585 255728 296618
rect 255686 296576 255742 296585
rect 255686 296511 255742 296520
rect 255780 295860 255832 295866
rect 255780 295802 255832 295808
rect 255688 293956 255740 293962
rect 255688 293898 255740 293904
rect 255700 293049 255728 293898
rect 255686 293040 255742 293049
rect 255686 292975 255742 292984
rect 255792 291553 255820 295802
rect 255778 291544 255834 291553
rect 255778 291479 255834 291488
rect 255688 291168 255740 291174
rect 255688 291110 255740 291116
rect 255700 290193 255728 291110
rect 255686 290184 255742 290193
rect 255686 290119 255742 290128
rect 255688 289808 255740 289814
rect 255688 289750 255740 289756
rect 255700 288833 255728 289750
rect 255686 288824 255742 288833
rect 255686 288759 255742 288768
rect 255688 288312 255740 288318
rect 255688 288254 255740 288260
rect 255700 287473 255728 288254
rect 255686 287464 255742 287473
rect 255686 287399 255742 287408
rect 255594 287056 255650 287065
rect 255504 287020 255556 287026
rect 255594 286991 255650 287000
rect 255504 286962 255556 286968
rect 255516 286521 255544 286962
rect 255502 286512 255558 286521
rect 255502 286447 255558 286456
rect 255410 285152 255466 285161
rect 255410 285087 255466 285096
rect 255596 284980 255648 284986
rect 255596 284922 255648 284928
rect 255410 284744 255466 284753
rect 255410 284679 255466 284688
rect 255424 284578 255452 284679
rect 255412 284572 255464 284578
rect 255412 284514 255464 284520
rect 255412 284300 255464 284306
rect 255412 284242 255464 284248
rect 255424 283393 255452 284242
rect 255410 283384 255466 283393
rect 255410 283319 255466 283328
rect 255504 282872 255556 282878
rect 255410 282840 255466 282849
rect 255504 282814 255556 282820
rect 255410 282775 255412 282784
rect 255464 282775 255466 282784
rect 255412 282746 255464 282752
rect 255516 282033 255544 282814
rect 255502 282024 255558 282033
rect 255502 281959 255558 281968
rect 255412 281512 255464 281518
rect 255412 281454 255464 281460
rect 255424 280673 255452 281454
rect 255502 281072 255558 281081
rect 255502 281007 255558 281016
rect 255410 280664 255466 280673
rect 255410 280599 255466 280608
rect 255240 280214 255360 280242
rect 255516 280226 255544 281007
rect 255504 280220 255556 280226
rect 255240 279154 255268 280214
rect 255504 280162 255556 280168
rect 255320 280152 255372 280158
rect 255320 280094 255372 280100
rect 255410 280120 255466 280129
rect 255332 279313 255360 280094
rect 255410 280055 255412 280064
rect 255464 280055 255466 280064
rect 255412 280026 255464 280032
rect 255608 279721 255636 284922
rect 255594 279712 255650 279721
rect 255594 279647 255650 279656
rect 255318 279304 255374 279313
rect 255318 279239 255374 279248
rect 255240 279126 255360 279154
rect 255332 278769 255360 279126
rect 255318 278760 255374 278769
rect 255318 278695 255374 278704
rect 255412 278520 255464 278526
rect 255412 278462 255464 278468
rect 255424 278361 255452 278462
rect 255410 278352 255466 278361
rect 255410 278287 255466 278296
rect 256606 278080 256662 278089
rect 256606 278015 256662 278024
rect 255410 277808 255466 277817
rect 255410 277743 255466 277752
rect 255424 277506 255452 277743
rect 255412 277500 255464 277506
rect 255412 277442 255464 277448
rect 255502 277400 255558 277409
rect 255502 277335 255558 277344
rect 255318 276992 255374 277001
rect 255318 276927 255374 276936
rect 255332 276078 255360 276927
rect 255516 276146 255544 277335
rect 256620 276457 256648 278015
rect 256606 276448 256662 276457
rect 256606 276383 256662 276392
rect 255504 276140 255556 276146
rect 255504 276082 255556 276088
rect 255320 276072 255372 276078
rect 255320 276014 255372 276020
rect 255412 276004 255464 276010
rect 255412 275946 255464 275952
rect 255424 275641 255452 275946
rect 255410 275632 255466 275641
rect 255410 275567 255466 275576
rect 255594 275088 255650 275097
rect 255594 275023 255650 275032
rect 255412 274644 255464 274650
rect 255412 274586 255464 274592
rect 255424 274281 255452 274586
rect 255410 274272 255466 274281
rect 255410 274207 255466 274216
rect 254030 273728 254086 273737
rect 254030 273663 254086 273672
rect 253938 273320 253994 273329
rect 253938 273255 253994 273264
rect 253938 272776 253994 272785
rect 253938 272711 253994 272720
rect 252926 269376 252982 269385
rect 252926 269311 252982 269320
rect 252834 267608 252890 267617
rect 252756 267566 252834 267594
rect 193402 258904 193458 258913
rect 193402 258839 193458 258848
rect 193416 258058 193444 258839
rect 193404 258052 193456 258058
rect 193404 257994 193456 258000
rect 193588 242956 193640 242962
rect 193588 242898 193640 242904
rect 193600 238754 193628 242898
rect 193678 242856 193734 242865
rect 193678 242791 193734 242800
rect 193692 241534 193720 242791
rect 251824 241936 251876 241942
rect 251824 241878 251876 241884
rect 250444 241868 250496 241874
rect 250444 241810 250496 241816
rect 193772 241596 193824 241602
rect 193772 241538 193824 241544
rect 193680 241528 193732 241534
rect 193680 241470 193732 241476
rect 193600 238726 193720 238754
rect 193692 234530 193720 238726
rect 193680 234524 193732 234530
rect 193680 234466 193732 234472
rect 193784 233238 193812 241538
rect 194796 240106 194824 241604
rect 194784 240100 194836 240106
rect 194784 240042 194836 240048
rect 197280 238678 197308 241604
rect 199764 241398 199792 241604
rect 199752 241392 199804 241398
rect 199752 241334 199804 241340
rect 197268 238672 197320 238678
rect 197268 238614 197320 238620
rect 193772 233232 193824 233238
rect 193772 233174 193824 233180
rect 199764 232558 199792 241334
rect 202248 235958 202276 241604
rect 204746 241590 204944 241618
rect 204916 240009 204944 241590
rect 204902 240000 204958 240009
rect 204902 239935 204958 239944
rect 206374 240000 206430 240009
rect 206374 239935 206430 239944
rect 202236 235952 202288 235958
rect 202236 235894 202288 235900
rect 202788 235952 202840 235958
rect 202788 235894 202840 235900
rect 202800 235278 202828 235894
rect 202788 235272 202840 235278
rect 202788 235214 202840 235220
rect 199752 232552 199804 232558
rect 199752 232494 199804 232500
rect 193220 229764 193272 229770
rect 193220 229706 193272 229712
rect 200762 227080 200818 227089
rect 200762 227015 200818 227024
rect 200776 213858 200804 227015
rect 200764 213852 200816 213858
rect 200764 213794 200816 213800
rect 195242 200696 195298 200705
rect 195242 200631 195298 200640
rect 193128 51740 193180 51746
rect 193128 51682 193180 51688
rect 188436 3460 188488 3466
rect 188436 3402 188488 3408
rect 152462 3360 152518 3369
rect 152462 3295 152518 3304
rect 195256 2106 195284 200631
rect 204916 185638 204944 239935
rect 206282 200696 206338 200705
rect 206282 200631 206338 200640
rect 204904 185632 204956 185638
rect 204904 185574 204956 185580
rect 198004 138712 198056 138718
rect 198004 138654 198056 138660
rect 198016 39370 198044 138654
rect 198096 100020 198148 100026
rect 198096 99962 198148 99968
rect 198004 39364 198056 39370
rect 198004 39306 198056 39312
rect 198108 6186 198136 99962
rect 206296 18698 206324 200631
rect 206388 61402 206416 239935
rect 207216 231742 207244 241604
rect 207204 231736 207256 231742
rect 207204 231678 207256 231684
rect 207664 231736 207716 231742
rect 207664 231678 207716 231684
rect 207676 230518 207704 231678
rect 207664 230512 207716 230518
rect 207664 230454 207716 230460
rect 207676 206990 207704 230454
rect 209792 227798 209820 241604
rect 212276 240038 212304 241604
rect 214760 241534 214788 241604
rect 217258 241590 217364 241618
rect 213920 241528 213972 241534
rect 213920 241470 213972 241476
rect 214748 241528 214800 241534
rect 214748 241470 214800 241476
rect 212264 240032 212316 240038
rect 212264 239974 212316 239980
rect 209780 227792 209832 227798
rect 209780 227734 209832 227740
rect 209792 220794 209820 227734
rect 209780 220788 209832 220794
rect 209780 220730 209832 220736
rect 213932 218754 213960 241470
rect 217336 234666 217364 241590
rect 217324 234660 217376 234666
rect 217324 234602 217376 234608
rect 213920 218748 213972 218754
rect 213920 218690 213972 218696
rect 217336 211070 217364 234602
rect 219728 234530 219756 241604
rect 220818 240136 220874 240145
rect 220818 240071 220874 240080
rect 219716 234524 219768 234530
rect 219716 234466 219768 234472
rect 217324 211064 217376 211070
rect 217324 211006 217376 211012
rect 207664 206984 207716 206990
rect 207664 206926 207716 206932
rect 213182 202872 213238 202881
rect 213182 202807 213238 202816
rect 206376 61396 206428 61402
rect 206376 61338 206428 61344
rect 213196 26926 213224 202807
rect 220084 98660 220136 98666
rect 220084 98602 220136 98608
rect 213184 26920 213236 26926
rect 213184 26862 213236 26868
rect 206284 18692 206336 18698
rect 206284 18634 206336 18640
rect 220096 18630 220124 98602
rect 220832 91769 220860 240071
rect 222212 223582 222240 241604
rect 224788 237318 224816 241604
rect 227272 240009 227300 241604
rect 227258 240000 227314 240009
rect 227258 239935 227314 239944
rect 224776 237312 224828 237318
rect 224776 237254 224828 237260
rect 229756 223650 229784 241604
rect 232240 238066 232268 241604
rect 234632 241590 234738 241618
rect 232228 238060 232280 238066
rect 232228 238002 232280 238008
rect 234632 228857 234660 241590
rect 234710 240136 234766 240145
rect 234710 240071 234766 240080
rect 234618 228848 234674 228857
rect 234618 228783 234674 228792
rect 234632 227050 234660 228783
rect 234620 227044 234672 227050
rect 234620 226986 234672 226992
rect 229744 223644 229796 223650
rect 229744 223586 229796 223592
rect 222200 223576 222252 223582
rect 222200 223518 222252 223524
rect 229756 205630 229784 223586
rect 234724 221474 234752 240071
rect 237208 233306 237236 241604
rect 239798 241590 240088 241618
rect 240060 238754 240088 241590
rect 240782 239456 240838 239465
rect 240782 239391 240838 239400
rect 240060 238726 240180 238754
rect 238666 238368 238722 238377
rect 238666 238303 238722 238312
rect 236644 233300 236696 233306
rect 236644 233242 236696 233248
rect 237196 233300 237248 233306
rect 237196 233242 237248 233248
rect 234712 221468 234764 221474
rect 234712 221410 234764 221416
rect 236656 208350 236684 233242
rect 238680 229129 238708 238303
rect 238666 229120 238722 229129
rect 238666 229055 238722 229064
rect 238666 228848 238722 228857
rect 238666 228783 238722 228792
rect 238680 219473 238708 228783
rect 238666 219464 238722 219473
rect 238666 219399 238722 219408
rect 238666 219056 238722 219065
rect 238666 218991 238722 219000
rect 238680 209817 238708 218991
rect 238666 209808 238722 209817
rect 238666 209743 238722 209752
rect 238666 209536 238722 209545
rect 238666 209471 238722 209480
rect 236644 208344 236696 208350
rect 236644 208286 236696 208292
rect 229744 205624 229796 205630
rect 229744 205566 229796 205572
rect 238680 200161 238708 209471
rect 240152 206242 240180 238726
rect 240796 222193 240824 239391
rect 241520 238060 241572 238066
rect 241520 238002 241572 238008
rect 240782 222184 240838 222193
rect 240782 222119 240838 222128
rect 241532 215218 241560 238002
rect 242268 222222 242296 241604
rect 243636 239420 243688 239426
rect 243636 239362 243688 239368
rect 243544 238060 243596 238066
rect 243544 238002 243596 238008
rect 242256 222216 242308 222222
rect 242256 222158 242308 222164
rect 242268 219434 242296 222158
rect 242176 219406 242296 219434
rect 242176 216578 242204 219406
rect 242164 216572 242216 216578
rect 242164 216514 242216 216520
rect 241520 215212 241572 215218
rect 241520 215154 241572 215160
rect 242164 215212 242216 215218
rect 242164 215154 242216 215160
rect 240140 206236 240192 206242
rect 240140 206178 240192 206184
rect 240784 206236 240836 206242
rect 240784 206178 240836 206184
rect 238666 200152 238722 200161
rect 238666 200087 238722 200096
rect 238666 199880 238722 199889
rect 238666 199815 238722 199824
rect 238680 190505 238708 199815
rect 238666 190496 238722 190505
rect 238666 190431 238722 190440
rect 238666 190360 238722 190369
rect 238666 190295 238722 190304
rect 238680 180849 238708 190295
rect 238666 180840 238722 180849
rect 238666 180775 238722 180784
rect 238666 180704 238722 180713
rect 238666 180639 238722 180648
rect 238680 171193 238708 180639
rect 238666 171184 238722 171193
rect 238666 171119 238722 171128
rect 238666 171048 238722 171057
rect 238666 170983 238722 170992
rect 238680 161537 238708 170983
rect 238666 161528 238722 161537
rect 238666 161463 238722 161472
rect 238666 161392 238722 161401
rect 238666 161327 238722 161336
rect 238680 151881 238708 161327
rect 238666 151872 238722 151881
rect 238666 151807 238722 151816
rect 238666 151736 238722 151745
rect 238666 151671 238722 151680
rect 238680 145625 238708 151671
rect 238666 145616 238722 145625
rect 238666 145551 238722 145560
rect 233148 101448 233200 101454
rect 233146 101416 233148 101425
rect 233200 101416 233202 101425
rect 233146 101351 233202 101360
rect 220818 91760 220874 91769
rect 220818 91695 220874 91704
rect 224224 53100 224276 53106
rect 224224 53042 224276 53048
rect 220084 18624 220136 18630
rect 220084 18566 220136 18572
rect 198096 6180 198148 6186
rect 198096 6122 198148 6128
rect 224236 3534 224264 53042
rect 231124 49020 231176 49026
rect 231124 48962 231176 48968
rect 231136 3913 231164 48962
rect 239310 4040 239366 4049
rect 239310 3975 239366 3984
rect 231122 3904 231178 3913
rect 231122 3839 231178 3848
rect 224224 3528 224276 3534
rect 224224 3470 224276 3476
rect 195244 2100 195296 2106
rect 195244 2042 195296 2048
rect 239324 480 239352 3975
rect 240506 3496 240562 3505
rect 240506 3431 240562 3440
rect 240520 480 240548 3431
rect 240796 2106 240824 206178
rect 241704 11756 241756 11762
rect 241704 11698 241756 11704
rect 240784 2100 240836 2106
rect 240784 2042 240836 2048
rect 241716 480 241744 11698
rect 242176 3369 242204 215154
rect 243556 213926 243584 238002
rect 243648 219434 243676 239362
rect 244278 237416 244334 237425
rect 244278 237351 244334 237360
rect 243636 219428 243688 219434
rect 243636 219370 243688 219376
rect 243544 213920 243596 213926
rect 243544 213862 243596 213868
rect 242992 51740 243044 51746
rect 242992 51682 243044 51688
rect 243004 16574 243032 51682
rect 243004 16546 244136 16574
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242162 3360 242218 3369
rect 242162 3295 242218 3304
rect 242912 480 242940 3402
rect 244108 480 244136 16546
rect 244292 3913 244320 237351
rect 244752 227730 244780 241604
rect 246394 239592 246450 239601
rect 246394 239527 246450 239536
rect 246304 235272 246356 235278
rect 246304 235214 246356 235220
rect 244740 227724 244792 227730
rect 244740 227666 244792 227672
rect 244752 221474 244780 227666
rect 244740 221468 244792 221474
rect 244740 221410 244792 221416
rect 244922 216744 244978 216753
rect 244922 216679 244978 216688
rect 244278 3904 244334 3913
rect 244278 3839 244334 3848
rect 244292 3641 244320 3839
rect 244278 3632 244334 3641
rect 244278 3567 244334 3576
rect 244936 3505 244964 216679
rect 245198 3632 245254 3641
rect 245198 3567 245254 3576
rect 244922 3496 244978 3505
rect 244922 3431 244978 3440
rect 245212 480 245240 3567
rect 246316 3466 246344 235214
rect 246408 216617 246436 239527
rect 247236 220794 247264 241604
rect 249168 241590 249734 241618
rect 249168 238814 249196 241590
rect 249248 241392 249300 241398
rect 249248 241334 249300 241340
rect 249156 238808 249208 238814
rect 249156 238750 249208 238756
rect 249062 237416 249118 237425
rect 249062 237351 249118 237360
rect 247224 220788 247276 220794
rect 247224 220730 247276 220736
rect 247684 220788 247736 220794
rect 247684 220730 247736 220736
rect 247696 219502 247724 220730
rect 247684 219496 247736 219502
rect 247684 219438 247736 219444
rect 246394 216608 246450 216617
rect 246394 216543 246450 216552
rect 247696 212498 247724 219438
rect 247684 212492 247736 212498
rect 247684 212434 247736 212440
rect 249076 198694 249104 237351
rect 249168 215966 249196 238750
rect 249260 227089 249288 241334
rect 250456 238513 250484 241810
rect 250534 241224 250590 241233
rect 250534 241159 250590 241168
rect 250442 238504 250498 238513
rect 250442 238439 250498 238448
rect 250444 232552 250496 232558
rect 250444 232494 250496 232500
rect 249246 227080 249302 227089
rect 249246 227015 249302 227024
rect 249156 215960 249208 215966
rect 249156 215902 249208 215908
rect 249064 198688 249116 198694
rect 249064 198630 249116 198636
rect 249062 138680 249118 138689
rect 249062 138615 249118 138624
rect 248420 48544 248472 48550
rect 248420 48486 248472 48492
rect 247592 6180 247644 6186
rect 247592 6122 247644 6128
rect 246396 3528 246448 3534
rect 246396 3470 246448 3476
rect 246304 3460 246356 3466
rect 246304 3402 246356 3408
rect 246408 480 246436 3470
rect 247604 480 247632 6122
rect 248432 490 248460 48486
rect 249076 42362 249104 138615
rect 249064 42356 249116 42362
rect 249064 42298 249116 42304
rect 249800 42356 249852 42362
rect 249800 42298 249852 42304
rect 249812 16574 249840 42298
rect 249812 16546 250024 16574
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 250456 3058 250484 232494
rect 250548 204241 250576 241159
rect 250628 240100 250680 240106
rect 250628 240042 250680 240048
rect 250640 212430 250668 240042
rect 251272 229764 251324 229770
rect 251272 229706 251324 229712
rect 250628 212424 250680 212430
rect 250628 212366 250680 212372
rect 250534 204232 250590 204241
rect 250534 204167 250590 204176
rect 251284 6914 251312 229706
rect 251836 226273 251864 241878
rect 252204 229094 252232 241604
rect 252652 239488 252704 239494
rect 252652 239430 252704 239436
rect 252664 238649 252692 239430
rect 252650 238640 252706 238649
rect 252650 238575 252706 238584
rect 251928 229066 252232 229094
rect 251822 226264 251878 226273
rect 251822 226199 251878 226208
rect 251928 225010 251956 229066
rect 251916 225004 251968 225010
rect 251916 224946 251968 224952
rect 251928 219337 251956 224946
rect 251914 219328 251970 219337
rect 251914 219263 251970 219272
rect 252756 208185 252784 267566
rect 252834 267543 252890 267552
rect 252940 258074 252968 269311
rect 252848 258046 252968 258074
rect 252848 237386 252876 258046
rect 252926 252512 252982 252521
rect 252926 252447 252982 252456
rect 252836 237380 252888 237386
rect 252836 237322 252888 237328
rect 252940 228410 252968 252447
rect 253202 247888 253258 247897
rect 253202 247823 253258 247832
rect 253110 246120 253166 246129
rect 253110 246055 253166 246064
rect 253018 243808 253074 243817
rect 253018 243743 253074 243752
rect 253032 242049 253060 243743
rect 253124 242894 253152 246055
rect 253216 245750 253244 247823
rect 253204 245744 253256 245750
rect 253204 245686 253256 245692
rect 253112 242888 253164 242894
rect 253112 242830 253164 242836
rect 253018 242040 253074 242049
rect 253018 241975 253074 241984
rect 253032 240106 253060 241975
rect 253124 241874 253152 242830
rect 253112 241868 253164 241874
rect 253112 241810 253164 241816
rect 253216 241398 253244 245686
rect 253204 241392 253256 241398
rect 253204 241334 253256 241340
rect 253020 240100 253072 240106
rect 253020 240042 253072 240048
rect 253204 236700 253256 236706
rect 253204 236642 253256 236648
rect 252928 228404 252980 228410
rect 252928 228346 252980 228352
rect 252742 208176 252798 208185
rect 252742 208111 252798 208120
rect 253216 77246 253244 236642
rect 253952 211138 253980 272711
rect 254044 234598 254072 273663
rect 255502 272368 255558 272377
rect 255502 272303 255558 272312
rect 255516 271998 255544 272303
rect 255504 271992 255556 271998
rect 255410 271960 255466 271969
rect 255504 271934 255556 271940
rect 255410 271895 255412 271904
rect 255464 271895 255466 271904
rect 255412 271866 255464 271872
rect 255320 271856 255372 271862
rect 255320 271798 255372 271804
rect 255332 271017 255360 271798
rect 255504 271652 255556 271658
rect 255504 271594 255556 271600
rect 255516 271425 255544 271594
rect 255502 271416 255558 271425
rect 255502 271351 255558 271360
rect 255318 271008 255374 271017
rect 255318 270943 255374 270952
rect 255410 270056 255466 270065
rect 255410 269991 255466 270000
rect 255424 269142 255452 269991
rect 255608 269822 255636 275023
rect 256606 274680 256662 274689
rect 256712 274666 256740 316678
rect 256804 295225 256832 328471
rect 258172 324352 258224 324358
rect 258172 324294 258224 324300
rect 256882 319424 256938 319433
rect 256882 319359 256938 319368
rect 256790 295216 256846 295225
rect 256790 295151 256846 295160
rect 256804 294098 256832 295151
rect 256792 294092 256844 294098
rect 256792 294034 256844 294040
rect 256896 285705 256924 319359
rect 258080 311908 258132 311914
rect 258080 311850 258132 311856
rect 256976 308440 257028 308446
rect 256976 308382 257028 308388
rect 256988 292126 257016 308382
rect 257344 294092 257396 294098
rect 257344 294034 257396 294040
rect 256976 292120 257028 292126
rect 256976 292062 257028 292068
rect 256882 285696 256938 285705
rect 256882 285631 256938 285640
rect 257356 276049 257384 294034
rect 258092 278526 258120 311850
rect 258184 290902 258212 324294
rect 258276 299402 258304 332551
rect 259644 329112 259696 329118
rect 259644 329054 259696 329060
rect 259552 321700 259604 321706
rect 259552 321642 259604 321648
rect 258356 314696 258408 314702
rect 258356 314638 258408 314644
rect 258264 299396 258316 299402
rect 258264 299338 258316 299344
rect 258172 290896 258224 290902
rect 258172 290838 258224 290844
rect 258368 282810 258396 314638
rect 259460 305652 259512 305658
rect 259460 305594 259512 305600
rect 259368 299396 259420 299402
rect 259368 299338 259420 299344
rect 259380 298790 259408 299338
rect 259368 298784 259420 298790
rect 259368 298726 259420 298732
rect 259368 295384 259420 295390
rect 259368 295326 259420 295332
rect 258356 282804 258408 282810
rect 258356 282746 258408 282752
rect 259380 278730 259408 295326
rect 259368 278724 259420 278730
rect 259368 278666 259420 278672
rect 258080 278520 258132 278526
rect 258080 278462 258132 278468
rect 258172 277500 258224 277506
rect 258172 277442 258224 277448
rect 257066 276040 257122 276049
rect 257066 275975 257122 275984
rect 257342 276040 257398 276049
rect 257342 275975 257398 275984
rect 258078 276040 258134 276049
rect 258078 275975 258134 275984
rect 256662 274638 256740 274666
rect 256606 274615 256662 274624
rect 255964 273964 256016 273970
rect 255964 273906 256016 273912
rect 255596 269816 255648 269822
rect 255596 269758 255648 269764
rect 255412 269136 255464 269142
rect 255412 269078 255464 269084
rect 255502 269104 255558 269113
rect 255502 269039 255558 269048
rect 255516 267782 255544 269039
rect 255504 267776 255556 267782
rect 255976 267734 256004 273906
rect 256698 272504 256754 272513
rect 256698 272439 256754 272448
rect 256514 269784 256570 269793
rect 256514 269719 256570 269728
rect 255504 267718 255556 267724
rect 255412 267708 255464 267714
rect 255412 267650 255464 267656
rect 255884 267706 256004 267734
rect 255424 267345 255452 267650
rect 255410 267336 255466 267345
rect 255410 267271 255466 267280
rect 255412 267028 255464 267034
rect 255412 266970 255464 266976
rect 255424 266937 255452 266970
rect 255410 266928 255466 266937
rect 255410 266863 255466 266872
rect 255502 266520 255558 266529
rect 255502 266455 255558 266464
rect 255320 266348 255372 266354
rect 255320 266290 255372 266296
rect 255332 265577 255360 266290
rect 255318 265568 255374 265577
rect 255318 265503 255374 265512
rect 255412 263696 255464 263702
rect 255410 263664 255412 263673
rect 255464 263664 255466 263673
rect 255410 263599 255466 263608
rect 255412 263560 255464 263566
rect 255412 263502 255464 263508
rect 255424 263265 255452 263502
rect 255410 263256 255466 263265
rect 255410 263191 255466 263200
rect 255410 259584 255466 259593
rect 255410 259519 255466 259528
rect 255424 259486 255452 259519
rect 255412 259480 255464 259486
rect 255412 259422 255464 259428
rect 255410 259040 255466 259049
rect 255410 258975 255466 258984
rect 255424 258126 255452 258975
rect 255516 258641 255544 266455
rect 255884 260001 255912 267706
rect 256528 266393 256556 269719
rect 256606 268696 256662 268705
rect 256712 268682 256740 272439
rect 256662 268654 256740 268682
rect 256606 268631 256662 268640
rect 256514 266384 256570 266393
rect 256514 266319 256570 266328
rect 255964 265668 256016 265674
rect 255964 265610 256016 265616
rect 255870 259992 255926 260001
rect 255870 259927 255926 259936
rect 255502 258632 255558 258641
rect 255502 258567 255558 258576
rect 255412 258120 255464 258126
rect 255412 258062 255464 258068
rect 255410 257680 255466 257689
rect 255410 257615 255466 257624
rect 255424 257446 255452 257615
rect 255412 257440 255464 257446
rect 255412 257382 255464 257388
rect 255688 257372 255740 257378
rect 255688 257314 255740 257320
rect 255504 256692 255556 256698
rect 255504 256634 255556 256640
rect 255410 256320 255466 256329
rect 255410 256255 255466 256264
rect 255424 256018 255452 256255
rect 255412 256012 255464 256018
rect 255412 255954 255464 255960
rect 255516 255921 255544 256634
rect 255502 255912 255558 255921
rect 255502 255847 255558 255856
rect 255410 254960 255466 254969
rect 255410 254895 255466 254904
rect 255424 254046 255452 254895
rect 255594 254552 255650 254561
rect 255594 254487 255650 254496
rect 255412 254040 255464 254046
rect 255412 253982 255464 253988
rect 255320 253972 255372 253978
rect 255320 253914 255372 253920
rect 255332 251297 255360 253914
rect 255502 253600 255558 253609
rect 255502 253535 255558 253544
rect 255410 253192 255466 253201
rect 255410 253127 255466 253136
rect 255424 252686 255452 253127
rect 255412 252680 255464 252686
rect 255412 252622 255464 252628
rect 255516 252618 255544 253535
rect 255504 252612 255556 252618
rect 255504 252554 255556 252560
rect 255502 252240 255558 252249
rect 255502 252175 255558 252184
rect 255410 251832 255466 251841
rect 255410 251767 255466 251776
rect 255424 251598 255452 251767
rect 255412 251592 255464 251598
rect 255412 251534 255464 251540
rect 255318 251288 255374 251297
rect 255516 251258 255544 252175
rect 255318 251223 255374 251232
rect 255504 251252 255556 251258
rect 255504 251194 255556 251200
rect 255318 250336 255374 250345
rect 255318 250271 255374 250280
rect 255332 249898 255360 250271
rect 255410 249928 255466 249937
rect 255320 249892 255372 249898
rect 255410 249863 255466 249872
rect 255320 249834 255372 249840
rect 255424 249830 255452 249863
rect 255412 249824 255464 249830
rect 255412 249766 255464 249772
rect 254582 249248 254638 249257
rect 254582 249183 254638 249192
rect 254596 247722 254624 249183
rect 255318 248976 255374 248985
rect 255318 248911 255374 248920
rect 255332 248538 255360 248911
rect 255320 248532 255372 248538
rect 255320 248474 255372 248480
rect 254584 247716 254636 247722
rect 254584 247658 254636 247664
rect 254124 244996 254176 245002
rect 254124 244938 254176 244944
rect 254136 241942 254164 244938
rect 254124 241936 254176 241942
rect 254124 241878 254176 241884
rect 254596 239426 254624 247658
rect 255410 247616 255466 247625
rect 255410 247551 255466 247560
rect 255424 247110 255452 247551
rect 255412 247104 255464 247110
rect 255412 247046 255464 247052
rect 255318 246800 255374 246809
rect 255318 246735 255374 246744
rect 255332 244361 255360 246735
rect 255424 245970 255452 247046
rect 255424 245942 255544 245970
rect 255410 245848 255466 245857
rect 255410 245783 255466 245792
rect 255424 245682 255452 245783
rect 255412 245676 255464 245682
rect 255412 245618 255464 245624
rect 255516 245426 255544 245942
rect 255424 245398 255544 245426
rect 255318 244352 255374 244361
rect 255318 244287 255374 244296
rect 255424 243658 255452 245398
rect 255502 245304 255558 245313
rect 255502 245239 255558 245248
rect 255332 243630 255452 243658
rect 255332 242842 255360 243630
rect 255516 243574 255544 245239
rect 255608 245002 255636 254487
rect 255700 252657 255728 257314
rect 255976 254561 256004 265610
rect 256606 264072 256662 264081
rect 256662 264030 256740 264058
rect 256606 264007 256662 264016
rect 256712 258074 256740 264030
rect 256882 261352 256938 261361
rect 256882 261287 256938 261296
rect 256712 258046 256832 258074
rect 255962 254552 256018 254561
rect 255962 254487 256018 254496
rect 255686 252648 255742 252657
rect 255686 252583 255742 252592
rect 255686 248568 255742 248577
rect 255686 248503 255742 248512
rect 255700 248470 255728 248503
rect 255688 248464 255740 248470
rect 255688 248406 255740 248412
rect 255596 244996 255648 245002
rect 255596 244938 255648 244944
rect 255594 244896 255650 244905
rect 255594 244831 255650 244840
rect 255504 243568 255556 243574
rect 255410 243536 255466 243545
rect 255504 243510 255556 243516
rect 255410 243471 255466 243480
rect 255424 242962 255452 243471
rect 255412 242956 255464 242962
rect 255412 242898 255464 242904
rect 255332 242814 255544 242842
rect 255318 242584 255374 242593
rect 255318 242519 255374 242528
rect 255332 241466 255360 242519
rect 255412 242208 255464 242214
rect 255412 242150 255464 242156
rect 255424 242049 255452 242150
rect 255410 242040 255466 242049
rect 255410 241975 255466 241984
rect 255410 241768 255466 241777
rect 255410 241703 255466 241712
rect 255424 241534 255452 241703
rect 255412 241528 255464 241534
rect 255412 241470 255464 241476
rect 255320 241460 255372 241466
rect 255320 241402 255372 241408
rect 255332 240786 255360 241402
rect 255516 241346 255544 242814
rect 255424 241318 255544 241346
rect 255320 240780 255372 240786
rect 255320 240722 255372 240728
rect 254584 239420 254636 239426
rect 254584 239362 254636 239368
rect 255424 235793 255452 241318
rect 255608 238754 255636 244831
rect 255688 244384 255740 244390
rect 255688 244326 255740 244332
rect 255700 242894 255728 244326
rect 255688 242888 255740 242894
rect 255688 242830 255740 242836
rect 255962 242176 256018 242185
rect 255962 242111 256018 242120
rect 255516 238726 255636 238754
rect 255410 235784 255466 235793
rect 255410 235719 255466 235728
rect 254032 234592 254084 234598
rect 254032 234534 254084 234540
rect 255516 230625 255544 238726
rect 255976 231878 256004 242111
rect 255964 231872 256016 231878
rect 255964 231814 256016 231820
rect 255502 230616 255558 230625
rect 255502 230551 255558 230560
rect 255516 228410 255544 230551
rect 255504 228404 255556 228410
rect 255504 228346 255556 228352
rect 255976 224942 256004 231814
rect 256804 231810 256832 258046
rect 256896 241369 256924 261287
rect 256882 241360 256938 241369
rect 256882 241295 256938 241304
rect 256792 231804 256844 231810
rect 256792 231746 256844 231752
rect 256056 227792 256108 227798
rect 256056 227734 256108 227740
rect 255964 224936 256016 224942
rect 255964 224878 256016 224884
rect 253940 211132 253992 211138
rect 253940 211074 253992 211080
rect 255320 113824 255372 113830
rect 255320 113766 255372 113772
rect 252560 77240 252612 77246
rect 252560 77182 252612 77188
rect 253204 77240 253256 77246
rect 253204 77182 253256 77188
rect 252572 48550 252600 77182
rect 253204 58676 253256 58682
rect 253204 58618 253256 58624
rect 252560 48544 252612 48550
rect 252560 48486 252612 48492
rect 253216 17270 253244 58618
rect 253204 17264 253256 17270
rect 253204 17206 253256 17212
rect 255332 16574 255360 113766
rect 255332 16546 255912 16574
rect 251192 6886 251312 6914
rect 250444 3052 250496 3058
rect 250444 2994 250496 3000
rect 251192 480 251220 6886
rect 254674 3496 254730 3505
rect 253480 3460 253532 3466
rect 254674 3431 254730 3440
rect 253480 3402 253532 3408
rect 252376 3052 252428 3058
rect 252376 2994 252428 3000
rect 252388 480 252416 2994
rect 253492 480 253520 3402
rect 254688 480 254716 3431
rect 255884 480 255912 16546
rect 256068 3466 256096 227734
rect 257080 206961 257108 275975
rect 257066 206952 257122 206961
rect 257066 206887 257122 206896
rect 258092 16574 258120 275975
rect 258184 238066 258212 277442
rect 259472 271658 259500 305594
rect 259564 288017 259592 321642
rect 259656 295390 259684 329054
rect 259736 310548 259788 310554
rect 259736 310490 259788 310496
rect 259644 295384 259696 295390
rect 259644 295326 259696 295332
rect 259550 288008 259606 288017
rect 259550 287943 259606 287952
rect 259552 284572 259604 284578
rect 259552 284514 259604 284520
rect 259460 271652 259512 271658
rect 259460 271594 259512 271600
rect 258356 256692 258408 256698
rect 258356 256634 258408 256640
rect 258368 256057 258396 256634
rect 258354 256048 258410 256057
rect 258354 255983 258410 255992
rect 258354 247208 258410 247217
rect 258354 247143 258410 247152
rect 258264 245676 258316 245682
rect 258264 245618 258316 245624
rect 258172 238060 258224 238066
rect 258172 238002 258224 238008
rect 258276 213897 258304 245618
rect 258368 238814 258396 247143
rect 258356 238808 258408 238814
rect 258356 238750 258408 238756
rect 258368 235929 258396 238750
rect 258354 235920 258410 235929
rect 258354 235855 258410 235864
rect 259564 233238 259592 284514
rect 259748 280090 259776 310490
rect 260116 305046 260144 349114
rect 261484 342304 261536 342310
rect 261484 342246 261536 342252
rect 260932 323604 260984 323610
rect 260932 323546 260984 323552
rect 260840 313948 260892 313954
rect 260840 313890 260892 313896
rect 260104 305040 260156 305046
rect 260104 304982 260156 304988
rect 259736 280084 259788 280090
rect 259736 280026 259788 280032
rect 259828 278724 259880 278730
rect 259828 278666 259880 278672
rect 259642 270600 259698 270609
rect 259642 270535 259698 270544
rect 259552 233232 259604 233238
rect 259552 233174 259604 233180
rect 259656 224913 259684 270535
rect 259736 251864 259788 251870
rect 259736 251806 259788 251812
rect 259748 239465 259776 251806
rect 259734 239456 259790 239465
rect 259734 239391 259790 239400
rect 259642 224904 259698 224913
rect 259642 224839 259698 224848
rect 258262 213888 258318 213897
rect 258262 213823 258318 213832
rect 259552 185632 259604 185638
rect 259552 185574 259604 185580
rect 258092 16546 258304 16574
rect 257068 4820 257120 4826
rect 257068 4762 257120 4768
rect 256056 3460 256108 3466
rect 256056 3402 256108 3408
rect 257080 480 257108 4762
rect 258276 480 258304 16546
rect 259564 6914 259592 185574
rect 259840 16574 259868 278666
rect 260852 274650 260880 313890
rect 260944 289746 260972 323546
rect 261024 310616 261076 310622
rect 261024 310558 261076 310564
rect 260932 289740 260984 289746
rect 260932 289682 260984 289688
rect 261036 284306 261064 310558
rect 261496 298042 261524 342246
rect 263690 332752 263746 332761
rect 263690 332687 263746 332696
rect 262402 331256 262458 331265
rect 262402 331191 262458 331200
rect 262310 320784 262366 320793
rect 262310 320719 262366 320728
rect 261484 298036 261536 298042
rect 261484 297978 261536 297984
rect 262220 298036 262272 298042
rect 262220 297978 262272 297984
rect 262128 297424 262180 297430
rect 262126 297392 262128 297401
rect 262180 297392 262182 297401
rect 262126 297327 262182 297336
rect 261482 296032 261538 296041
rect 261482 295967 261538 295976
rect 261024 284300 261076 284306
rect 261024 284242 261076 284248
rect 261496 275398 261524 295967
rect 262232 293894 262260 297978
rect 262220 293888 262272 293894
rect 262220 293830 262272 293836
rect 261484 275392 261536 275398
rect 261484 275334 261536 275340
rect 260840 274644 260892 274650
rect 260840 274586 260892 274592
rect 260932 269136 260984 269142
rect 260932 269078 260984 269084
rect 260840 259480 260892 259486
rect 260840 259422 260892 259428
rect 260746 244352 260802 244361
rect 260746 244287 260748 244296
rect 260800 244287 260802 244296
rect 260748 244258 260800 244264
rect 260852 211041 260880 259422
rect 260944 233073 260972 269078
rect 261116 267776 261168 267782
rect 261116 267718 261168 267724
rect 261024 243024 261076 243030
rect 261024 242966 261076 242972
rect 260930 233064 260986 233073
rect 260930 232999 260986 233008
rect 261036 215286 261064 242966
rect 261128 239494 261156 267718
rect 262220 267028 262272 267034
rect 262220 266970 262272 266976
rect 262232 266529 262260 266970
rect 262218 266520 262274 266529
rect 262218 266455 262274 266464
rect 262220 263696 262272 263702
rect 262220 263638 262272 263644
rect 261116 239488 261168 239494
rect 261116 239430 261168 239436
rect 261024 215280 261076 215286
rect 261024 215222 261076 215228
rect 262232 212537 262260 263638
rect 262324 263566 262352 320719
rect 262416 297401 262444 331191
rect 263600 320204 263652 320210
rect 263600 320146 263652 320152
rect 262496 307828 262548 307834
rect 262496 307770 262548 307776
rect 262402 297392 262458 297401
rect 262402 297327 262458 297336
rect 262508 281518 262536 307770
rect 262588 301164 262640 301170
rect 262588 301106 262640 301112
rect 262496 281512 262548 281518
rect 262496 281454 262548 281460
rect 262312 263560 262364 263566
rect 262312 263502 262364 263508
rect 262494 251832 262550 251841
rect 262494 251767 262550 251776
rect 262508 251258 262536 251767
rect 262496 251252 262548 251258
rect 262496 251194 262548 251200
rect 262404 243568 262456 243574
rect 262404 243510 262456 243516
rect 262416 242962 262444 243510
rect 262404 242956 262456 242962
rect 262404 242898 262456 242904
rect 262218 212528 262274 212537
rect 262218 212463 262274 212472
rect 260838 211032 260894 211041
rect 260838 210967 260894 210976
rect 262416 204270 262444 242898
rect 262508 228993 262536 251194
rect 262494 228984 262550 228993
rect 262494 228919 262550 228928
rect 262404 204264 262456 204270
rect 262404 204206 262456 204212
rect 259840 16546 260696 16574
rect 259472 6886 259592 6914
rect 259472 480 259500 6886
rect 260668 480 260696 16546
rect 261760 6180 261812 6186
rect 261760 6122 261812 6128
rect 261772 480 261800 6122
rect 262600 490 262628 301106
rect 263612 282305 263640 320146
rect 263704 299470 263732 332687
rect 265164 321632 265216 321638
rect 265070 321600 265126 321609
rect 265164 321574 265216 321580
rect 265070 321535 265126 321544
rect 264980 316056 265032 316062
rect 264980 315998 265032 316004
rect 263782 312080 263838 312089
rect 263782 312015 263838 312024
rect 263692 299464 263744 299470
rect 263692 299406 263744 299412
rect 263704 298178 263732 299406
rect 263692 298172 263744 298178
rect 263692 298114 263744 298120
rect 263692 294024 263744 294030
rect 263692 293966 263744 293972
rect 263598 282296 263654 282305
rect 263598 282231 263654 282240
rect 263600 276140 263652 276146
rect 263600 276082 263652 276088
rect 262680 258052 262732 258058
rect 262680 257994 262732 258000
rect 262692 257446 262720 257994
rect 262680 257440 262732 257446
rect 262680 257382 262732 257388
rect 262692 256737 262720 257382
rect 262678 256728 262734 256737
rect 262678 256663 262734 256672
rect 263612 205562 263640 276082
rect 263704 236706 263732 293966
rect 263796 280158 263824 312015
rect 263876 305040 263928 305046
rect 263876 304982 263928 304988
rect 263888 293962 263916 304982
rect 263876 293956 263928 293962
rect 263876 293898 263928 293904
rect 263784 280152 263836 280158
rect 263784 280094 263836 280100
rect 264992 276010 265020 315998
rect 265084 287026 265112 321535
rect 265176 288318 265204 321574
rect 266372 309806 266400 697546
rect 266452 339516 266504 339522
rect 266452 339458 266504 339464
rect 266360 309800 266412 309806
rect 266360 309742 266412 309748
rect 265164 288312 265216 288318
rect 265164 288254 265216 288260
rect 265072 287020 265124 287026
rect 265072 286962 265124 286968
rect 265256 276072 265308 276078
rect 265256 276014 265308 276020
rect 264980 276004 265032 276010
rect 264980 275946 265032 275952
rect 265072 271924 265124 271930
rect 265072 271866 265124 271872
rect 263876 252340 263928 252346
rect 263876 252282 263928 252288
rect 263888 250617 263916 252282
rect 263874 250608 263930 250617
rect 263874 250543 263930 250552
rect 263784 241528 263836 241534
rect 263784 241470 263836 241476
rect 263692 236700 263744 236706
rect 263692 236642 263744 236648
rect 263600 205556 263652 205562
rect 263600 205498 263652 205504
rect 263796 202842 263824 241470
rect 263888 230450 263916 250543
rect 263876 230444 263928 230450
rect 263876 230386 263928 230392
rect 265084 226302 265112 271866
rect 265164 250504 265216 250510
rect 265164 250446 265216 250452
rect 265176 249898 265204 250446
rect 265164 249892 265216 249898
rect 265164 249834 265216 249840
rect 265072 226296 265124 226302
rect 265072 226238 265124 226244
rect 265176 223514 265204 249834
rect 265164 223508 265216 223514
rect 265164 223450 265216 223456
rect 265268 208282 265296 276014
rect 266372 272513 266400 309742
rect 266358 272504 266414 272513
rect 266358 272439 266414 272448
rect 266464 269793 266492 339458
rect 267832 329860 267884 329866
rect 267832 329802 267884 329808
rect 266544 327140 266596 327146
rect 266544 327082 266596 327088
rect 266556 271862 266584 327082
rect 267740 320272 267792 320278
rect 267740 320214 267792 320220
rect 266636 313336 266688 313342
rect 266636 313278 266688 313284
rect 266648 282878 266676 313278
rect 267752 284986 267780 320214
rect 267844 296682 267872 329802
rect 267832 296676 267884 296682
rect 267832 296618 267884 296624
rect 267740 284980 267792 284986
rect 267740 284922 267792 284928
rect 266636 282872 266688 282878
rect 266636 282814 266688 282820
rect 267004 271924 267056 271930
rect 267004 271866 267056 271872
rect 266544 271856 266596 271862
rect 266544 271798 266596 271804
rect 266450 269784 266506 269793
rect 266450 269719 266506 269728
rect 266358 264344 266414 264353
rect 266358 264279 266414 264288
rect 266372 215257 266400 264279
rect 266636 258800 266688 258806
rect 266636 258742 266688 258748
rect 266648 258126 266676 258742
rect 266636 258120 266688 258126
rect 267016 258074 267044 271866
rect 268396 264897 268424 702986
rect 269764 700324 269816 700330
rect 269764 700266 269816 700272
rect 269120 343732 269172 343738
rect 269120 343674 269172 343680
rect 268476 298172 268528 298178
rect 268476 298114 268528 298120
rect 268382 264888 268438 264897
rect 268382 264823 268438 264832
rect 268384 262880 268436 262886
rect 268384 262822 268436 262828
rect 267924 258732 267976 258738
rect 267924 258674 267976 258680
rect 266636 258062 266688 258068
rect 266452 252680 266504 252686
rect 266452 252622 266504 252628
rect 266358 215248 266414 215257
rect 266358 215183 266414 215192
rect 266464 209098 266492 252622
rect 266544 249824 266596 249830
rect 266544 249766 266596 249772
rect 266556 222154 266584 249766
rect 266648 240825 266676 258062
rect 266924 258046 267044 258074
rect 266924 252346 266952 258046
rect 267830 257272 267886 257281
rect 267830 257207 267886 257216
rect 267740 254040 267792 254046
rect 267740 253982 267792 253988
rect 267004 253904 267056 253910
rect 267004 253846 267056 253852
rect 267016 252686 267044 253846
rect 267004 252680 267056 252686
rect 267004 252622 267056 252628
rect 266912 252340 266964 252346
rect 266912 252282 266964 252288
rect 266634 240816 266690 240825
rect 266634 240751 266690 240760
rect 267004 234660 267056 234666
rect 267004 234602 267056 234608
rect 266544 222148 266596 222154
rect 266544 222090 266596 222096
rect 266452 209092 266504 209098
rect 266452 209034 266504 209040
rect 265256 208276 265308 208282
rect 265256 208218 265308 208224
rect 263784 202836 263836 202842
rect 263784 202778 263836 202784
rect 264244 112464 264296 112470
rect 264244 112406 264296 112412
rect 262864 39364 262916 39370
rect 262864 39306 262916 39312
rect 262876 11762 262904 39306
rect 262864 11756 262916 11762
rect 262864 11698 262916 11704
rect 264256 4826 264284 112406
rect 266360 54528 266412 54534
rect 266360 54470 266412 54476
rect 266372 16574 266400 54470
rect 266372 16546 266584 16574
rect 264244 4820 264296 4826
rect 264244 4762 264296 4768
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262600 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 3470
rect 265348 3460 265400 3466
rect 265348 3402 265400 3408
rect 265360 480 265388 3402
rect 266556 480 266584 16546
rect 267016 3466 267044 234602
rect 267752 216646 267780 253982
rect 267740 216640 267792 216646
rect 267740 216582 267792 216588
rect 267844 194546 267872 257207
rect 267936 254561 267964 258674
rect 267922 254552 267978 254561
rect 267922 254487 267978 254496
rect 267936 220833 267964 254487
rect 268396 253910 268424 262822
rect 268488 261526 268516 298114
rect 269028 296676 269080 296682
rect 269028 296618 269080 296624
rect 269040 296002 269068 296618
rect 269028 295996 269080 296002
rect 269028 295938 269080 295944
rect 269132 288386 269160 343674
rect 269212 331288 269264 331294
rect 269212 331230 269264 331236
rect 269224 298110 269252 331230
rect 269212 298104 269264 298110
rect 269212 298046 269264 298052
rect 269120 288380 269172 288386
rect 269120 288322 269172 288328
rect 269120 275392 269172 275398
rect 269120 275334 269172 275340
rect 268566 264208 268622 264217
rect 268566 264143 268622 264152
rect 268476 261520 268528 261526
rect 268476 261462 268528 261468
rect 268580 257281 268608 264143
rect 268566 257272 268622 257281
rect 268566 257207 268622 257216
rect 269028 254584 269080 254590
rect 269028 254526 269080 254532
rect 269040 254046 269068 254526
rect 269028 254040 269080 254046
rect 269028 253982 269080 253988
rect 268384 253904 268436 253910
rect 268384 253846 268436 253852
rect 268016 248532 268068 248538
rect 268016 248474 268068 248480
rect 268028 224777 268056 248474
rect 268014 224768 268070 224777
rect 268014 224703 268070 224712
rect 268382 224768 268438 224777
rect 268382 224703 268438 224712
rect 267922 220824 267978 220833
rect 267922 220759 267978 220768
rect 268396 219434 268424 224703
rect 268384 219428 268436 219434
rect 268384 219370 268436 219376
rect 267924 218748 267976 218754
rect 267924 218690 267976 218696
rect 267832 194540 267884 194546
rect 267832 194482 267884 194488
rect 267832 133204 267884 133210
rect 267832 133146 267884 133152
rect 267844 6914 267872 133146
rect 267936 16574 267964 218690
rect 269132 56574 269160 275334
rect 269212 271992 269264 271998
rect 269212 271934 269264 271940
rect 269224 195974 269252 271934
rect 269776 268433 269804 700266
rect 270592 345092 270644 345098
rect 270592 345034 270644 345040
rect 270500 300892 270552 300898
rect 270500 300834 270552 300840
rect 270408 298104 270460 298110
rect 270408 298046 270460 298052
rect 270420 297430 270448 298046
rect 270408 297424 270460 297430
rect 270408 297366 270460 297372
rect 269762 268424 269818 268433
rect 269762 268359 269818 268368
rect 269302 260128 269358 260137
rect 269302 260063 269358 260072
rect 269316 219201 269344 260063
rect 269776 258074 269804 268359
rect 269408 258046 269804 258074
rect 269408 230489 269436 258046
rect 269394 230480 269450 230489
rect 269394 230415 269450 230424
rect 269302 219192 269358 219201
rect 269302 219127 269358 219136
rect 269212 195968 269264 195974
rect 269212 195910 269264 195916
rect 269120 56568 269172 56574
rect 269120 56510 269172 56516
rect 269132 16574 269160 56510
rect 267936 16546 268424 16574
rect 269132 16546 270080 16574
rect 267752 6886 267872 6914
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267752 480 267780 6886
rect 268396 490 268424 16546
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 16546
rect 270512 6186 270540 300834
rect 270604 289814 270632 345034
rect 270592 289808 270644 289814
rect 270592 289750 270644 289756
rect 271156 265577 271184 703122
rect 276664 703112 276716 703118
rect 276664 703054 276716 703060
rect 272064 346452 272116 346458
rect 272064 346394 272116 346400
rect 271972 341012 272024 341018
rect 271972 340954 272024 340960
rect 271984 291174 272012 340954
rect 271972 291168 272024 291174
rect 271972 291110 272024 291116
rect 271880 280220 271932 280226
rect 271880 280162 271932 280168
rect 271142 265568 271198 265577
rect 271142 265503 271198 265512
rect 271788 260160 271840 260166
rect 271788 260102 271840 260108
rect 270776 256012 270828 256018
rect 270776 255954 270828 255960
rect 270788 255542 270816 255954
rect 271800 255542 271828 260102
rect 270776 255536 270828 255542
rect 270776 255478 270828 255484
rect 271788 255536 271840 255542
rect 271788 255478 271840 255484
rect 270684 252612 270736 252618
rect 270684 252554 270736 252560
rect 270592 230512 270644 230518
rect 270592 230454 270644 230460
rect 270500 6180 270552 6186
rect 270500 6122 270552 6128
rect 270604 3534 270632 230454
rect 270696 205601 270724 252554
rect 270788 223553 270816 255478
rect 271788 253224 271840 253230
rect 271788 253166 271840 253172
rect 271800 252618 271828 253166
rect 271788 252612 271840 252618
rect 271788 252554 271840 252560
rect 270774 223544 270830 223553
rect 270774 223479 270830 223488
rect 271892 209166 271920 280162
rect 272076 278089 272104 346394
rect 276676 310457 276704 703054
rect 283852 700330 283880 703520
rect 300136 702982 300164 703520
rect 300124 702976 300176 702982
rect 300124 702918 300176 702924
rect 332520 700330 332548 703520
rect 348804 702681 348832 703520
rect 364996 702914 365024 703520
rect 397472 703186 397500 703520
rect 397460 703180 397512 703186
rect 397460 703122 397512 703128
rect 413664 703118 413692 703520
rect 413652 703112 413704 703118
rect 413652 703054 413704 703060
rect 364984 702908 365036 702914
rect 364984 702850 365036 702856
rect 429856 702846 429884 703520
rect 462332 703050 462360 703520
rect 462320 703044 462372 703050
rect 462320 702986 462372 702992
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 478524 702778 478552 703520
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 494808 702710 494836 703520
rect 494796 702704 494848 702710
rect 348790 702672 348846 702681
rect 494796 702646 494848 702652
rect 527192 702642 527220 703520
rect 348790 702607 348846 702616
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 543476 702545 543504 703520
rect 543462 702536 543518 702545
rect 559668 702506 559696 703520
rect 582472 702568 582524 702574
rect 582472 702510 582524 702516
rect 543462 702471 543518 702480
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 286324 700324 286376 700330
rect 286324 700266 286376 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 276018 310448 276074 310457
rect 276018 310383 276074 310392
rect 276662 310448 276718 310457
rect 276662 310383 276718 310392
rect 276032 309369 276060 310383
rect 276018 309360 276074 309369
rect 276018 309295 276074 309304
rect 273260 302932 273312 302938
rect 273260 302874 273312 302880
rect 272062 278080 272118 278089
rect 272062 278015 272118 278024
rect 271972 248464 272024 248470
rect 271972 248406 272024 248412
rect 271880 209160 271932 209166
rect 271880 209102 271932 209108
rect 270682 205592 270738 205601
rect 270682 205527 270738 205536
rect 271984 201482 272012 248406
rect 271972 201476 272024 201482
rect 271972 201418 272024 201424
rect 273272 159390 273300 302874
rect 274640 299600 274692 299606
rect 274640 299542 274692 299548
rect 273352 269816 273404 269822
rect 273352 269758 273404 269764
rect 273364 208321 273392 269758
rect 273442 267064 273498 267073
rect 273442 266999 273498 267008
rect 273456 266393 273484 266999
rect 273442 266384 273498 266393
rect 273442 266319 273498 266328
rect 273456 218006 273484 266319
rect 273444 218000 273496 218006
rect 273444 217942 273496 217948
rect 273350 208312 273406 208321
rect 273350 208247 273406 208256
rect 273260 159384 273312 159390
rect 273260 159326 273312 159332
rect 270592 3528 270644 3534
rect 270592 3470 270644 3476
rect 271236 3460 271288 3466
rect 271236 3402 271288 3408
rect 271248 480 271276 3402
rect 272432 3256 272484 3262
rect 272432 3198 272484 3204
rect 272444 480 272472 3198
rect 273272 490 273300 159326
rect 273904 109744 273956 109750
rect 273904 109686 273956 109692
rect 273916 13122 273944 109686
rect 274652 84153 274680 299542
rect 276032 266354 276060 309295
rect 286336 309097 286364 700266
rect 582484 670721 582512 702510
rect 583574 696960 583630 696969
rect 583574 696895 583630 696904
rect 582654 683904 582710 683913
rect 582654 683839 582710 683848
rect 582470 670712 582526 670721
rect 582470 670647 582526 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 309784 643136 309836 643142
rect 309784 643078 309836 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 307024 590708 307076 590714
rect 307024 590650 307076 590656
rect 304264 536852 304316 536858
rect 304264 536794 304316 536800
rect 291844 324352 291896 324358
rect 291844 324294 291896 324300
rect 285678 309088 285734 309097
rect 285678 309023 285734 309032
rect 286322 309088 286378 309097
rect 286322 309023 286378 309032
rect 276662 306504 276718 306513
rect 276662 306439 276718 306448
rect 276020 266348 276072 266354
rect 276020 266290 276072 266296
rect 276020 254652 276072 254658
rect 276020 254594 276072 254600
rect 276032 253978 276060 254594
rect 276020 253972 276072 253978
rect 276020 253914 276072 253920
rect 276032 197334 276060 253914
rect 276020 197328 276072 197334
rect 276020 197270 276072 197276
rect 276676 149054 276704 306439
rect 277398 305008 277454 305017
rect 277398 304943 277454 304952
rect 276664 149048 276716 149054
rect 276664 148990 276716 148996
rect 276020 135312 276072 135318
rect 276020 135254 276072 135260
rect 274638 84144 274694 84153
rect 274638 84079 274694 84088
rect 274652 83473 274680 84079
rect 274638 83464 274694 83473
rect 274638 83399 274694 83408
rect 274640 43444 274692 43450
rect 274640 43386 274692 43392
rect 274652 16574 274680 43386
rect 274652 16546 274864 16574
rect 273904 13116 273956 13122
rect 273904 13058 273956 13064
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 16546
rect 276032 3602 276060 135254
rect 276112 95940 276164 95946
rect 276112 95882 276164 95888
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276124 3482 276152 95882
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 277136 480 277164 3538
rect 277412 3262 277440 304943
rect 282184 299532 282236 299538
rect 282184 299474 282236 299480
rect 280896 298784 280948 298790
rect 280896 298726 280948 298732
rect 280802 297392 280858 297401
rect 280802 297327 280858 297336
rect 280160 79348 280212 79354
rect 280160 79290 280212 79296
rect 277492 21412 277544 21418
rect 277492 21354 277544 21360
rect 277504 16574 277532 21354
rect 280172 16574 280200 79290
rect 280816 22778 280844 297327
rect 280908 217326 280936 298726
rect 282196 297430 282224 299474
rect 284298 297528 284354 297537
rect 284298 297463 284354 297472
rect 282092 297424 282144 297430
rect 282092 297366 282144 297372
rect 282184 297424 282236 297430
rect 282184 297366 282236 297372
rect 282104 296714 282132 297366
rect 282104 296686 282224 296714
rect 280896 217320 280948 217326
rect 280896 217262 280948 217268
rect 280804 22772 280856 22778
rect 280804 22714 280856 22720
rect 277504 16546 278360 16574
rect 280172 16546 280752 16574
rect 277400 3256 277452 3262
rect 277400 3198 277452 3204
rect 278332 480 278360 16546
rect 279516 4820 279568 4826
rect 279516 4762 279568 4768
rect 279528 480 279556 4762
rect 280724 480 280752 16546
rect 281908 4820 281960 4826
rect 281908 4762 281960 4768
rect 281920 480 281948 4762
rect 282196 3534 282224 296686
rect 282184 3528 282236 3534
rect 282184 3470 282236 3476
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 283116 480 283144 3470
rect 284312 480 284340 297463
rect 285692 267714 285720 309023
rect 289084 303748 289136 303754
rect 289084 303690 289136 303696
rect 287060 295996 287112 296002
rect 287060 295938 287112 295944
rect 285680 267708 285732 267714
rect 285680 267650 285732 267656
rect 285678 236600 285734 236609
rect 285678 236535 285734 236544
rect 284392 42084 284444 42090
rect 284392 42026 284444 42032
rect 284404 16574 284432 42026
rect 285692 16574 285720 236535
rect 284404 16546 284984 16574
rect 285692 16546 286640 16574
rect 284956 490 284984 16546
rect 285232 598 285444 626
rect 285232 490 285260 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 284956 462 285260 490
rect 285416 480 285444 598
rect 286612 480 286640 16546
rect 287072 4826 287100 295938
rect 288440 223644 288492 223650
rect 288440 223586 288492 223592
rect 287152 17264 287204 17270
rect 287152 17206 287204 17212
rect 287164 16574 287192 17206
rect 288452 16574 288480 223586
rect 289096 184210 289124 303690
rect 291856 251841 291884 324294
rect 295982 302832 296038 302841
rect 295982 302767 296038 302776
rect 291842 251832 291898 251841
rect 291842 251767 291898 251776
rect 291936 241528 291988 241534
rect 291936 241470 291988 241476
rect 291948 227050 291976 241470
rect 291844 227044 291896 227050
rect 291844 226986 291896 226992
rect 291936 227044 291988 227050
rect 291936 226986 291988 226992
rect 289084 184204 289136 184210
rect 289084 184146 289136 184152
rect 291200 60036 291252 60042
rect 291200 59978 291252 59984
rect 289084 50380 289136 50386
rect 289084 50322 289136 50328
rect 287164 16546 287376 16574
rect 288452 16546 289032 16574
rect 287060 4820 287112 4826
rect 287060 4762 287112 4768
rect 287348 490 287376 16546
rect 287624 598 287836 626
rect 287624 490 287652 598
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287348 462 287652 490
rect 287808 480 287836 598
rect 289004 480 289032 16546
rect 289096 3398 289124 50322
rect 291212 16574 291240 59978
rect 291212 16546 291424 16574
rect 289084 3392 289136 3398
rect 289084 3334 289136 3340
rect 290186 3360 290242 3369
rect 290186 3295 290242 3304
rect 290200 480 290228 3295
rect 291396 480 291424 16546
rect 291856 3534 291884 226986
rect 295338 141400 295394 141409
rect 295338 141335 295394 141344
rect 292672 22772 292724 22778
rect 292672 22714 292724 22720
rect 292684 16574 292712 22714
rect 295352 16574 295380 141335
rect 295996 22778 296024 302767
rect 298744 298172 298796 298178
rect 298744 298114 298796 298120
rect 298756 254658 298784 298114
rect 299478 294536 299534 294545
rect 299478 294471 299534 294480
rect 298744 254652 298796 254658
rect 298744 254594 298796 254600
rect 298100 233300 298152 233306
rect 298100 233242 298152 233248
rect 295984 22772 296036 22778
rect 295984 22714 296036 22720
rect 292684 16546 293264 16574
rect 295352 16546 295656 16574
rect 291844 3528 291896 3534
rect 291844 3470 291896 3476
rect 292580 3528 292632 3534
rect 292580 3470 292632 3476
rect 292592 480 292620 3470
rect 293236 490 293264 16546
rect 294880 3392 294932 3398
rect 294880 3334 294932 3340
rect 293512 598 293724 626
rect 293512 490 293540 598
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 462 293540 490
rect 293696 480 293724 598
rect 294892 480 294920 3334
rect 295628 490 295656 16546
rect 297272 3528 297324 3534
rect 297272 3470 297324 3476
rect 295904 598 296116 626
rect 295904 490 295932 598
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 462 295932 490
rect 296088 480 296116 598
rect 297284 480 297312 3470
rect 298112 490 298140 233242
rect 299492 3534 299520 294471
rect 302240 261520 302292 261526
rect 302240 261462 302292 261468
rect 300860 184204 300912 184210
rect 300860 184146 300912 184152
rect 300872 16574 300900 184146
rect 300872 16546 301544 16574
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 299664 3188 299716 3194
rect 299664 3130 299716 3136
rect 298296 598 298508 626
rect 298296 490 298324 598
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 462 298324 490
rect 298480 480 298508 598
rect 299676 480 299704 3130
rect 300768 2100 300820 2106
rect 300768 2042 300820 2048
rect 300780 480 300808 2042
rect 301516 490 301544 16546
rect 302252 3194 302280 261462
rect 304276 258058 304304 536794
rect 305642 307864 305698 307873
rect 305642 307799 305698 307808
rect 304264 258052 304316 258058
rect 304264 257994 304316 258000
rect 304264 243024 304316 243030
rect 304264 242966 304316 242972
rect 303620 217320 303672 217326
rect 303620 217262 303672 217268
rect 302332 44872 302384 44878
rect 302332 44814 302384 44820
rect 302344 16574 302372 44814
rect 303632 16574 303660 217262
rect 304276 60722 304304 242966
rect 304264 60716 304316 60722
rect 304264 60658 304316 60664
rect 304264 57248 304316 57254
rect 304264 57190 304316 57196
rect 302344 16546 302832 16574
rect 303632 16546 303936 16574
rect 302240 3188 302292 3194
rect 302240 3130 302292 3136
rect 302804 2938 302832 16546
rect 302884 11756 302936 11762
rect 302884 11698 302936 11704
rect 302896 3126 302924 11698
rect 302884 3120 302936 3126
rect 302884 3062 302936 3068
rect 302804 2910 303200 2938
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 2910
rect 303908 490 303936 16546
rect 304276 4010 304304 57190
rect 305656 6186 305684 307799
rect 307036 258806 307064 590650
rect 309796 260137 309824 643078
rect 582470 630864 582526 630873
rect 582470 630799 582526 630808
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 511320 580226 511329
rect 580170 511255 580172 511264
rect 580224 511255 580226 511264
rect 580172 511226 580224 511232
rect 582378 458144 582434 458153
rect 582378 458079 582434 458088
rect 582392 436762 582420 458079
rect 582380 436756 582432 436762
rect 582380 436698 582432 436704
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 321558 307048 321614 307057
rect 321558 306983 321614 306992
rect 317420 297424 317472 297430
rect 317420 297366 317472 297372
rect 309782 260128 309838 260137
rect 309782 260063 309838 260072
rect 307024 258800 307076 258806
rect 307024 258742 307076 258748
rect 313924 245744 313976 245750
rect 313924 245686 313976 245692
rect 306380 222216 306432 222222
rect 306380 222158 306432 222164
rect 305644 6180 305696 6186
rect 305644 6122 305696 6128
rect 304264 4004 304316 4010
rect 304264 3946 304316 3952
rect 305552 3120 305604 3126
rect 305552 3062 305604 3068
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 3062
rect 306392 490 306420 222158
rect 309784 221468 309836 221474
rect 309784 221410 309836 221416
rect 307852 40724 307904 40730
rect 307852 40666 307904 40672
rect 307864 16250 307892 40666
rect 307852 16244 307904 16250
rect 307852 16186 307904 16192
rect 309048 16244 309100 16250
rect 309048 16186 309100 16192
rect 307944 4004 307996 4010
rect 307944 3946 307996 3952
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3946
rect 309060 480 309088 16186
rect 309796 3534 309824 221410
rect 313936 193186 313964 245686
rect 313924 193180 313976 193186
rect 313924 193122 313976 193128
rect 316040 156664 316092 156670
rect 316040 156606 316092 156612
rect 313280 149116 313332 149122
rect 313280 149058 313332 149064
rect 311900 62824 311952 62830
rect 311900 62766 311952 62772
rect 311912 16574 311940 62766
rect 311912 16546 312216 16574
rect 311440 6180 311492 6186
rect 311440 6122 311492 6128
rect 310244 5568 310296 5574
rect 310244 5510 310296 5516
rect 309784 3528 309836 3534
rect 309784 3470 309836 3476
rect 310256 480 310284 5510
rect 311452 480 311480 6122
rect 312188 490 312216 16546
rect 313292 5574 313320 149058
rect 316052 16574 316080 156606
rect 317432 16574 317460 297366
rect 318798 124808 318854 124817
rect 318798 124743 318854 124752
rect 318812 16574 318840 124743
rect 320178 83464 320234 83473
rect 320178 83399 320234 83408
rect 320192 16574 320220 83399
rect 321572 16574 321600 306983
rect 336004 303680 336056 303686
rect 336004 303622 336056 303628
rect 327078 302288 327134 302297
rect 327078 302223 327134 302232
rect 324962 300520 325018 300529
rect 324962 300455 325018 300464
rect 322204 46232 322256 46238
rect 322204 46174 322256 46180
rect 316052 16546 316264 16574
rect 317432 16546 318104 16574
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 313280 5568 313332 5574
rect 313280 5510 313332 5516
rect 313832 3528 313884 3534
rect 313832 3470 313884 3476
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 3470
rect 315028 3460 315080 3466
rect 315028 3402 315080 3408
rect 315040 480 315068 3402
rect 316236 480 316264 16546
rect 317328 7608 317380 7614
rect 317328 7550 317380 7556
rect 317340 480 317368 7550
rect 318076 490 318104 16546
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 16546
rect 320468 490 320496 16546
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 322216 3534 322244 46174
rect 322940 15904 322992 15910
rect 322940 15846 322992 15852
rect 322204 3528 322256 3534
rect 322204 3470 322256 3476
rect 322952 490 322980 15846
rect 324872 13116 324924 13122
rect 324872 13058 324924 13064
rect 324412 3528 324464 3534
rect 324412 3470 324464 3476
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 3470
rect 324884 3210 324912 13058
rect 324976 3369 325004 300455
rect 325700 19984 325752 19990
rect 325700 19926 325752 19932
rect 325712 16574 325740 19926
rect 325712 16546 326384 16574
rect 324962 3360 325018 3369
rect 324962 3295 325018 3304
rect 324884 3182 325648 3210
rect 325620 480 325648 3182
rect 326356 490 326384 16546
rect 327092 3466 327120 302223
rect 333978 289096 334034 289105
rect 333978 289031 334034 289040
rect 331220 219496 331272 219502
rect 331220 219438 331272 219444
rect 327172 82136 327224 82142
rect 327172 82078 327224 82084
rect 327184 16574 327212 82078
rect 327184 16546 328040 16574
rect 327080 3460 327132 3466
rect 327080 3402 327132 3408
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 16546
rect 331232 3534 331260 219438
rect 332600 66904 332652 66910
rect 332600 66846 332652 66852
rect 331312 18624 331364 18630
rect 331312 18566 331364 18572
rect 331324 16574 331352 18566
rect 331324 16546 331628 16574
rect 329196 3528 329248 3534
rect 329196 3470 329248 3476
rect 331220 3528 331272 3534
rect 331220 3470 331272 3476
rect 329208 480 329236 3470
rect 330392 3460 330444 3466
rect 330392 3402 330444 3408
rect 330404 480 330432 3402
rect 331600 480 331628 16546
rect 332612 3534 332640 66846
rect 333992 11014 334020 289031
rect 335360 22772 335412 22778
rect 335360 22714 335412 22720
rect 335372 16574 335400 22714
rect 335372 16546 335952 16574
rect 333980 11008 334032 11014
rect 333980 10950 334032 10956
rect 334624 11008 334676 11014
rect 334624 10950 334676 10956
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 332690 3360 332746 3369
rect 332690 3295 332746 3304
rect 332704 480 332732 3295
rect 333900 480 333928 3470
rect 334636 490 334664 10950
rect 335924 3210 335952 16546
rect 336016 3369 336044 303622
rect 345018 301744 345074 301753
rect 345018 301679 345074 301688
rect 342258 284880 342314 284889
rect 342258 284815 342314 284824
rect 339498 283520 339554 283529
rect 339498 283455 339554 283464
rect 338120 215960 338172 215966
rect 338120 215902 338172 215908
rect 337016 14476 337068 14482
rect 337016 14418 337068 14424
rect 336002 3360 336058 3369
rect 336002 3295 336058 3304
rect 335924 3182 336320 3210
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3182
rect 337028 490 337056 14418
rect 338132 3466 338160 215902
rect 338212 84856 338264 84862
rect 338212 84798 338264 84804
rect 338224 16574 338252 84798
rect 338224 16546 338712 16574
rect 338120 3460 338172 3466
rect 338120 3402 338172 3408
rect 337304 598 337516 626
rect 337304 490 337332 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 462 337332 490
rect 337488 480 337516 598
rect 338684 480 338712 16546
rect 339512 490 339540 283455
rect 341524 247104 341576 247110
rect 341524 247046 341576 247052
rect 341536 179382 341564 247046
rect 341524 179376 341576 179382
rect 341524 179318 341576 179324
rect 340880 77988 340932 77994
rect 340880 77930 340932 77936
rect 340892 16574 340920 77930
rect 342272 16574 342300 284815
rect 343640 69692 343692 69698
rect 343640 69634 343692 69640
rect 343652 16574 343680 69634
rect 340892 16546 341012 16574
rect 342272 16546 342944 16574
rect 343652 16546 344600 16574
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 16546
rect 342168 3732 342220 3738
rect 342168 3674 342220 3680
rect 342180 480 342208 3674
rect 342916 490 342944 16546
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 16546
rect 345032 3738 345060 301679
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580276 262886 580304 365055
rect 582378 312080 582434 312089
rect 582378 312015 582434 312024
rect 580264 262880 580316 262886
rect 580264 262822 580316 262828
rect 582392 251870 582420 312015
rect 582484 273970 582512 630799
rect 582562 617536 582618 617545
rect 582562 617471 582618 617480
rect 582576 585818 582604 617471
rect 582564 585812 582616 585818
rect 582564 585754 582616 585760
rect 582562 577688 582618 577697
rect 582562 577623 582618 577632
rect 582472 273964 582524 273970
rect 582472 273906 582524 273912
rect 582576 267073 582604 577623
rect 582668 570654 582696 683839
rect 582746 582448 582802 582457
rect 582746 582383 582802 582392
rect 582656 570648 582708 570654
rect 582656 570590 582708 570596
rect 582760 564369 582788 582383
rect 582746 564360 582802 564369
rect 582746 564295 582802 564304
rect 582654 524512 582710 524521
rect 582654 524447 582710 524456
rect 582562 267064 582618 267073
rect 582562 266999 582618 267008
rect 582668 264217 582696 524447
rect 582746 484664 582802 484673
rect 582746 484599 582802 484608
rect 582654 264208 582710 264217
rect 582654 264143 582710 264152
rect 582760 260166 582788 484599
rect 582838 471472 582894 471481
rect 582838 471407 582894 471416
rect 582748 260160 582800 260166
rect 582748 260102 582800 260108
rect 582470 258904 582526 258913
rect 582470 258839 582526 258848
rect 582380 251864 582432 251870
rect 582380 251806 582432 251812
rect 582484 250510 582512 258839
rect 582852 256698 582880 471407
rect 583114 431624 583170 431633
rect 583114 431559 583170 431568
rect 582930 293176 582986 293185
rect 582930 293111 582986 293120
rect 582840 256692 582892 256698
rect 582840 256634 582892 256640
rect 582472 250504 582524 250510
rect 582472 250446 582524 250452
rect 582380 249824 582432 249830
rect 582380 249766 582432 249772
rect 582392 245585 582420 249766
rect 582564 248464 582616 248470
rect 582564 248406 582616 248412
rect 582472 247716 582524 247722
rect 582472 247658 582524 247664
rect 582378 245576 582434 245585
rect 582378 245511 582434 245520
rect 582484 245426 582512 247658
rect 582392 245398 582512 245426
rect 349804 244384 349856 244390
rect 349804 244326 349856 244332
rect 349816 139398 349844 244326
rect 580264 240780 580316 240786
rect 580264 240722 580316 240728
rect 351920 225004 351972 225010
rect 351920 224946 351972 224952
rect 349804 139392 349856 139398
rect 349804 139334 349856 139340
rect 349160 80708 349212 80714
rect 349160 80650 349212 80656
rect 346952 8968 347004 8974
rect 346952 8910 347004 8916
rect 345020 3732 345072 3738
rect 345020 3674 345072 3680
rect 345756 3392 345808 3398
rect 345756 3334 345808 3340
rect 345768 480 345796 3334
rect 346964 480 346992 8910
rect 349172 6914 349200 80650
rect 349080 6886 349200 6914
rect 348054 4040 348110 4049
rect 348054 3975 348110 3984
rect 348068 480 348096 3975
rect 349080 3482 349108 6886
rect 349080 3454 349292 3482
rect 349264 480 349292 3454
rect 351644 3460 351696 3466
rect 351644 3402 351696 3408
rect 350446 3360 350502 3369
rect 350446 3295 350502 3304
rect 350460 480 350488 3295
rect 351656 480 351684 3402
rect 351932 3398 351960 224946
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 356060 122120 356112 122126
rect 356060 122062 356112 122068
rect 356072 4049 356100 122062
rect 357438 86184 357494 86193
rect 357438 86119 357494 86128
rect 356058 4040 356114 4049
rect 356058 3975 356114 3984
rect 357452 3466 357480 86119
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580276 33153 580304 240722
rect 580356 238808 580408 238814
rect 580356 238750 580408 238756
rect 580368 165889 580396 238750
rect 582392 232393 582420 245398
rect 582576 238754 582604 248406
rect 582748 242208 582800 242214
rect 582748 242150 582800 242156
rect 582484 238726 582604 238754
rect 582378 232384 582434 232393
rect 582378 232319 582434 232328
rect 582380 227044 582432 227050
rect 582380 226986 582432 226992
rect 580354 165880 580410 165889
rect 580354 165815 580410 165824
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 582392 6633 582420 226986
rect 582484 205737 582512 238726
rect 582654 234696 582710 234705
rect 582654 234631 582710 234640
rect 582564 231872 582616 231878
rect 582564 231814 582616 231820
rect 582470 205728 582526 205737
rect 582470 205663 582526 205672
rect 582576 19825 582604 231814
rect 582668 46345 582696 234631
rect 582760 73001 582788 242150
rect 582838 237960 582894 237969
rect 582838 237895 582894 237904
rect 582852 86193 582880 237895
rect 582838 86184 582894 86193
rect 582838 86119 582894 86128
rect 582746 72992 582802 73001
rect 582746 72927 582802 72936
rect 582654 46336 582710 46345
rect 582654 46271 582710 46280
rect 582562 19816 582618 19825
rect 582562 19751 582618 19760
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 582944 3534 582972 293111
rect 583022 279440 583078 279449
rect 583022 279375 583078 279384
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 582932 3528 582984 3534
rect 582932 3470 582984 3476
rect 357440 3460 357492 3466
rect 357440 3402 357492 3408
rect 351920 3392 351972 3398
rect 351920 3334 351972 3340
rect 581000 2916 581052 2922
rect 581000 2858 581052 2864
rect 581012 480 581040 2858
rect 582208 480 582236 3470
rect 583036 2922 583064 279375
rect 583128 254590 583156 431559
rect 583206 418296 583262 418305
rect 583206 418231 583262 418240
rect 583220 265674 583248 418231
rect 583298 404968 583354 404977
rect 583298 404903 583354 404912
rect 583208 265668 583260 265674
rect 583208 265610 583260 265616
rect 583312 258738 583340 404903
rect 583390 378448 583446 378457
rect 583390 378383 583446 378392
rect 583300 258732 583352 258738
rect 583300 258674 583352 258680
rect 583116 254584 583168 254590
rect 583116 254526 583168 254532
rect 583404 253230 583432 378383
rect 583482 351656 583538 351665
rect 583482 351591 583538 351600
rect 583496 257378 583524 351591
rect 583588 271153 583616 696895
rect 583574 271144 583630 271153
rect 583574 271079 583630 271088
rect 583484 257372 583536 257378
rect 583484 257314 583536 257320
rect 583392 253224 583444 253230
rect 583392 253166 583444 253172
rect 583300 245676 583352 245682
rect 583300 245618 583352 245624
rect 583116 242956 583168 242962
rect 583116 242898 583168 242904
rect 583128 112849 583156 242898
rect 583208 228404 583260 228410
rect 583208 228346 583260 228352
rect 583114 112840 583170 112849
rect 583114 112775 583170 112784
rect 583220 99521 583248 228346
rect 583312 126041 583340 245618
rect 583392 244316 583444 244322
rect 583392 244258 583444 244264
rect 583404 152697 583432 244258
rect 583482 213208 583538 213217
rect 583482 213143 583538 213152
rect 583390 152688 583446 152697
rect 583390 152623 583446 152632
rect 583298 126032 583354 126041
rect 583298 125967 583354 125976
rect 583206 99512 583262 99521
rect 583206 99447 583262 99456
rect 583496 6914 583524 213143
rect 583404 6886 583524 6914
rect 583024 2916 583076 2922
rect 583024 2858 583076 2864
rect 583404 480 583432 6886
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 2778 671200 2834 671256
rect 3422 658144 3478 658200
rect 3422 632032 3478 632088
rect 3330 579944 3386 580000
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3514 566888 3570 566944
rect 3422 553832 3478 553888
rect 4802 541048 4858 541104
rect 3514 527876 3570 527912
rect 3514 527856 3516 527876
rect 3516 527856 3568 527876
rect 3568 527856 3570 527876
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 3422 501744 3478 501800
rect 2962 475668 2964 475688
rect 2964 475668 3016 475688
rect 3016 475668 3018 475688
rect 2962 475632 3018 475668
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 2778 423580 2780 423600
rect 2780 423580 2832 423600
rect 2832 423580 2834 423600
rect 2778 423544 2834 423580
rect 2870 410488 2926 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 4066 392128 4122 392184
rect 17222 397432 17278 397488
rect 7562 391856 7618 391912
rect 3422 371320 3478 371376
rect 3330 358400 3386 358456
rect 3330 345344 3386 345400
rect 3882 319252 3938 319288
rect 3882 319232 3884 319252
rect 3884 319232 3936 319252
rect 3936 319232 3938 319252
rect 3422 306176 3478 306232
rect 3514 293120 3570 293176
rect 3054 267144 3110 267200
rect 29642 388728 29698 388784
rect 17222 314744 17278 314800
rect 16486 310528 16542 310584
rect 3422 254088 3478 254144
rect 2778 241032 2834 241088
rect 15106 235184 15162 235240
rect 4066 222808 4122 222864
rect 3146 214920 3202 214976
rect 3238 201864 3294 201920
rect 2778 188844 2780 188864
rect 2780 188844 2832 188864
rect 2832 188844 2834 188864
rect 2778 188808 2834 188844
rect 3422 162832 3478 162888
rect 2962 149776 3018 149832
rect 3238 136720 3294 136776
rect 3146 110608 3202 110664
rect 3054 97552 3110 97608
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3422 58520 3478 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 5446 188264 5502 188320
rect 6826 39208 6882 39264
rect 16394 151000 16450 151056
rect 8758 3304 8814 3360
rect 16486 3984 16542 4040
rect 22742 311888 22798 311944
rect 18602 310664 18658 310720
rect 18234 3984 18290 4040
rect 17222 3304 17278 3360
rect 22006 298696 22062 298752
rect 21362 185544 21418 185600
rect 29642 309168 29698 309224
rect 26146 306448 26202 306504
rect 23386 33768 23442 33824
rect 27526 21256 27582 21312
rect 32954 275168 33010 275224
rect 34426 313248 34482 313304
rect 34242 261432 34298 261488
rect 33046 232464 33102 232520
rect 37094 531936 37150 531992
rect 35806 316104 35862 316160
rect 38566 214512 38622 214568
rect 31298 3304 31354 3360
rect 41234 406952 41290 407008
rect 41050 267824 41106 267880
rect 40682 153720 40738 153776
rect 43810 338680 43866 338736
rect 42614 216552 42670 216608
rect 43994 384240 44050 384296
rect 43902 321544 43958 321600
rect 44086 284824 44142 284880
rect 43994 239808 44050 239864
rect 42706 35128 42762 35184
rect 41326 22616 41382 22672
rect 45282 234504 45338 234560
rect 45466 267824 45522 267880
rect 49606 393488 49662 393544
rect 48226 264968 48282 265024
rect 48042 244432 48098 244488
rect 47950 237360 48006 237416
rect 48226 238584 48282 238640
rect 48226 237360 48282 237416
rect 49514 254496 49570 254552
rect 49422 223488 49478 223544
rect 48042 216552 48098 216608
rect 50710 285776 50766 285832
rect 49606 223488 49662 223544
rect 49514 209616 49570 209672
rect 48226 146920 48282 146976
rect 45466 36488 45522 36544
rect 53746 578856 53802 578912
rect 52182 436192 52238 436248
rect 50894 389136 50950 389192
rect 50894 387640 50950 387696
rect 53562 433608 53618 433664
rect 52182 306312 52238 306368
rect 52182 304952 52238 305008
rect 50710 220768 50766 220824
rect 50342 149640 50398 149696
rect 52090 228928 52146 228984
rect 52458 276120 52514 276176
rect 52182 224848 52238 224904
rect 52458 247152 52514 247208
rect 52090 137264 52146 137320
rect 50986 90752 51042 90808
rect 53746 420144 53802 420200
rect 53562 282104 53618 282160
rect 53470 271904 53526 271960
rect 53562 247152 53618 247208
rect 54850 264152 54906 264208
rect 55126 387912 55182 387968
rect 55126 386416 55182 386472
rect 55218 248376 55274 248432
rect 59266 581032 59322 581088
rect 56598 406952 56654 407008
rect 56414 264152 56470 264208
rect 58990 533296 59046 533352
rect 57702 331200 57758 331256
rect 57518 275848 57574 275904
rect 57518 275168 57574 275224
rect 56506 248376 56562 248432
rect 54482 91704 54538 91760
rect 53746 24112 53802 24168
rect 57702 246200 57758 246256
rect 57610 222128 57666 222184
rect 57702 205536 57758 205592
rect 58990 393488 59046 393544
rect 60462 283464 60518 283520
rect 59082 237224 59138 237280
rect 57702 90888 57758 90944
rect 58622 88984 58678 89040
rect 57886 86264 57942 86320
rect 54482 3304 54538 3360
rect 60370 253952 60426 254008
rect 61934 418240 61990 418296
rect 61842 318008 61898 318064
rect 60554 273264 60610 273320
rect 60554 269184 60610 269240
rect 60462 226208 60518 226264
rect 62026 389272 62082 389328
rect 61934 295296 61990 295352
rect 61842 284824 61898 284880
rect 61750 270680 61806 270736
rect 58990 88168 59046 88224
rect 61934 263608 61990 263664
rect 61842 252728 61898 252784
rect 63130 287272 63186 287328
rect 62854 273128 62910 273184
rect 66074 567568 66130 567624
rect 66534 579944 66590 580000
rect 66902 578584 66958 578640
rect 66442 575864 66498 575920
rect 66626 573144 66682 573200
rect 66718 571784 66774 571840
rect 66810 564712 66866 564768
rect 66534 564168 66590 564224
rect 66810 561992 66866 562048
rect 66810 560632 66866 560688
rect 66810 559272 66866 559328
rect 66810 557912 66866 557968
rect 66718 555192 66774 555248
rect 66810 553560 66866 553616
rect 66810 549480 66866 549536
rect 66534 546760 66590 546816
rect 66258 545944 66314 546000
rect 66350 544448 66406 544504
rect 66626 543088 66682 543144
rect 64786 411304 64842 411360
rect 63406 263472 63462 263528
rect 63314 251232 63370 251288
rect 63314 135904 63370 135960
rect 63130 120128 63186 120184
rect 64142 240760 64198 240816
rect 65890 401512 65946 401568
rect 66626 539960 66682 540016
rect 66074 433880 66130 433936
rect 65890 334056 65946 334112
rect 65890 294072 65946 294128
rect 64786 252728 64842 252784
rect 64602 113192 64658 113248
rect 64878 249872 64934 249928
rect 64786 241576 64842 241632
rect 66350 433336 66406 433392
rect 66810 432520 66866 432576
rect 66810 431432 66866 431488
rect 66810 430344 66866 430400
rect 66258 429276 66314 429312
rect 66258 429256 66260 429276
rect 66260 429256 66312 429276
rect 66312 429256 66314 429276
rect 66166 428168 66222 428224
rect 65982 240080 66038 240136
rect 66810 427352 66866 427408
rect 66534 425176 66590 425232
rect 66626 424088 66682 424144
rect 66810 423272 66866 423328
rect 66810 421096 66866 421152
rect 66810 420008 66866 420064
rect 66810 417016 66866 417072
rect 66718 415928 66774 415984
rect 66718 414840 66774 414896
rect 66258 412936 66314 412992
rect 66810 410760 66866 410816
rect 66626 408856 66682 408912
rect 66810 407768 66866 407824
rect 66442 405592 66498 405648
rect 66350 402600 66406 402656
rect 66810 404504 66866 404560
rect 67546 577224 67602 577280
rect 66994 570152 67050 570208
rect 67454 552200 67510 552256
rect 67454 433236 67456 433256
rect 67456 433236 67508 433256
rect 67508 433236 67510 433256
rect 67454 433200 67510 433236
rect 66994 418140 66996 418160
rect 66996 418140 67048 418160
rect 67048 418140 67050 418160
rect 66994 418104 67050 418140
rect 67454 409672 67510 409728
rect 66810 403688 66866 403744
rect 66810 400424 66866 400480
rect 66810 399608 66866 399664
rect 66810 398520 66866 398576
rect 66902 397432 66958 397488
rect 66810 396344 66866 396400
rect 66810 395292 66812 395312
rect 66812 395292 66864 395312
rect 66864 395292 66866 395312
rect 66810 395256 66866 395292
rect 66810 394440 66866 394496
rect 66810 392264 66866 392320
rect 66810 391176 66866 391232
rect 66810 387504 66866 387560
rect 72422 585112 72478 585168
rect 71778 584840 71834 584896
rect 69478 582392 69534 582448
rect 70214 582392 70270 582448
rect 79966 587968 80022 588024
rect 75366 581032 75422 581088
rect 79046 582664 79102 582720
rect 78126 581032 78182 581088
rect 82726 583752 82782 583808
rect 83002 581168 83058 581224
rect 70950 580760 71006 580816
rect 84198 580760 84254 580816
rect 89718 582664 89774 582720
rect 88246 582528 88302 582584
rect 89718 581576 89774 581632
rect 92110 582392 92166 582448
rect 88706 580760 88762 580816
rect 68650 578856 68706 578912
rect 67730 575320 67786 575376
rect 67730 568792 67786 568848
rect 67638 566616 67694 566672
rect 67638 556552 67694 556608
rect 67822 550840 67878 550896
rect 69110 539824 69166 539880
rect 68466 436192 68522 436248
rect 93858 539844 93914 539880
rect 93858 539824 93860 539844
rect 93860 539824 93912 539844
rect 93912 539824 93914 539844
rect 76470 536696 76526 536752
rect 76470 535608 76526 535664
rect 75918 535472 75974 535528
rect 77206 535608 77262 535664
rect 76746 535472 76802 535528
rect 75458 434424 75514 434480
rect 74722 434288 74778 434344
rect 76194 434288 76250 434344
rect 77390 436192 77446 436248
rect 77482 435376 77538 435432
rect 81346 520920 81402 520976
rect 80058 453192 80114 453248
rect 77942 434696 77998 434752
rect 80242 434288 80298 434344
rect 81346 444896 81402 444952
rect 80426 434832 80482 434888
rect 80978 434288 81034 434344
rect 83462 443536 83518 443592
rect 86222 449112 86278 449168
rect 83186 436056 83242 436112
rect 82910 434696 82966 434752
rect 81898 434288 81954 434344
rect 67730 414044 67786 414080
rect 67730 414024 67732 414044
rect 67732 414024 67784 414044
rect 67784 414024 67786 414044
rect 67546 405592 67602 405648
rect 67546 326304 67602 326360
rect 67546 281288 67602 281344
rect 66626 279656 66682 279712
rect 66810 278840 66866 278896
rect 66810 278044 66866 278080
rect 66810 278024 66812 278044
rect 66812 278024 66864 278044
rect 66864 278024 66866 278044
rect 66810 276392 66866 276448
rect 66902 275576 66958 275632
rect 66534 273944 66590 274000
rect 66258 273128 66314 273184
rect 66810 272312 66866 272368
rect 66258 271904 66314 271960
rect 66166 271496 66222 271552
rect 66166 270680 66222 270736
rect 66810 270680 66866 270736
rect 66166 268232 66222 268288
rect 65982 128968 66038 129024
rect 65522 123800 65578 123856
rect 66810 267416 66866 267472
rect 66258 266464 66314 266520
rect 66810 264968 66866 265024
rect 66626 263336 66682 263392
rect 66902 262520 66958 262576
rect 66718 260888 66774 260944
rect 66442 260072 66498 260128
rect 66626 257624 66682 257680
rect 66350 256808 66406 256864
rect 66810 255992 66866 256048
rect 66810 255176 66866 255232
rect 66994 253544 67050 253600
rect 66810 251096 66866 251152
rect 66718 249464 66774 249520
rect 66994 246200 67050 246256
rect 66902 244568 66958 244624
rect 66810 243752 66866 243808
rect 67454 247052 67456 247072
rect 67456 247052 67508 247072
rect 67508 247052 67510 247072
rect 67454 247016 67510 247052
rect 66166 145560 66222 145616
rect 66074 125976 66130 126032
rect 66074 119176 66130 119232
rect 66258 134408 66314 134464
rect 66258 133592 66314 133648
rect 66258 131960 66314 132016
rect 66350 131144 66406 131200
rect 66442 128152 66498 128208
rect 66718 126792 66774 126848
rect 66258 124344 66314 124400
rect 66718 120536 66774 120592
rect 66258 119176 66314 119232
rect 66166 117544 66222 117600
rect 66626 113192 66682 113248
rect 66258 110200 66314 110256
rect 66718 106392 66774 106448
rect 66258 104796 66260 104816
rect 66260 104796 66312 104816
rect 66312 104796 66314 104816
rect 66258 104760 66314 104796
rect 66902 127608 66958 127664
rect 66902 125160 66958 125216
rect 66902 122984 66958 123040
rect 66902 122168 66958 122224
rect 66902 120028 66904 120048
rect 66904 120028 66956 120048
rect 66956 120028 66958 120048
rect 66902 119992 66958 120028
rect 66902 118360 66958 118416
rect 66902 117000 66958 117056
rect 66902 115368 66958 115424
rect 67178 114588 67180 114608
rect 67180 114588 67232 114608
rect 67232 114588 67234 114608
rect 67178 114552 67234 114588
rect 66902 112376 66958 112432
rect 66902 110744 66958 110800
rect 66902 109384 66958 109440
rect 66902 108568 66958 108624
rect 66994 107752 67050 107808
rect 66902 106936 66958 106992
rect 66902 105576 66958 105632
rect 66902 103128 66958 103184
rect 66810 101768 66866 101824
rect 66442 100952 66498 101008
rect 66810 100136 66866 100192
rect 66810 99592 66866 99648
rect 66810 98776 66866 98832
rect 66258 96328 66314 96384
rect 66902 97144 66958 97200
rect 66810 95784 66866 95840
rect 66442 94968 66498 95024
rect 66810 93336 66866 93392
rect 67362 103944 67418 104000
rect 85762 437552 85818 437608
rect 84474 434560 84530 434616
rect 83738 434424 83794 434480
rect 86866 437552 86922 437608
rect 88430 462984 88486 463040
rect 90454 468424 90510 468480
rect 88338 440952 88394 441008
rect 87326 436056 87382 436112
rect 88246 436056 88302 436112
rect 85854 434288 85910 434344
rect 87142 434288 87198 434344
rect 95330 575320 95386 575376
rect 95238 563624 95294 563680
rect 94778 555464 94834 555520
rect 94686 538192 94742 538248
rect 94778 518064 94834 518120
rect 91098 436192 91154 436248
rect 95422 567160 95478 567216
rect 97538 577496 97594 577552
rect 97906 576716 97908 576736
rect 97908 576716 97960 576736
rect 97960 576716 97962 576736
rect 97906 576680 97962 576716
rect 97630 575320 97686 575376
rect 97446 573416 97502 573472
rect 97078 571396 97134 571432
rect 97078 571376 97080 571396
rect 97080 571376 97132 571396
rect 97132 571376 97134 571396
rect 97906 570288 97962 570344
rect 96802 569064 96858 569120
rect 97906 569064 97962 569120
rect 97906 565800 97962 565856
rect 96802 562264 96858 562320
rect 96894 560904 96950 560960
rect 96802 559544 96858 559600
rect 96710 558728 96766 558784
rect 96802 556824 96858 556880
rect 95514 552472 95570 552528
rect 96618 552472 96674 552528
rect 96710 542952 96766 543008
rect 96618 538872 96674 538928
rect 95422 527720 95478 527776
rect 97170 558748 97226 558784
rect 97170 558728 97172 558748
rect 97172 558728 97224 558748
rect 97224 558728 97226 558748
rect 96986 552744 97042 552800
rect 97906 550704 97962 550760
rect 97078 549364 97134 549400
rect 97078 549344 97080 549364
rect 97080 549344 97132 549364
rect 97132 549344 97134 549364
rect 96986 545672 97042 545728
rect 97354 544312 97410 544368
rect 96986 461488 97042 461544
rect 95238 454688 95294 454744
rect 96618 444216 96674 444272
rect 96618 442992 96674 443048
rect 92662 434696 92718 434752
rect 94226 434288 94282 434344
rect 101402 585112 101458 585168
rect 99286 572600 99342 572656
rect 100022 547848 100078 547904
rect 98642 439456 98698 439512
rect 100114 507864 100170 507920
rect 104162 582528 104218 582584
rect 102782 581576 102838 581632
rect 101402 446392 101458 446448
rect 100022 434968 100078 435024
rect 101218 434832 101274 434888
rect 97170 434288 97226 434344
rect 102598 434288 102654 434344
rect 106922 458768 106978 458824
rect 104162 435240 104218 435296
rect 104162 434288 104218 434344
rect 106738 436328 106794 436384
rect 107658 436056 107714 436112
rect 109130 436192 109186 436248
rect 108210 436056 108266 436112
rect 108210 434288 108266 434344
rect 71226 433880 71282 433936
rect 100574 433880 100630 433936
rect 110418 436056 110474 436112
rect 110970 436056 111026 436112
rect 109590 433880 109646 433936
rect 70858 433744 70914 433800
rect 87970 433744 88026 433800
rect 98458 433744 98514 433800
rect 73434 433608 73490 433664
rect 78402 433608 78458 433664
rect 79598 433608 79654 433664
rect 87326 433608 87382 433664
rect 89994 433608 90050 433664
rect 91466 433608 91522 433664
rect 93490 433608 93546 433664
rect 95146 433608 95202 433664
rect 98366 433608 98422 433664
rect 99838 433608 99894 433664
rect 105174 433608 105230 433664
rect 110418 433608 110474 433664
rect 111706 433608 111762 433664
rect 70306 385056 70362 385112
rect 69662 338000 69718 338056
rect 69110 314880 69166 314936
rect 69018 284824 69074 284880
rect 70306 314880 70362 314936
rect 68282 277364 68338 277400
rect 68282 277344 68284 277364
rect 68284 277344 68336 277364
rect 68336 277344 68338 277364
rect 68190 258712 68246 258768
rect 67638 241304 67694 241360
rect 67546 129784 67602 129840
rect 67546 102584 67602 102640
rect 67546 102176 67602 102232
rect 67454 97960 67510 98016
rect 63222 3304 63278 3360
rect 68558 241732 68614 241768
rect 68558 241712 68560 241732
rect 68560 241712 68612 241732
rect 68612 241712 68614 241732
rect 68374 241440 68430 241496
rect 72422 390360 72478 390416
rect 71870 389000 71926 389056
rect 72974 384376 73030 384432
rect 71686 380840 71742 380896
rect 70490 328480 70546 328536
rect 72422 319368 72478 319424
rect 71686 318008 71742 318064
rect 70398 288360 70454 288416
rect 72606 318824 72662 318880
rect 72974 318844 73030 318880
rect 72974 318824 72976 318844
rect 72976 318824 73028 318844
rect 73028 318824 73030 318844
rect 71180 283736 71236 283792
rect 71042 283192 71098 283248
rect 71870 283464 71926 283520
rect 73802 343712 73858 343768
rect 73250 300192 73306 300248
rect 73802 300192 73858 300248
rect 73802 287680 73858 287736
rect 74078 285776 74134 285832
rect 73526 283464 73582 283520
rect 75826 386280 75882 386336
rect 75182 379480 75238 379536
rect 75274 340892 75276 340912
rect 75276 340892 75328 340912
rect 75328 340892 75330 340912
rect 75274 340856 75330 340892
rect 74262 284144 74318 284200
rect 75826 312432 75882 312488
rect 77206 390360 77262 390416
rect 76010 389000 76066 389056
rect 76746 389000 76802 389056
rect 75826 301416 75882 301472
rect 77482 390632 77538 390688
rect 78954 389000 79010 389056
rect 78586 383696 78642 383752
rect 77298 338680 77354 338736
rect 76746 322904 76802 322960
rect 76654 318688 76710 318744
rect 77942 320728 77998 320784
rect 80058 387912 80114 387968
rect 82082 391040 82138 391096
rect 85486 391040 85542 391096
rect 81530 388728 81586 388784
rect 80978 387640 81034 387696
rect 79966 385056 80022 385112
rect 79874 304136 79930 304192
rect 81254 377304 81310 377360
rect 78770 292576 78826 292632
rect 79874 292576 79930 292632
rect 77390 283600 77446 283656
rect 82726 387640 82782 387696
rect 82634 333240 82690 333296
rect 81346 319504 81402 319560
rect 80794 287272 80850 287328
rect 85394 380160 85450 380216
rect 85302 378664 85358 378720
rect 83554 339516 83610 339552
rect 83554 339496 83556 339516
rect 83556 339496 83608 339516
rect 83608 339496 83610 339516
rect 84106 329024 84162 329080
rect 83462 323584 83518 323640
rect 82634 285912 82690 285968
rect 84106 289040 84162 289096
rect 86222 389000 86278 389056
rect 86866 382336 86922 382392
rect 86222 369008 86278 369064
rect 85670 320864 85726 320920
rect 85486 291352 85542 291408
rect 85302 287272 85358 287328
rect 89672 391040 89728 391096
rect 92754 391040 92810 391096
rect 88246 373224 88302 373280
rect 89166 389000 89222 389056
rect 89626 387096 89682 387152
rect 89534 385600 89590 385656
rect 88154 319368 88210 319424
rect 88062 291216 88118 291272
rect 87510 285368 87566 285424
rect 89166 287408 89222 287464
rect 89442 287408 89498 287464
rect 93214 389000 93270 389056
rect 91098 382336 91154 382392
rect 93858 388864 93914 388920
rect 93766 386960 93822 387016
rect 93674 364928 93730 364984
rect 92386 332696 92442 332752
rect 92386 322088 92442 322144
rect 91190 312024 91246 312080
rect 92386 312024 92442 312080
rect 91006 308352 91062 308408
rect 89718 292576 89774 292632
rect 89626 288496 89682 288552
rect 90822 289856 90878 289912
rect 93674 304136 93730 304192
rect 94594 388864 94650 388920
rect 98458 389272 98514 389328
rect 97814 385600 97870 385656
rect 97998 381520 98054 381576
rect 95054 285640 95110 285696
rect 94134 285504 94190 285560
rect 94962 285504 95018 285560
rect 94134 284416 94190 284472
rect 95698 283464 95754 283520
rect 97722 321000 97778 321056
rect 96710 285504 96766 285560
rect 97722 285504 97778 285560
rect 96710 284280 96766 284336
rect 96802 283464 96858 283520
rect 69018 282376 69074 282432
rect 100666 390904 100722 390960
rect 99746 389000 99802 389056
rect 100114 389000 100170 389056
rect 99470 388320 99526 388376
rect 99286 329876 99288 329896
rect 99288 329876 99340 329896
rect 99340 329876 99342 329896
rect 99286 329840 99342 329876
rect 100666 388456 100722 388512
rect 102046 387096 102102 387152
rect 100022 285640 100078 285696
rect 99378 280200 99434 280256
rect 99194 273264 99250 273320
rect 99194 272040 99250 272096
rect 98734 267008 98790 267064
rect 98090 262112 98146 262168
rect 98642 262112 98698 262168
rect 98642 261024 98698 261080
rect 98090 259528 98146 259584
rect 68788 241304 68844 241360
rect 68650 232600 68706 232656
rect 68558 140800 68614 140856
rect 69386 240080 69442 240136
rect 70122 241712 70178 241768
rect 71134 241712 71190 241768
rect 70582 240760 70638 240816
rect 70398 240080 70454 240136
rect 70398 239808 70454 239864
rect 69846 136856 69902 136912
rect 71042 240080 71098 240136
rect 71686 233824 71742 233880
rect 71686 134680 71742 134736
rect 71962 140800 72018 140856
rect 72790 241712 72846 241768
rect 74262 241712 74318 241768
rect 91558 241712 91614 241768
rect 72422 239944 72478 240000
rect 72698 239944 72754 240000
rect 74262 238720 74318 238776
rect 74630 238720 74686 238776
rect 72422 230560 72478 230616
rect 72146 138080 72202 138136
rect 74538 230560 74594 230616
rect 73250 135904 73306 135960
rect 73802 137264 73858 137320
rect 76562 225528 76618 225584
rect 76884 241440 76940 241496
rect 78034 240216 78090 240272
rect 78770 234504 78826 234560
rect 77574 232600 77630 232656
rect 78586 226888 78642 226944
rect 82082 240080 82138 240136
rect 81438 237904 81494 237960
rect 79322 228248 79378 228304
rect 78862 224168 78918 224224
rect 81070 138624 81126 138680
rect 80426 137420 80482 137456
rect 80426 137400 80428 137420
rect 80428 137400 80480 137420
rect 80480 137400 80482 137420
rect 81530 226072 81586 226128
rect 85486 239944 85542 240000
rect 84014 210296 84070 210352
rect 83094 206216 83150 206272
rect 84198 207576 84254 207632
rect 84474 141344 84530 141400
rect 86866 239944 86922 240000
rect 86774 234096 86830 234152
rect 85670 233280 85726 233336
rect 86774 233280 86830 233336
rect 85578 231240 85634 231296
rect 85578 231104 85634 231160
rect 86222 213152 86278 213208
rect 88338 235320 88394 235376
rect 86866 137284 86922 137320
rect 86866 137264 86868 137284
rect 86868 137264 86920 137284
rect 86920 137264 86922 137284
rect 87326 136720 87382 136776
rect 90914 237360 90970 237416
rect 89718 237088 89774 237144
rect 88798 139984 88854 140040
rect 90822 211792 90878 211848
rect 90914 206352 90970 206408
rect 91190 237360 91246 237416
rect 92294 227704 92350 227760
rect 92294 227024 92350 227080
rect 92662 235456 92718 235512
rect 92478 220632 92534 220688
rect 92478 148280 92534 148336
rect 92386 135224 92442 135280
rect 93858 233824 93914 233880
rect 93766 207712 93822 207768
rect 92754 200640 92810 200696
rect 94686 227704 94742 227760
rect 94962 241576 95018 241632
rect 94962 137400 95018 137456
rect 94870 134544 94926 134600
rect 95882 241712 95938 241768
rect 95882 217232 95938 217288
rect 95330 216688 95386 216744
rect 95882 216688 95938 216744
rect 95238 124072 95294 124128
rect 69570 92656 69626 92712
rect 69708 92656 69764 92712
rect 70812 92622 70868 92678
rect 68558 92384 68614 92440
rect 70306 92520 70362 92576
rect 72238 91024 72294 91080
rect 71134 90888 71190 90944
rect 69846 84088 69902 84144
rect 67546 47504 67602 47560
rect 70214 11600 70270 11656
rect 74814 88168 74870 88224
rect 75734 92384 75790 92440
rect 77942 90752 77998 90808
rect 77482 90616 77538 90672
rect 74446 28192 74502 28248
rect 72514 25472 72570 25528
rect 80610 90752 80666 90808
rect 81438 90888 81494 90944
rect 82082 89664 82138 89720
rect 83002 88032 83058 88088
rect 79506 85448 79562 85504
rect 77206 73752 77262 73808
rect 84658 86808 84714 86864
rect 83554 85312 83610 85368
rect 77390 4800 77446 4856
rect 83462 72392 83518 72448
rect 85486 29552 85542 29608
rect 87602 76472 87658 76528
rect 89810 92248 89866 92304
rect 91282 92384 91338 92440
rect 90730 90888 90786 90944
rect 92570 91432 92626 91488
rect 95146 94288 95202 94344
rect 92754 91024 92810 91080
rect 92570 90616 92626 90672
rect 89534 89528 89590 89584
rect 88706 88168 88762 88224
rect 89534 88168 89590 88224
rect 89534 87896 89590 87952
rect 85670 3440 85726 3496
rect 88982 3304 89038 3360
rect 93858 92384 93914 92440
rect 95054 91432 95110 91488
rect 91006 71032 91062 71088
rect 92386 30912 92442 30968
rect 97814 240080 97870 240136
rect 97906 234640 97962 234696
rect 97446 230288 97502 230344
rect 96710 220224 96766 220280
rect 97354 204856 97410 204912
rect 96710 133048 96766 133104
rect 96618 132232 96674 132288
rect 97446 133864 97502 133920
rect 97354 131416 97410 131472
rect 97262 130872 97318 130928
rect 96710 129240 96766 129296
rect 97170 127608 97226 127664
rect 96802 125432 96858 125488
rect 96618 123972 96620 123992
rect 96620 123972 96672 123992
rect 96672 123972 96674 123992
rect 96618 123936 96674 123972
rect 96618 117036 96620 117056
rect 96620 117036 96672 117056
rect 96672 117036 96674 117056
rect 96618 117000 96674 117036
rect 96618 114008 96674 114064
rect 95974 111832 96030 111888
rect 95974 101360 96030 101416
rect 95974 88032 96030 88088
rect 97170 104216 97226 104272
rect 97170 102856 97226 102912
rect 97538 127064 97594 127120
rect 97814 126248 97870 126304
rect 97446 124616 97502 124672
rect 97814 123256 97870 123312
rect 97814 122440 97870 122496
rect 97814 120808 97870 120864
rect 97814 120264 97870 120320
rect 97814 117816 97870 117872
rect 97814 116456 97870 116512
rect 97814 115640 97870 115696
rect 97722 114824 97778 114880
rect 97814 112648 97870 112704
rect 98642 233824 98698 233880
rect 99102 233824 99158 233880
rect 97998 232600 98054 232656
rect 97906 111016 97962 111072
rect 97906 110200 97962 110256
rect 97814 109656 97870 109712
rect 97722 108024 97778 108080
rect 97538 106664 97594 106720
rect 97906 108840 97962 108896
rect 97906 105848 97962 105904
rect 97630 105032 97686 105088
rect 97354 100000 97410 100056
rect 97906 102076 97908 102096
rect 97908 102076 97960 102096
rect 97960 102076 97962 102096
rect 97906 102040 97962 102076
rect 97814 101224 97870 101280
rect 97906 100408 97962 100464
rect 97722 99592 97778 99648
rect 97538 98232 97594 98288
rect 97906 97416 97962 97472
rect 97538 96600 97594 96656
rect 97906 95240 97962 95296
rect 97906 94424 97962 94480
rect 97906 93608 97962 93664
rect 97354 92792 97410 92848
rect 99102 214648 99158 214704
rect 98642 115096 98698 115152
rect 98734 111016 98790 111072
rect 100574 287408 100630 287464
rect 100574 283464 100630 283520
rect 100666 282376 100722 282432
rect 100758 281016 100814 281072
rect 100758 278704 100814 278760
rect 100758 275324 100814 275360
rect 100758 275304 100760 275324
rect 100760 275304 100812 275324
rect 100812 275304 100814 275324
rect 100850 274488 100906 274544
rect 100758 273672 100814 273728
rect 101494 280200 101550 280256
rect 101586 279384 101642 279440
rect 101954 278568 102010 278624
rect 103518 389136 103574 389192
rect 102322 388456 102378 388512
rect 103794 389136 103850 389192
rect 102230 335416 102286 335472
rect 102138 326984 102194 327040
rect 102782 323584 102838 323640
rect 102046 277752 102102 277808
rect 102046 276120 102102 276176
rect 101954 275848 102010 275904
rect 101402 272040 101458 272096
rect 101678 271224 101734 271280
rect 100758 269592 100814 269648
rect 100850 268776 100906 268832
rect 100758 267960 100814 268016
rect 101402 267144 101458 267200
rect 100022 265512 100078 265568
rect 99470 252456 99526 252512
rect 99470 234640 99526 234696
rect 100758 264696 100814 264752
rect 100758 263880 100814 263936
rect 100758 263064 100814 263120
rect 100850 262248 100906 262304
rect 100758 261468 100760 261488
rect 100760 261468 100812 261488
rect 100812 261468 100814 261488
rect 100758 261432 100814 261468
rect 100850 260616 100906 260672
rect 100850 258984 100906 259040
rect 100758 258168 100814 258224
rect 100390 252492 100392 252512
rect 100392 252492 100444 252512
rect 100444 252492 100446 252512
rect 100390 252456 100446 252492
rect 100022 233960 100078 234016
rect 100574 229744 100630 229800
rect 100574 218592 100630 218648
rect 100850 257352 100906 257408
rect 101034 257216 101090 257272
rect 100942 256536 100998 256592
rect 100850 255720 100906 255776
rect 101034 254088 101090 254144
rect 100850 250824 100906 250880
rect 100850 250008 100906 250064
rect 100850 249192 100906 249248
rect 100942 248376 100998 248432
rect 100850 247560 100906 247616
rect 100850 246744 100906 246800
rect 100850 245928 100906 245984
rect 100850 245112 100906 245168
rect 100942 244296 100998 244352
rect 100850 242700 100852 242720
rect 100852 242700 100904 242720
rect 100904 242700 100906 242720
rect 100850 242664 100906 242700
rect 100850 241848 100906 241904
rect 101494 254904 101550 254960
rect 101402 235456 101458 235512
rect 103426 318144 103482 318200
rect 102322 273264 102378 273320
rect 103518 289040 103574 289096
rect 104254 304136 104310 304192
rect 104438 304136 104494 304192
rect 104346 271088 104402 271144
rect 103978 270408 104034 270464
rect 104346 262112 104402 262168
rect 105266 390360 105322 390416
rect 104898 383560 104954 383616
rect 104898 382336 104954 382392
rect 104162 240080 104218 240136
rect 102782 237088 102838 237144
rect 99378 204856 99434 204912
rect 98642 90888 98698 90944
rect 100758 134544 100814 134600
rect 103426 225936 103482 225992
rect 102874 199960 102930 200016
rect 102874 128424 102930 128480
rect 102046 104080 102102 104136
rect 101034 7520 101090 7576
rect 98642 3576 98698 3632
rect 102230 87896 102286 87952
rect 104806 228248 104862 228304
rect 104162 137264 104218 137320
rect 104162 124752 104218 124808
rect 103610 85448 103666 85504
rect 105082 262112 105138 262168
rect 104990 207576 105046 207632
rect 106186 322088 106242 322144
rect 105634 270408 105690 270464
rect 106094 256264 106150 256320
rect 113270 440952 113326 441008
rect 113270 431160 113326 431216
rect 113178 429256 113234 429312
rect 113178 420008 113234 420064
rect 107750 390632 107806 390688
rect 108762 390632 108818 390688
rect 111706 390632 111762 390688
rect 106738 390360 106794 390416
rect 105542 236544 105598 236600
rect 106830 269184 106886 269240
rect 107750 389000 107806 389056
rect 108946 389000 109002 389056
rect 107014 284144 107070 284200
rect 107566 284144 107622 284200
rect 106646 249076 106702 249112
rect 106646 249056 106648 249076
rect 106648 249056 106700 249076
rect 106700 249056 106702 249076
rect 107658 239944 107714 240000
rect 107658 237904 107714 237960
rect 105634 85312 105690 85368
rect 105726 8880 105782 8936
rect 105542 3440 105598 3496
rect 110694 387776 110750 387832
rect 109682 324944 109738 325000
rect 109038 246200 109094 246256
rect 109038 207712 109094 207768
rect 109682 273128 109738 273184
rect 111706 330384 111762 330440
rect 109314 206216 109370 206272
rect 109314 101360 109370 101416
rect 113454 430072 113510 430128
rect 113362 416744 113418 416800
rect 113822 429256 113878 429312
rect 111706 186904 111762 186960
rect 109038 91024 109094 91080
rect 111890 214648 111946 214704
rect 112258 271924 112314 271960
rect 112258 271904 112260 271924
rect 112260 271904 112312 271924
rect 112312 271904 112314 271924
rect 114098 424904 114154 424960
rect 115202 435240 115258 435296
rect 114742 432248 114798 432304
rect 114742 431160 114798 431216
rect 114650 424088 114706 424144
rect 115386 428168 115442 428224
rect 115846 425992 115902 426048
rect 115846 424088 115902 424144
rect 115846 423000 115902 423056
rect 114742 418920 114798 418976
rect 114650 417832 114706 417888
rect 114558 406408 114614 406464
rect 115846 421948 115848 421968
rect 115848 421948 115900 421968
rect 115900 421948 115902 421968
rect 115846 421912 115902 421948
rect 115846 416780 115848 416800
rect 115848 416780 115900 416800
rect 115900 416780 115902 416800
rect 115846 416744 115902 416780
rect 115202 415692 115204 415712
rect 115204 415692 115256 415712
rect 115256 415692 115258 415712
rect 115202 415656 115258 415692
rect 115846 414876 115848 414896
rect 115848 414876 115900 414896
rect 115900 414876 115902 414896
rect 115846 414840 115902 414876
rect 115846 413752 115902 413808
rect 115202 412664 115258 412720
rect 115846 411576 115902 411632
rect 115846 410524 115848 410544
rect 115848 410524 115900 410544
rect 115900 410524 115902 410544
rect 115846 410488 115902 410524
rect 115846 409672 115902 409728
rect 115846 407496 115902 407552
rect 114926 406408 114982 406464
rect 115846 405592 115902 405648
rect 115570 404504 115626 404560
rect 115846 403416 115902 403472
rect 115662 401240 115718 401296
rect 115018 400444 115074 400480
rect 115018 400424 115020 400444
rect 115020 400424 115072 400444
rect 115072 400424 115074 400444
rect 115202 399336 115258 399392
rect 115846 398248 115902 398304
rect 115846 397160 115902 397216
rect 115846 396344 115902 396400
rect 115846 395256 115902 395312
rect 115570 394168 115626 394224
rect 115846 393116 115848 393136
rect 115848 393116 115900 393136
rect 115900 393116 115902 393136
rect 115846 393080 115902 393116
rect 115846 392012 115902 392048
rect 115846 391992 115848 392012
rect 115848 391992 115900 392012
rect 115900 391992 115902 392012
rect 116582 536696 116638 536752
rect 114742 318144 114798 318200
rect 114650 307808 114706 307864
rect 114650 285912 114706 285968
rect 114558 283464 114614 283520
rect 115018 263608 115074 263664
rect 115846 285912 115902 285968
rect 114650 234504 114706 234560
rect 114558 206352 114614 206408
rect 110510 3440 110566 3496
rect 109314 3304 109370 3360
rect 114558 92248 114614 92304
rect 117318 442992 117374 443048
rect 116122 402328 116178 402384
rect 117502 439456 117558 439512
rect 117502 383560 117558 383616
rect 116030 291796 116032 291816
rect 116032 291796 116084 291816
rect 116084 291796 116086 291816
rect 116030 291760 116086 291796
rect 116030 287272 116086 287328
rect 115846 224168 115902 224224
rect 114650 86808 114706 86864
rect 115754 86808 115810 86864
rect 115754 86128 115810 86184
rect 116582 288496 116638 288552
rect 116122 284144 116178 284200
rect 116858 271904 116914 271960
rect 120078 437552 120134 437608
rect 118882 320864 118938 320920
rect 118790 275984 118846 276040
rect 118790 274624 118846 274680
rect 117962 237904 118018 237960
rect 117686 235320 117742 235376
rect 117410 206896 117466 206952
rect 117410 206352 117466 206408
rect 117318 138624 117374 138680
rect 116766 111016 116822 111072
rect 116398 3576 116454 3632
rect 112810 3440 112866 3496
rect 119342 324944 119398 325000
rect 122838 582392 122894 582448
rect 121458 389000 121514 389056
rect 120078 320728 120134 320784
rect 120170 282920 120226 282976
rect 119066 208256 119122 208312
rect 119066 207576 119122 207632
rect 120170 246200 120226 246256
rect 120354 210976 120410 211032
rect 120722 210976 120778 211032
rect 120354 210296 120410 210352
rect 124402 434696 124458 434752
rect 124126 396616 124182 396672
rect 121642 304136 121698 304192
rect 122102 292576 122158 292632
rect 121642 291216 121698 291272
rect 121550 275848 121606 275904
rect 121550 274624 121606 274680
rect 121458 206216 121514 206272
rect 121642 141344 121698 141400
rect 120262 121488 120318 121544
rect 122930 234504 122986 234560
rect 122930 233824 122986 233880
rect 124402 322088 124458 322144
rect 125506 322088 125562 322144
rect 125598 312024 125654 312080
rect 124310 244316 124366 244352
rect 124310 244296 124312 244316
rect 124312 244296 124364 244316
rect 124364 244296 124366 244316
rect 124310 212472 124366 212528
rect 126886 383696 126942 383752
rect 125782 251776 125838 251832
rect 125690 218592 125746 218648
rect 125598 139984 125654 140040
rect 126242 241304 126298 241360
rect 126886 221992 126942 222048
rect 127070 263608 127126 263664
rect 128450 309032 128506 309088
rect 128450 308352 128506 308408
rect 128358 208120 128414 208176
rect 128358 207712 128414 207768
rect 127254 95512 127310 95568
rect 129738 234504 129794 234560
rect 129738 232600 129794 232656
rect 128634 211792 128690 211848
rect 129002 108296 129058 108352
rect 131118 219136 131174 219192
rect 131118 218592 131174 218648
rect 132590 396616 132646 396672
rect 132590 258712 132646 258768
rect 135258 278704 135314 278760
rect 133786 258732 133842 258768
rect 133786 258712 133788 258732
rect 133788 258712 133840 258732
rect 133840 258712 133842 258732
rect 134522 215872 134578 215928
rect 133878 113328 133934 113384
rect 126242 3440 126298 3496
rect 135350 244840 135406 244896
rect 136638 192480 136694 192536
rect 136454 4936 136510 4992
rect 138018 220224 138074 220280
rect 141422 323584 141478 323640
rect 140778 235320 140834 235376
rect 141422 225528 141478 225584
rect 139490 213832 139546 213888
rect 139490 213152 139546 213208
rect 142986 251776 143042 251832
rect 143538 248240 143594 248296
rect 143538 247560 143594 247616
rect 142894 241304 142950 241360
rect 146298 233008 146354 233064
rect 151082 302504 151138 302560
rect 180154 313384 180210 313440
rect 152462 307808 152518 307864
rect 178774 306584 178830 306640
rect 156602 276664 156658 276720
rect 157982 257216 158038 257272
rect 166354 298832 166410 298888
rect 166262 291760 166318 291816
rect 160926 242800 160982 242856
rect 173346 237224 173402 237280
rect 178682 301552 178738 301608
rect 179418 295296 179474 295352
rect 178682 241576 178738 241632
rect 185674 309304 185730 309360
rect 185582 305088 185638 305144
rect 181534 261024 181590 261080
rect 186318 301416 186374 301472
rect 185674 284824 185730 284880
rect 187054 306720 187110 306776
rect 184294 257216 184350 257272
rect 184386 247016 184442 247072
rect 188342 317464 188398 317520
rect 188526 310800 188582 310856
rect 188342 309440 188398 309496
rect 188526 306312 188582 306368
rect 188434 301280 188490 301336
rect 189814 304952 189870 305008
rect 191378 307944 191434 308000
rect 191286 302368 191342 302424
rect 191194 300872 191250 300928
rect 191102 299920 191158 299976
rect 191194 292168 191250 292224
rect 190826 287408 190882 287464
rect 190366 284280 190422 284336
rect 191746 298968 191802 299024
rect 191470 297472 191526 297528
rect 191470 296792 191526 296848
rect 191746 296112 191802 296168
rect 191654 294208 191710 294264
rect 191746 293120 191802 293176
rect 191378 291760 191434 291816
rect 191286 282784 191342 282840
rect 191654 291216 191710 291272
rect 201590 320184 201646 320240
rect 193770 316240 193826 316296
rect 200302 311888 200358 311944
rect 199658 306448 199714 306504
rect 192574 301688 192630 301744
rect 191746 290264 191802 290320
rect 191746 289312 191802 289368
rect 191654 289040 191710 289096
rect 195518 303864 195574 303920
rect 197910 303592 197966 303648
rect 197542 301688 197598 301744
rect 200394 310664 200450 310720
rect 203246 313248 203302 313304
rect 207754 307944 207810 308000
rect 204258 306584 204314 306640
rect 206006 305088 206062 305144
rect 208398 306720 208454 306776
rect 222198 316104 222254 316160
rect 214562 314880 214618 314936
rect 213182 313384 213238 313440
rect 209778 309440 209834 309496
rect 211894 304952 211950 305008
rect 218518 314744 218574 314800
rect 219622 310528 219678 310584
rect 220818 309168 220874 309224
rect 227718 317464 227774 317520
rect 226982 315288 227038 315344
rect 226982 304952 227038 305008
rect 234618 307808 234674 307864
rect 229374 303728 229430 303784
rect 230478 303592 230534 303648
rect 238666 303864 238722 303920
rect 238022 302232 238078 302288
rect 194230 301416 194286 301472
rect 197542 301416 197598 301472
rect 194506 301144 194562 301200
rect 212814 301144 212870 301200
rect 224958 301144 225014 301200
rect 210422 301008 210478 301064
rect 216310 301008 216366 301064
rect 220358 301008 220414 301064
rect 222750 301008 222806 301064
rect 224406 301008 224462 301064
rect 231398 301008 231454 301064
rect 232594 301008 232650 301064
rect 233790 301008 233846 301064
rect 235446 301008 235502 301064
rect 196070 300872 196126 300928
rect 198186 300872 198242 300928
rect 198830 300872 198886 300928
rect 202326 300872 202382 300928
rect 203062 300872 203118 300928
rect 204626 300872 204682 300928
rect 206282 300872 206338 300928
rect 207110 300872 207166 300928
rect 209318 300872 209374 300928
rect 212170 300872 212226 300928
rect 214286 300872 214342 300928
rect 215114 300872 215170 300928
rect 216678 300872 216734 300928
rect 217322 300872 217378 300928
rect 219530 300872 219586 300928
rect 221462 300872 221518 300928
rect 223210 300872 223266 300928
rect 224038 300872 224094 300928
rect 225602 300872 225658 300928
rect 226338 300872 226394 300928
rect 227258 300872 227314 300928
rect 228454 300872 228510 300928
rect 229742 300872 229798 300928
rect 231030 300872 231086 300928
rect 232318 300872 232374 300928
rect 233330 300872 233386 300928
rect 234894 300872 234950 300928
rect 236734 300872 236790 300928
rect 237838 300872 237894 300928
rect 238850 300872 238906 300928
rect 248418 338680 248474 338736
rect 246302 335416 246358 335472
rect 244922 334056 244978 334112
rect 242162 304952 242218 305008
rect 245014 326304 245070 326360
rect 244922 308896 244978 308952
rect 246210 308896 246266 308952
rect 246210 307808 246266 307864
rect 245658 306448 245714 306504
rect 244830 301416 244886 301472
rect 248418 306992 248474 307048
rect 247682 304136 247738 304192
rect 246854 302504 246910 302560
rect 246854 302232 246910 302288
rect 249706 303592 249762 303648
rect 248878 302776 248934 302832
rect 247774 301552 247830 301608
rect 249798 302776 249854 302832
rect 250902 303728 250958 303784
rect 250350 301688 250406 301744
rect 252650 302368 252706 302424
rect 246486 301416 246542 301472
rect 251822 301280 251878 301336
rect 240046 300872 240102 300928
rect 193678 300192 193734 300248
rect 192574 287000 192630 287056
rect 191746 286456 191802 286512
rect 191654 285504 191710 285560
rect 191746 284416 191802 284472
rect 191654 284280 191710 284336
rect 191746 283464 191802 283520
rect 192482 282512 192538 282568
rect 191470 281560 191526 281616
rect 191562 280608 191618 280664
rect 191746 279656 191802 279712
rect 191654 278704 191710 278760
rect 191746 277752 191802 277808
rect 191102 276800 191158 276856
rect 191654 275712 191710 275768
rect 191746 274760 191802 274816
rect 188526 267824 188582 267880
rect 187146 239944 187202 240000
rect 188526 236680 188582 236736
rect 191746 272856 191802 272912
rect 191194 271940 191196 271960
rect 191196 271940 191248 271960
rect 191248 271940 191250 271960
rect 191194 271904 191250 271940
rect 191102 270952 191158 271008
rect 191010 264152 191066 264208
rect 191010 262268 191066 262304
rect 191010 262248 191012 262268
rect 191012 262248 191064 262268
rect 191064 262248 191066 262268
rect 190642 258304 190698 258360
rect 189722 255720 189778 255776
rect 188986 213152 189042 213208
rect 188342 86264 188398 86320
rect 191010 253544 191066 253600
rect 190642 249600 190698 249656
rect 189814 248512 189870 248568
rect 189906 245656 189962 245712
rect 191746 270000 191802 270056
rect 191654 269048 191710 269104
rect 253202 304136 253258 304192
rect 252834 286320 252890 286376
rect 258262 332560 258318 332616
rect 256790 328480 256846 328536
rect 253938 312432 253994 312488
rect 253294 301552 253350 301608
rect 253478 301416 253534 301472
rect 253202 300464 253258 300520
rect 253478 298696 253534 298752
rect 252926 284144 252982 284200
rect 252834 281288 252890 281344
rect 193218 276800 193274 276856
rect 193126 273808 193182 273864
rect 191470 267008 191526 267064
rect 191746 266056 191802 266112
rect 191286 265104 191342 265160
rect 191194 263200 191250 263256
rect 189906 232464 189962 232520
rect 191378 261296 191434 261352
rect 191746 260344 191802 260400
rect 191746 257352 191802 257408
rect 191746 255448 191802 255504
rect 191562 254496 191618 254552
rect 191746 252612 191802 252648
rect 191746 252592 191748 252612
rect 191748 252592 191800 252612
rect 191800 252592 191802 252612
rect 191562 251640 191618 251696
rect 191746 250688 191802 250744
rect 191746 247696 191802 247752
rect 191562 245792 191618 245848
rect 191746 243888 191802 243944
rect 191838 239808 191894 239864
rect 191378 236544 191434 236600
rect 192482 236544 192538 236600
rect 254030 292440 254086 292496
rect 254214 289312 254270 289368
rect 254122 284280 254178 284336
rect 255410 295704 255466 295760
rect 255410 294752 255466 294808
rect 255410 293392 255466 293448
rect 255410 292068 255412 292088
rect 255412 292068 255464 292088
rect 255464 292068 255466 292088
rect 255410 292032 255466 292068
rect 255410 290672 255466 290728
rect 255410 289740 255466 289776
rect 255410 289720 255412 289740
rect 255412 289720 255464 289740
rect 255464 289720 255466 289740
rect 255410 288380 255466 288416
rect 255410 288360 255412 288380
rect 255412 288360 255464 288380
rect 255464 288360 255466 288380
rect 255686 300736 255742 300792
rect 255870 300192 255926 300248
rect 255686 299396 255742 299432
rect 255686 299376 255688 299396
rect 255688 299376 255740 299396
rect 255740 299376 255742 299396
rect 255778 298832 255834 298888
rect 255686 298016 255742 298072
rect 255778 297064 255834 297120
rect 255686 296520 255742 296576
rect 255686 292984 255742 293040
rect 255778 291488 255834 291544
rect 255686 290128 255742 290184
rect 255686 288768 255742 288824
rect 255686 287408 255742 287464
rect 255594 287000 255650 287056
rect 255502 286456 255558 286512
rect 255410 285096 255466 285152
rect 255410 284688 255466 284744
rect 255410 283328 255466 283384
rect 255410 282804 255466 282840
rect 255410 282784 255412 282804
rect 255412 282784 255464 282804
rect 255464 282784 255466 282804
rect 255502 281968 255558 282024
rect 255502 281016 255558 281072
rect 255410 280608 255466 280664
rect 255410 280084 255466 280120
rect 255410 280064 255412 280084
rect 255412 280064 255464 280084
rect 255464 280064 255466 280084
rect 255594 279656 255650 279712
rect 255318 279248 255374 279304
rect 255318 278704 255374 278760
rect 255410 278296 255466 278352
rect 256606 278024 256662 278080
rect 255410 277752 255466 277808
rect 255502 277344 255558 277400
rect 255318 276936 255374 276992
rect 256606 276392 256662 276448
rect 255410 275576 255466 275632
rect 255594 275032 255650 275088
rect 255410 274216 255466 274272
rect 254030 273672 254086 273728
rect 253938 273264 253994 273320
rect 253938 272720 253994 272776
rect 252926 269320 252982 269376
rect 193402 258848 193458 258904
rect 193678 242800 193734 242856
rect 204902 239944 204958 240000
rect 206374 239944 206430 240000
rect 200762 227024 200818 227080
rect 195242 200640 195298 200696
rect 152462 3304 152518 3360
rect 206282 200640 206338 200696
rect 220818 240080 220874 240136
rect 213182 202816 213238 202872
rect 227258 239944 227314 240000
rect 234710 240080 234766 240136
rect 234618 228792 234674 228848
rect 240782 239400 240838 239456
rect 238666 238312 238722 238368
rect 238666 229064 238722 229120
rect 238666 228792 238722 228848
rect 238666 219408 238722 219464
rect 238666 219000 238722 219056
rect 238666 209752 238722 209808
rect 238666 209480 238722 209536
rect 240782 222128 240838 222184
rect 238666 200096 238722 200152
rect 238666 199824 238722 199880
rect 238666 190440 238722 190496
rect 238666 190304 238722 190360
rect 238666 180784 238722 180840
rect 238666 180648 238722 180704
rect 238666 171128 238722 171184
rect 238666 170992 238722 171048
rect 238666 161472 238722 161528
rect 238666 161336 238722 161392
rect 238666 151816 238722 151872
rect 238666 151680 238722 151736
rect 238666 145560 238722 145616
rect 233146 101396 233148 101416
rect 233148 101396 233200 101416
rect 233200 101396 233202 101416
rect 233146 101360 233202 101396
rect 220818 91704 220874 91760
rect 239310 3984 239366 4040
rect 231122 3848 231178 3904
rect 240506 3440 240562 3496
rect 244278 237360 244334 237416
rect 242162 3304 242218 3360
rect 246394 239536 246450 239592
rect 244922 216688 244978 216744
rect 244278 3848 244334 3904
rect 244278 3576 244334 3632
rect 245198 3576 245254 3632
rect 244922 3440 244978 3496
rect 249062 237360 249118 237416
rect 246394 216552 246450 216608
rect 250534 241168 250590 241224
rect 250442 238448 250498 238504
rect 249246 227024 249302 227080
rect 249062 138624 249118 138680
rect 250534 204176 250590 204232
rect 252650 238584 252706 238640
rect 251822 226208 251878 226264
rect 251914 219272 251970 219328
rect 252834 267552 252890 267608
rect 252926 252456 252982 252512
rect 253202 247832 253258 247888
rect 253110 246064 253166 246120
rect 253018 243752 253074 243808
rect 253018 241984 253074 242040
rect 252742 208120 252798 208176
rect 255502 272312 255558 272368
rect 255410 271924 255466 271960
rect 255410 271904 255412 271924
rect 255412 271904 255464 271924
rect 255464 271904 255466 271924
rect 255502 271360 255558 271416
rect 255318 270952 255374 271008
rect 255410 270000 255466 270056
rect 256606 274624 256662 274680
rect 256882 319368 256938 319424
rect 256790 295160 256846 295216
rect 256882 285640 256938 285696
rect 257066 275984 257122 276040
rect 257342 275984 257398 276040
rect 258078 275984 258134 276040
rect 255502 269048 255558 269104
rect 256698 272448 256754 272504
rect 256514 269728 256570 269784
rect 255410 267280 255466 267336
rect 255410 266872 255466 266928
rect 255502 266464 255558 266520
rect 255318 265512 255374 265568
rect 255410 263644 255412 263664
rect 255412 263644 255464 263664
rect 255464 263644 255466 263664
rect 255410 263608 255466 263644
rect 255410 263200 255466 263256
rect 255410 259528 255466 259584
rect 255410 258984 255466 259040
rect 256606 268640 256662 268696
rect 256514 266328 256570 266384
rect 255870 259936 255926 259992
rect 255502 258576 255558 258632
rect 255410 257624 255466 257680
rect 255410 256264 255466 256320
rect 255502 255856 255558 255912
rect 255410 254904 255466 254960
rect 255594 254496 255650 254552
rect 255502 253544 255558 253600
rect 255410 253136 255466 253192
rect 255502 252184 255558 252240
rect 255410 251776 255466 251832
rect 255318 251232 255374 251288
rect 255318 250280 255374 250336
rect 255410 249872 255466 249928
rect 254582 249192 254638 249248
rect 255318 248920 255374 248976
rect 255410 247560 255466 247616
rect 255318 246744 255374 246800
rect 255410 245792 255466 245848
rect 255318 244296 255374 244352
rect 255502 245248 255558 245304
rect 256606 264016 256662 264072
rect 256882 261296 256938 261352
rect 255962 254496 256018 254552
rect 255686 252592 255742 252648
rect 255686 248512 255742 248568
rect 255594 244840 255650 244896
rect 255410 243480 255466 243536
rect 255318 242528 255374 242584
rect 255410 241984 255466 242040
rect 255410 241712 255466 241768
rect 255962 242120 256018 242176
rect 255410 235728 255466 235784
rect 255502 230560 255558 230616
rect 256882 241304 256938 241360
rect 254674 3440 254730 3496
rect 257066 206896 257122 206952
rect 259550 287952 259606 288008
rect 258354 255992 258410 256048
rect 258354 247152 258410 247208
rect 258354 235864 258410 235920
rect 259642 270544 259698 270600
rect 259734 239400 259790 239456
rect 259642 224848 259698 224904
rect 258262 213832 258318 213888
rect 263690 332696 263746 332752
rect 262402 331200 262458 331256
rect 262310 320728 262366 320784
rect 262126 297372 262128 297392
rect 262128 297372 262180 297392
rect 262180 297372 262182 297392
rect 262126 297336 262182 297372
rect 261482 295976 261538 296032
rect 260746 244316 260802 244352
rect 260746 244296 260748 244316
rect 260748 244296 260800 244316
rect 260800 244296 260802 244316
rect 260930 233008 260986 233064
rect 262218 266464 262274 266520
rect 262402 297336 262458 297392
rect 262494 251776 262550 251832
rect 262218 212472 262274 212528
rect 260838 210976 260894 211032
rect 262494 228928 262550 228984
rect 265070 321544 265126 321600
rect 263782 312024 263838 312080
rect 263598 282240 263654 282296
rect 262678 256672 262734 256728
rect 263874 250552 263930 250608
rect 266358 272448 266414 272504
rect 266450 269728 266506 269784
rect 266358 264288 266414 264344
rect 268382 264832 268438 264888
rect 266358 215192 266414 215248
rect 267830 257216 267886 257272
rect 266634 240760 266690 240816
rect 267922 254496 267978 254552
rect 268566 264152 268622 264208
rect 268566 257216 268622 257272
rect 268014 224712 268070 224768
rect 268382 224712 268438 224768
rect 267922 220768 267978 220824
rect 269762 268368 269818 268424
rect 269302 260072 269358 260128
rect 269394 230424 269450 230480
rect 269302 219136 269358 219192
rect 271142 265512 271198 265568
rect 270774 223488 270830 223544
rect 348790 702616 348846 702672
rect 543462 702480 543518 702536
rect 276018 310392 276074 310448
rect 276662 310392 276718 310448
rect 276018 309304 276074 309360
rect 272062 278024 272118 278080
rect 270682 205536 270738 205592
rect 273442 267008 273498 267064
rect 273442 266328 273498 266384
rect 273350 208256 273406 208312
rect 583574 696904 583630 696960
rect 582654 683848 582710 683904
rect 582470 670656 582526 670712
rect 580170 644000 580226 644056
rect 285678 309032 285734 309088
rect 286322 309032 286378 309088
rect 276662 306448 276718 306504
rect 277398 304952 277454 305008
rect 274638 84088 274694 84144
rect 274638 83408 274694 83464
rect 280802 297336 280858 297392
rect 284298 297472 284354 297528
rect 285678 236544 285734 236600
rect 295982 302776 296038 302832
rect 291842 251776 291898 251832
rect 290186 3304 290242 3360
rect 295338 141344 295394 141400
rect 299478 294480 299534 294536
rect 305642 307808 305698 307864
rect 582470 630808 582526 630864
rect 579802 590960 579858 591016
rect 580170 537784 580226 537840
rect 580170 511284 580226 511320
rect 580170 511264 580172 511284
rect 580172 511264 580224 511284
rect 580224 511264 580226 511284
rect 582378 458088 582434 458144
rect 580262 365064 580318 365120
rect 580170 325216 580226 325272
rect 321558 306992 321614 307048
rect 309782 260072 309838 260128
rect 318798 124752 318854 124808
rect 320178 83408 320234 83464
rect 327078 302232 327134 302288
rect 324962 300464 325018 300520
rect 324962 3304 325018 3360
rect 333978 289040 334034 289096
rect 332690 3304 332746 3360
rect 345018 301688 345074 301744
rect 342258 284824 342314 284880
rect 339498 283464 339554 283520
rect 336002 3304 336058 3360
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 582378 312024 582434 312080
rect 582562 617480 582618 617536
rect 582562 577632 582618 577688
rect 582746 582392 582802 582448
rect 582746 564304 582802 564360
rect 582654 524456 582710 524512
rect 582562 267008 582618 267064
rect 582746 484608 582802 484664
rect 582654 264152 582710 264208
rect 582838 471416 582894 471472
rect 582470 258848 582526 258904
rect 583114 431568 583170 431624
rect 582930 293120 582986 293176
rect 582378 245520 582434 245576
rect 348054 3984 348110 4040
rect 350446 3304 350502 3360
rect 580170 219000 580226 219056
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 357438 86128 357494 86184
rect 356058 3984 356114 4040
rect 580170 59608 580226 59664
rect 582378 232328 582434 232384
rect 580354 165824 580410 165880
rect 580262 33088 580318 33144
rect 582654 234640 582710 234696
rect 582470 205672 582526 205728
rect 582838 237904 582894 237960
rect 582838 86128 582894 86184
rect 582746 72936 582802 72992
rect 582654 46280 582710 46336
rect 582562 19760 582618 19816
rect 582378 6568 582434 6624
rect 583022 279384 583078 279440
rect 583206 418240 583262 418296
rect 583298 404912 583354 404968
rect 583390 378392 583446 378448
rect 583482 351600 583538 351656
rect 583574 271088 583630 271144
rect 583114 112784 583170 112840
rect 583482 213152 583538 213208
rect 583390 152632 583446 152688
rect 583298 125976 583354 126032
rect 583206 99456 583262 99512
<< metal3 >>
rect 263358 702612 263364 702676
rect 263428 702674 263434 702676
rect 348785 702674 348851 702677
rect 263428 702672 348851 702674
rect 263428 702616 348790 702672
rect 348846 702616 348851 702672
rect 263428 702614 348851 702616
rect 263428 702612 263434 702614
rect 348785 702611 348851 702614
rect 264094 702476 264100 702540
rect 264164 702538 264170 702540
rect 543457 702538 543523 702541
rect 264164 702536 543523 702538
rect 264164 702480 543462 702536
rect 543518 702480 543523 702536
rect 264164 702478 543523 702480
rect 264164 702476 264170 702478
rect 543457 702475 543523 702478
rect -960 697220 480 697460
rect 583520 697234 584960 697324
rect 583342 697174 584960 697234
rect 583342 697098 583402 697174
rect 583520 697098 584960 697174
rect 583342 697084 584960 697098
rect 583342 697038 583586 697084
rect 583526 696965 583586 697038
rect 583526 696960 583635 696965
rect 583526 696904 583574 696960
rect 583630 696904 583635 696960
rect 583526 696902 583635 696904
rect 583569 696899 583635 696902
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582649 683906 582715 683909
rect 583520 683906 584960 683996
rect 582649 683904 584960 683906
rect 582649 683848 582654 683904
rect 582710 683848 584960 683904
rect 582649 683846 584960 683848
rect 582649 683843 582715 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 582465 670714 582531 670717
rect 583520 670714 584960 670804
rect 582465 670712 584960 670714
rect 582465 670656 582470 670712
rect 582526 670656 584960 670712
rect 582465 670654 584960 670656
rect 582465 670651 582531 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582465 630866 582531 630869
rect 583520 630866 584960 630956
rect 582465 630864 584960 630866
rect 582465 630808 582470 630864
rect 582526 630808 584960 630864
rect 582465 630806 584960 630808
rect 582465 630803 582531 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 582557 617538 582623 617541
rect 583520 617538 584960 617628
rect 582557 617536 584960 617538
rect 582557 617480 582562 617536
rect 582618 617480 584960 617536
rect 582557 617478 584960 617480
rect 582557 617475 582623 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 79961 588026 80027 588029
rect 124254 588026 124260 588028
rect 79961 588024 124260 588026
rect 79961 587968 79966 588024
rect 80022 587968 124260 588024
rect 79961 587966 124260 587968
rect 79961 587963 80027 587966
rect 124254 587964 124260 587966
rect 124324 587964 124330 588028
rect 72417 585170 72483 585173
rect 101397 585170 101463 585173
rect 72417 585168 101463 585170
rect 72417 585112 72422 585168
rect 72478 585112 101402 585168
rect 101458 585112 101463 585168
rect 72417 585110 101463 585112
rect 72417 585107 72483 585110
rect 101397 585107 101463 585110
rect 71773 584898 71839 584901
rect 75862 584898 75868 584900
rect 71773 584896 75868 584898
rect 71773 584840 71778 584896
rect 71834 584840 75868 584896
rect 71773 584838 75868 584840
rect 71773 584835 71839 584838
rect 75862 584836 75868 584838
rect 75932 584836 75938 584900
rect 82721 583810 82787 583813
rect 111742 583810 111748 583812
rect 82721 583808 111748 583810
rect 82721 583752 82726 583808
rect 82782 583752 111748 583808
rect 82721 583750 111748 583752
rect 82721 583747 82787 583750
rect 111742 583748 111748 583750
rect 111812 583748 111818 583812
rect 79041 582722 79107 582725
rect 89713 582722 89779 582725
rect 79041 582720 89779 582722
rect 79041 582664 79046 582720
rect 79102 582664 89718 582720
rect 89774 582664 89779 582720
rect 79041 582662 89779 582664
rect 79041 582659 79107 582662
rect 89713 582659 89779 582662
rect 88241 582586 88307 582589
rect 104157 582586 104223 582589
rect 88241 582584 104223 582586
rect 88241 582528 88246 582584
rect 88302 582528 104162 582584
rect 104218 582528 104223 582584
rect 88241 582526 104223 582528
rect 88241 582523 88307 582526
rect 104157 582523 104223 582526
rect 69473 582450 69539 582453
rect 70209 582450 70275 582453
rect 69473 582448 70275 582450
rect 69473 582392 69478 582448
rect 69534 582392 70214 582448
rect 70270 582392 70275 582448
rect 69473 582390 70275 582392
rect 69473 582387 69539 582390
rect 70209 582387 70275 582390
rect 92105 582450 92171 582453
rect 122833 582450 122899 582453
rect 582741 582450 582807 582453
rect 92105 582448 582807 582450
rect 92105 582392 92110 582448
rect 92166 582392 122838 582448
rect 122894 582392 582746 582448
rect 582802 582392 582807 582448
rect 92105 582390 582807 582392
rect 92105 582387 92171 582390
rect 122833 582387 122899 582390
rect 582741 582387 582807 582390
rect 89713 581634 89779 581637
rect 102777 581634 102843 581637
rect 89713 581632 102843 581634
rect 89713 581576 89718 581632
rect 89774 581576 102782 581632
rect 102838 581576 102843 581632
rect 89713 581574 102843 581576
rect 89713 581571 89779 581574
rect 102777 581571 102843 581574
rect 82997 581226 83063 581229
rect 64830 581224 83063 581226
rect 64830 581168 83002 581224
rect 83058 581168 83063 581224
rect 64830 581166 83063 581168
rect 59261 581090 59327 581093
rect 64830 581090 64890 581166
rect 82997 581163 83063 581166
rect 59261 581088 64890 581090
rect 59261 581032 59266 581088
rect 59322 581032 64890 581088
rect 59261 581030 64890 581032
rect 75361 581090 75427 581093
rect 75678 581090 75684 581092
rect 75361 581088 75684 581090
rect 75361 581032 75366 581088
rect 75422 581032 75684 581088
rect 75361 581030 75684 581032
rect 59261 581027 59327 581030
rect 75361 581027 75427 581030
rect 75678 581028 75684 581030
rect 75748 581028 75754 581092
rect 78121 581090 78187 581093
rect 78438 581090 78444 581092
rect 78121 581088 78444 581090
rect 78121 581032 78126 581088
rect 78182 581032 78444 581088
rect 78121 581030 78444 581032
rect 78121 581027 78187 581030
rect 78438 581028 78444 581030
rect 78508 581028 78514 581092
rect 70945 580820 71011 580821
rect 70894 580818 70900 580820
rect 70854 580758 70900 580818
rect 70964 580816 71011 580820
rect 71006 580760 71011 580816
rect 70894 580756 70900 580758
rect 70964 580756 71011 580760
rect 83958 580756 83964 580820
rect 84028 580818 84034 580820
rect 84193 580818 84259 580821
rect 84028 580816 84259 580818
rect 84028 580760 84198 580816
rect 84254 580760 84259 580816
rect 84028 580758 84259 580760
rect 84028 580756 84034 580758
rect 70945 580755 71011 580756
rect 84193 580755 84259 580758
rect 88374 580756 88380 580820
rect 88444 580818 88450 580820
rect 88701 580818 88767 580821
rect 88444 580816 88767 580818
rect 88444 580760 88706 580816
rect 88762 580760 88767 580816
rect 88444 580758 88767 580760
rect 88444 580756 88450 580758
rect 88701 580755 88767 580758
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 66529 580002 66595 580005
rect 68878 580002 68938 580584
rect 66529 580000 68938 580002
rect 66529 579944 66534 580000
rect 66590 579944 68938 580000
rect 66529 579942 68938 579944
rect 66529 579939 66595 579942
rect 53741 578914 53807 578917
rect 68645 578914 68711 578917
rect 53741 578912 68711 578914
rect 53741 578856 53746 578912
rect 53802 578856 68650 578912
rect 68706 578856 68711 578912
rect 53741 578854 68711 578856
rect 53741 578851 53807 578854
rect 68645 578851 68711 578854
rect 66897 578642 66963 578645
rect 68878 578642 68938 579224
rect 94638 578778 94698 579496
rect 94638 578718 103530 578778
rect 66897 578640 68938 578642
rect 66897 578584 66902 578640
rect 66958 578584 68938 578640
rect 66897 578582 68938 578584
rect 66897 578579 66963 578582
rect 103470 578370 103530 578718
rect 130326 578370 130332 578372
rect 103470 578310 130332 578370
rect 130326 578308 130332 578310
rect 130396 578308 130402 578372
rect 67541 577282 67607 577285
rect 68878 577282 68938 577864
rect 94638 577554 94698 578136
rect 582557 577690 582623 577693
rect 583520 577690 584960 577780
rect 582557 577688 584960 577690
rect 582557 577632 582562 577688
rect 582618 577632 584960 577688
rect 582557 577630 584960 577632
rect 582557 577627 582623 577630
rect 97533 577554 97599 577557
rect 94638 577552 97599 577554
rect 94638 577496 97538 577552
rect 97594 577496 97599 577552
rect 583520 577540 584960 577630
rect 94638 577494 97599 577496
rect 97533 577491 97599 577494
rect 67541 577280 68938 577282
rect 67541 577224 67546 577280
rect 67602 577224 68938 577280
rect 67541 577222 68938 577224
rect 67541 577219 67607 577222
rect 94638 576738 94698 576776
rect 97901 576738 97967 576741
rect 94638 576736 97967 576738
rect 94638 576680 97906 576736
rect 97962 576680 97967 576736
rect 94638 576678 97967 576680
rect 97901 576675 97967 576678
rect 66437 575922 66503 575925
rect 68878 575922 68938 576504
rect 66437 575920 68938 575922
rect 66437 575864 66442 575920
rect 66498 575864 68938 575920
rect 66437 575862 68938 575864
rect 66437 575859 66503 575862
rect 67725 575378 67791 575381
rect 94638 575378 94698 575416
rect 95325 575378 95391 575381
rect 97625 575378 97691 575381
rect 67725 575376 68938 575378
rect 67725 575320 67730 575376
rect 67786 575320 68938 575376
rect 67725 575318 68938 575320
rect 94638 575376 97691 575378
rect 94638 575320 95330 575376
rect 95386 575320 97630 575376
rect 97686 575320 97691 575376
rect 94638 575318 97691 575320
rect 67725 575315 67791 575318
rect 68878 575144 68938 575318
rect 95325 575315 95391 575318
rect 97625 575315 97691 575318
rect 66621 573202 66687 573205
rect 68878 573202 68938 573784
rect 94638 573474 94698 574056
rect 97441 573474 97507 573477
rect 94638 573472 97507 573474
rect 94638 573416 97446 573472
rect 97502 573416 97507 573472
rect 94638 573414 97507 573416
rect 97441 573411 97507 573414
rect 66621 573200 68938 573202
rect 66621 573144 66626 573200
rect 66682 573144 68938 573200
rect 66621 573142 68938 573144
rect 66621 573139 66687 573142
rect 94638 572658 94698 572696
rect 99281 572658 99347 572661
rect 94638 572656 99347 572658
rect 94638 572600 99286 572656
rect 99342 572600 99347 572656
rect 94638 572598 99347 572600
rect 99281 572595 99347 572598
rect 66713 571842 66779 571845
rect 68878 571842 68938 572424
rect 66713 571840 68938 571842
rect 66713 571784 66718 571840
rect 66774 571784 68938 571840
rect 66713 571782 68938 571784
rect 66713 571779 66779 571782
rect 97073 571434 97139 571437
rect 94638 571432 97139 571434
rect 94638 571376 97078 571432
rect 97134 571376 97139 571432
rect 94638 571374 97139 571376
rect 94638 571336 94698 571374
rect 97073 571371 97139 571374
rect 66989 570210 67055 570213
rect 68878 570210 68938 570792
rect 97901 570346 97967 570349
rect 66989 570208 68938 570210
rect 66989 570152 66994 570208
rect 67050 570152 68938 570208
rect 66989 570150 68938 570152
rect 94638 570344 97967 570346
rect 94638 570288 97906 570344
rect 97962 570288 97967 570344
rect 94638 570286 97967 570288
rect 66989 570147 67055 570150
rect 94638 569976 94698 570286
rect 97901 570283 97967 570286
rect 67725 568850 67791 568853
rect 68878 568850 68938 569432
rect 96797 569122 96863 569125
rect 97901 569122 97967 569125
rect 67725 568848 68938 568850
rect 67725 568792 67730 568848
rect 67786 568792 68938 568848
rect 67725 568790 68938 568792
rect 94638 569120 97967 569122
rect 94638 569064 96802 569120
rect 96858 569064 97906 569120
rect 97962 569064 97967 569120
rect 94638 569062 97967 569064
rect 67725 568787 67791 568790
rect 94638 568616 94698 569062
rect 96797 569059 96863 569062
rect 97901 569059 97967 569062
rect 66069 567626 66135 567629
rect 68878 567626 68938 568072
rect 66069 567624 68938 567626
rect 66069 567568 66074 567624
rect 66130 567568 68938 567624
rect 66069 567566 68938 567568
rect 66069 567563 66135 567566
rect 94638 567218 94698 567256
rect 95417 567218 95483 567221
rect 94638 567216 95483 567218
rect 94638 567160 95422 567216
rect 95478 567160 95483 567216
rect 94638 567158 95483 567160
rect 95417 567155 95483 567158
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 67633 566674 67699 566677
rect 68878 566674 68938 566712
rect 67633 566672 68938 566674
rect 67633 566616 67638 566672
rect 67694 566616 68938 566672
rect 67633 566614 68938 566616
rect 67633 566611 67699 566614
rect 94638 565858 94698 565896
rect 97901 565858 97967 565861
rect 94638 565856 97967 565858
rect 94638 565800 97906 565856
rect 97962 565800 97967 565856
rect 94638 565798 97967 565800
rect 97901 565795 97967 565798
rect 66805 564770 66871 564773
rect 68878 564770 68938 565352
rect 66805 564768 68938 564770
rect 66805 564712 66810 564768
rect 66866 564712 68938 564768
rect 66805 564710 68938 564712
rect 66805 564707 66871 564710
rect 582741 564362 582807 564365
rect 583520 564362 584960 564452
rect 582741 564360 584960 564362
rect 582741 564304 582746 564360
rect 582802 564304 584960 564360
rect 582741 564302 584960 564304
rect 582741 564299 582807 564302
rect 66529 564226 66595 564229
rect 66529 564224 68938 564226
rect 66529 564168 66534 564224
rect 66590 564168 68938 564224
rect 66529 564166 68938 564168
rect 66529 564163 66595 564166
rect 68878 563992 68938 564166
rect 94638 563682 94698 564264
rect 583520 564212 584960 564302
rect 95233 563682 95299 563685
rect 94638 563680 95299 563682
rect 94638 563624 95238 563680
rect 95294 563624 95299 563680
rect 94638 563622 95299 563624
rect 95233 563619 95299 563622
rect 66805 562050 66871 562053
rect 68878 562050 68938 562632
rect 94638 562322 94698 562904
rect 96797 562322 96863 562325
rect 94638 562320 96863 562322
rect 94638 562264 96802 562320
rect 96858 562264 96863 562320
rect 94638 562262 96863 562264
rect 96797 562259 96863 562262
rect 66805 562048 68938 562050
rect 66805 561992 66810 562048
rect 66866 561992 68938 562048
rect 66805 561990 68938 561992
rect 66805 561987 66871 561990
rect 66805 560690 66871 560693
rect 68878 560690 68938 561272
rect 94638 560962 94698 561544
rect 96889 560962 96955 560965
rect 94638 560960 96955 560962
rect 94638 560904 96894 560960
rect 96950 560904 96955 560960
rect 94638 560902 96955 560904
rect 96889 560899 96955 560902
rect 66805 560688 68938 560690
rect 66805 560632 66810 560688
rect 66866 560632 68938 560688
rect 66805 560630 68938 560632
rect 66805 560627 66871 560630
rect 66805 559330 66871 559333
rect 68878 559330 68938 559912
rect 94638 559602 94698 560184
rect 96797 559602 96863 559605
rect 94638 559600 96863 559602
rect 94638 559544 96802 559600
rect 96858 559544 96863 559600
rect 94638 559542 96863 559544
rect 96797 559539 96863 559542
rect 66805 559328 68938 559330
rect 66805 559272 66810 559328
rect 66866 559272 68938 559328
rect 66805 559270 68938 559272
rect 66805 559267 66871 559270
rect 94638 558786 94698 558824
rect 96705 558786 96771 558789
rect 97165 558786 97231 558789
rect 94638 558784 97231 558786
rect 94638 558728 96710 558784
rect 96766 558728 97170 558784
rect 97226 558728 97231 558784
rect 94638 558726 97231 558728
rect 96705 558723 96771 558726
rect 97165 558723 97231 558726
rect 66805 557970 66871 557973
rect 68878 557970 68938 558552
rect 66805 557968 68938 557970
rect 66805 557912 66810 557968
rect 66866 557912 68938 557968
rect 66805 557910 68938 557912
rect 66805 557907 66871 557910
rect 67633 556610 67699 556613
rect 68878 556610 68938 557192
rect 94638 556882 94698 557464
rect 96797 556882 96863 556885
rect 94638 556880 96863 556882
rect 94638 556824 96802 556880
rect 96858 556824 96863 556880
rect 94638 556822 96863 556824
rect 96797 556819 96863 556822
rect 67633 556608 68938 556610
rect 67633 556552 67638 556608
rect 67694 556552 68938 556608
rect 67633 556550 68938 556552
rect 67633 556547 67699 556550
rect 66713 555250 66779 555253
rect 68878 555250 68938 555832
rect 94638 555522 94698 556104
rect 94773 555522 94839 555525
rect 94638 555520 94839 555522
rect 94638 555464 94778 555520
rect 94834 555464 94839 555520
rect 94638 555462 94839 555464
rect 94773 555459 94839 555462
rect 66713 555248 68938 555250
rect 66713 555192 66718 555248
rect 66774 555192 68938 555248
rect 66713 555190 68938 555192
rect 66713 555187 66779 555190
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 66805 553618 66871 553621
rect 68878 553618 68938 554200
rect 94638 554162 94698 554744
rect 97206 554162 97212 554164
rect 94638 554102 97212 554162
rect 97206 554100 97212 554102
rect 97276 554100 97282 554164
rect 66805 553616 68938 553618
rect 66805 553560 66810 553616
rect 66866 553560 68938 553616
rect 66805 553558 68938 553560
rect 66805 553555 66871 553558
rect 67449 552258 67515 552261
rect 68878 552258 68938 552840
rect 94638 552802 94698 553384
rect 96981 552802 97047 552805
rect 94638 552800 97047 552802
rect 94638 552744 96986 552800
rect 97042 552744 97047 552800
rect 94638 552742 97047 552744
rect 96981 552739 97047 552742
rect 95509 552530 95575 552533
rect 96613 552530 96679 552533
rect 67449 552256 68938 552258
rect 67449 552200 67454 552256
rect 67510 552200 68938 552256
rect 67449 552198 68938 552200
rect 94638 552528 96679 552530
rect 94638 552472 95514 552528
rect 95570 552472 96618 552528
rect 96674 552472 96679 552528
rect 94638 552470 96679 552472
rect 67449 552195 67515 552198
rect 94638 552024 94698 552470
rect 95509 552467 95575 552470
rect 96613 552467 96679 552470
rect 67817 550898 67883 550901
rect 68878 550898 68938 551480
rect 583520 551020 584960 551260
rect 67817 550896 68938 550898
rect 67817 550840 67822 550896
rect 67878 550840 68938 550896
rect 67817 550838 68938 550840
rect 67817 550835 67883 550838
rect 97901 550762 97967 550765
rect 94638 550760 97967 550762
rect 94638 550704 97906 550760
rect 97962 550704 97967 550760
rect 94638 550702 97967 550704
rect 94638 550664 94698 550702
rect 97901 550699 97967 550702
rect 66805 549538 66871 549541
rect 68878 549538 68938 550120
rect 66805 549536 68938 549538
rect 66805 549480 66810 549536
rect 66866 549480 68938 549536
rect 66805 549478 68938 549480
rect 66805 549475 66871 549478
rect 97073 549402 97139 549405
rect 94638 549400 97139 549402
rect 94638 549344 97078 549400
rect 97134 549344 97139 549400
rect 94638 549342 97139 549344
rect 94638 549304 94698 549342
rect 97073 549339 97139 549342
rect 67766 548252 67772 548316
rect 67836 548314 67842 548316
rect 68878 548314 68938 548760
rect 67836 548254 68938 548314
rect 67836 548252 67842 548254
rect 100017 547906 100083 547909
rect 104934 547906 104940 547908
rect 100017 547904 104940 547906
rect 100017 547848 100022 547904
rect 100078 547848 104940 547904
rect 100017 547846 104940 547848
rect 100017 547843 100083 547846
rect 104934 547844 104940 547846
rect 105004 547844 105010 547908
rect 66529 546818 66595 546821
rect 68878 546818 68938 547400
rect 94638 547090 94698 547672
rect 96654 547090 96660 547092
rect 94638 547030 96660 547090
rect 96654 547028 96660 547030
rect 96724 547028 96730 547092
rect 66529 546816 68938 546818
rect 66529 546760 66534 546816
rect 66590 546760 68938 546816
rect 66529 546758 68938 546760
rect 66529 546755 66595 546758
rect 66253 546002 66319 546005
rect 68878 546002 68938 546040
rect 66253 546000 68938 546002
rect 66253 545944 66258 546000
rect 66314 545944 68938 546000
rect 66253 545942 68938 545944
rect 66253 545939 66319 545942
rect 94638 545730 94698 546312
rect 96981 545730 97047 545733
rect 94638 545728 97047 545730
rect 94638 545672 96986 545728
rect 97042 545672 97047 545728
rect 94638 545670 97047 545672
rect 96981 545667 97047 545670
rect 66345 544506 66411 544509
rect 68878 544506 68938 544680
rect 66345 544504 68938 544506
rect 66345 544448 66350 544504
rect 66406 544448 68938 544504
rect 66345 544446 68938 544448
rect 66345 544443 66411 544446
rect 94638 544370 94698 544952
rect 97349 544370 97415 544373
rect 94638 544368 97415 544370
rect 94638 544312 97354 544368
rect 97410 544312 97415 544368
rect 94638 544310 97415 544312
rect 97349 544307 97415 544310
rect 66621 543146 66687 543149
rect 68878 543146 68938 543320
rect 66621 543144 68938 543146
rect 66621 543088 66626 543144
rect 66682 543088 68938 543144
rect 66621 543086 68938 543088
rect 66621 543083 66687 543086
rect 94638 543010 94698 543592
rect 96705 543010 96771 543013
rect 94638 543008 96771 543010
rect 94638 542952 96710 543008
rect 96766 542952 96771 543008
rect 94638 542950 96771 542952
rect 96705 542947 96771 542950
rect 69422 542132 69428 542196
rect 69492 542132 69498 542196
rect 4797 541106 4863 541109
rect 69430 541106 69490 542132
rect 94086 541652 94146 542232
rect 94078 541588 94084 541652
rect 94148 541588 94154 541652
rect 4797 541104 69490 541106
rect 4797 541048 4802 541104
rect 4858 541048 69490 541104
rect 4797 541046 69490 541048
rect 4797 541043 4863 541046
rect -960 540684 480 540924
rect 66621 540018 66687 540021
rect 68878 540018 68938 540600
rect 66621 540016 68938 540018
rect 66621 539960 66626 540016
rect 66682 539960 68938 540016
rect 66621 539958 68938 539960
rect 66621 539955 66687 539958
rect 67766 539820 67772 539884
rect 67836 539882 67842 539884
rect 69105 539882 69171 539885
rect 67836 539880 69171 539882
rect 67836 539824 69110 539880
rect 69166 539824 69171 539880
rect 67836 539822 69171 539824
rect 67836 539820 67842 539822
rect 69105 539819 69171 539822
rect 93853 539882 93919 539885
rect 94086 539882 94146 540872
rect 93853 539880 94146 539882
rect 93853 539824 93858 539880
rect 93914 539824 94146 539880
rect 93853 539822 94146 539824
rect 93853 539819 93919 539822
rect 94638 538930 94698 539512
rect 96613 538930 96679 538933
rect 94638 538928 96679 538930
rect 94638 538872 96618 538928
rect 96674 538872 96679 538928
rect 94638 538870 96679 538872
rect 96613 538867 96679 538870
rect 91502 538188 91508 538252
rect 91572 538250 91578 538252
rect 94681 538250 94747 538253
rect 91572 538248 94747 538250
rect 91572 538192 94686 538248
rect 94742 538192 94747 538248
rect 91572 538190 94747 538192
rect 91572 538188 91578 538190
rect 94681 538187 94747 538190
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 76465 536754 76531 536757
rect 116577 536754 116643 536757
rect 76465 536752 116643 536754
rect 76465 536696 76470 536752
rect 76526 536696 116582 536752
rect 116638 536696 116643 536752
rect 76465 536694 116643 536696
rect 76465 536691 76531 536694
rect 116577 536691 116643 536694
rect 76465 535666 76531 535669
rect 77201 535666 77267 535669
rect 76465 535664 77267 535666
rect 76465 535608 76470 535664
rect 76526 535608 77206 535664
rect 77262 535608 77267 535664
rect 76465 535606 77267 535608
rect 76465 535603 76531 535606
rect 77201 535603 77267 535606
rect 75913 535532 75979 535533
rect 75862 535530 75868 535532
rect 75786 535470 75868 535530
rect 75932 535530 75979 535532
rect 76741 535530 76807 535533
rect 75932 535528 76807 535530
rect 75974 535472 76746 535528
rect 76802 535472 76807 535528
rect 75862 535468 75868 535470
rect 75932 535470 76807 535472
rect 75932 535468 75979 535470
rect 75913 535467 75979 535468
rect 76741 535467 76807 535470
rect 58985 533354 59051 533357
rect 96654 533354 96660 533356
rect 58985 533352 96660 533354
rect 58985 533296 58990 533352
rect 59046 533296 96660 533352
rect 58985 533294 96660 533296
rect 58985 533291 59051 533294
rect 96654 533292 96660 533294
rect 96724 533292 96730 533356
rect 37089 531994 37155 531997
rect 94078 531994 94084 531996
rect 37089 531992 94084 531994
rect 37089 531936 37094 531992
rect 37150 531936 94084 531992
rect 37089 531934 94084 531936
rect 37089 531931 37155 531934
rect 94078 531932 94084 531934
rect 94148 531932 94154 531996
rect -960 527914 480 528004
rect 3509 527914 3575 527917
rect -960 527912 3575 527914
rect -960 527856 3514 527912
rect 3570 527856 3575 527912
rect -960 527854 3575 527856
rect -960 527764 480 527854
rect 3509 527851 3575 527854
rect 79910 527716 79916 527780
rect 79980 527778 79986 527780
rect 95417 527778 95483 527781
rect 79980 527776 95483 527778
rect 79980 527720 95422 527776
rect 95478 527720 95483 527776
rect 79980 527718 95483 527720
rect 79980 527716 79986 527718
rect 95417 527715 95483 527718
rect 582649 524514 582715 524517
rect 583520 524514 584960 524604
rect 582649 524512 584960 524514
rect 582649 524456 582654 524512
rect 582710 524456 584960 524512
rect 582649 524454 584960 524456
rect 582649 524451 582715 524454
rect 583520 524364 584960 524454
rect 81341 520978 81407 520981
rect 94446 520978 94452 520980
rect 81341 520976 94452 520978
rect 81341 520920 81346 520976
rect 81402 520920 94452 520976
rect 81341 520918 94452 520920
rect 81341 520915 81407 520918
rect 94446 520916 94452 520918
rect 94516 520916 94522 520980
rect 77150 518060 77156 518124
rect 77220 518122 77226 518124
rect 94773 518122 94839 518125
rect 77220 518120 94839 518122
rect 77220 518064 94778 518120
rect 94834 518064 94839 518120
rect 77220 518062 94839 518064
rect 77220 518060 77226 518062
rect 94773 518059 94839 518062
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 100109 507922 100175 507925
rect 100702 507922 100708 507924
rect 100109 507920 100708 507922
rect 100109 507864 100114 507920
rect 100170 507864 100708 507920
rect 100109 507862 100708 507864
rect 100109 507859 100175 507862
rect 100702 507860 100708 507862
rect 100772 507860 100778 507924
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 582741 484666 582807 484669
rect 583520 484666 584960 484756
rect 582741 484664 584960 484666
rect 582741 484608 582746 484664
rect 582802 484608 584960 484664
rect 582741 484606 584960 484608
rect 582741 484603 582807 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 2957 475690 3023 475693
rect -960 475688 3023 475690
rect -960 475632 2962 475688
rect 3018 475632 3023 475688
rect -960 475630 3023 475632
rect -960 475540 480 475630
rect 2957 475627 3023 475630
rect 582833 471474 582899 471477
rect 583520 471474 584960 471564
rect 582833 471472 584960 471474
rect 582833 471416 582838 471472
rect 582894 471416 584960 471472
rect 582833 471414 584960 471416
rect 582833 471411 582899 471414
rect 583520 471324 584960 471414
rect 75678 468420 75684 468484
rect 75748 468482 75754 468484
rect 90449 468482 90515 468485
rect 75748 468480 90515 468482
rect 75748 468424 90454 468480
rect 90510 468424 90515 468480
rect 75748 468422 90515 468424
rect 75748 468420 75754 468422
rect 90449 468419 90515 468422
rect 88425 463042 88491 463045
rect 106406 463042 106412 463044
rect 88425 463040 106412 463042
rect 88425 462984 88430 463040
rect 88486 462984 106412 463040
rect 88425 462982 106412 462984
rect 88425 462979 88491 462982
rect 106406 462980 106412 462982
rect 106476 462980 106482 463044
rect 69606 462844 69612 462908
rect 69676 462906 69682 462908
rect 88742 462906 88748 462908
rect 69676 462846 88748 462906
rect 69676 462844 69682 462846
rect 88742 462844 88748 462846
rect 88812 462844 88818 462908
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 69606 461484 69612 461548
rect 69676 461546 69682 461548
rect 96981 461546 97047 461549
rect 69676 461544 97047 461546
rect 69676 461488 96986 461544
rect 97042 461488 97047 461544
rect 69676 461486 97047 461488
rect 69676 461484 69682 461486
rect 96981 461483 97047 461486
rect 78438 460124 78444 460188
rect 78508 460186 78514 460188
rect 92606 460186 92612 460188
rect 78508 460126 92612 460186
rect 78508 460124 78514 460126
rect 92606 460124 92612 460126
rect 92676 460124 92682 460188
rect 106917 458826 106983 458829
rect 114502 458826 114508 458828
rect 106917 458824 114508 458826
rect 106917 458768 106922 458824
rect 106978 458768 114508 458824
rect 106917 458766 114508 458768
rect 106917 458763 106983 458766
rect 114502 458764 114508 458766
rect 114572 458764 114578 458828
rect 582373 458146 582439 458149
rect 583520 458146 584960 458236
rect 582373 458144 584960 458146
rect 582373 458088 582378 458144
rect 582434 458088 584960 458144
rect 582373 458086 584960 458088
rect 582373 458083 582439 458086
rect 583520 457996 584960 458086
rect 72550 454684 72556 454748
rect 72620 454746 72626 454748
rect 95233 454746 95299 454749
rect 72620 454744 95299 454746
rect 72620 454688 95238 454744
rect 95294 454688 95299 454744
rect 72620 454686 95299 454688
rect 72620 454684 72626 454686
rect 95233 454683 95299 454686
rect 80053 453250 80119 453253
rect 113214 453250 113220 453252
rect 80053 453248 113220 453250
rect 80053 453192 80058 453248
rect 80114 453192 113220 453248
rect 80053 453190 113220 453192
rect 80053 453187 80119 453190
rect 113214 453188 113220 453190
rect 113284 453188 113290 453252
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 86217 449170 86283 449173
rect 107694 449170 107700 449172
rect 86217 449168 107700 449170
rect 86217 449112 86222 449168
rect 86278 449112 107700 449168
rect 86217 449110 107700 449112
rect 86217 449107 86283 449110
rect 107694 449108 107700 449110
rect 107764 449108 107770 449172
rect 101397 446450 101463 446453
rect 123334 446450 123340 446452
rect 101397 446448 123340 446450
rect 101397 446392 101402 446448
rect 101458 446392 123340 446448
rect 101397 446390 123340 446392
rect 101397 446387 101463 446390
rect 123334 446388 123340 446390
rect 123404 446388 123410 446452
rect 81341 444954 81407 444957
rect 88374 444954 88380 444956
rect 81341 444952 88380 444954
rect 81341 444896 81346 444952
rect 81402 444896 88380 444952
rect 81341 444894 88380 444896
rect 81341 444891 81407 444894
rect 88374 444892 88380 444894
rect 88444 444892 88450 444956
rect 583520 444668 584960 444908
rect 96613 444274 96679 444277
rect 97206 444274 97212 444276
rect 96613 444272 97212 444274
rect 96613 444216 96618 444272
rect 96674 444216 97212 444272
rect 96613 444214 97212 444216
rect 96613 444211 96679 444214
rect 97206 444212 97212 444214
rect 97276 444212 97282 444276
rect 66110 443532 66116 443596
rect 66180 443594 66186 443596
rect 83457 443594 83523 443597
rect 66180 443592 83523 443594
rect 66180 443536 83462 443592
rect 83518 443536 83523 443592
rect 66180 443534 83523 443536
rect 66180 443532 66186 443534
rect 83457 443531 83523 443534
rect 96613 443050 96679 443053
rect 117313 443050 117379 443053
rect 96613 443048 117379 443050
rect 96613 442992 96618 443048
rect 96674 442992 117318 443048
rect 117374 442992 117379 443048
rect 96613 442990 117379 442992
rect 96613 442987 96679 442990
rect 117313 442987 117379 442990
rect 88333 441010 88399 441013
rect 113265 441010 113331 441013
rect 88333 441008 113331 441010
rect 88333 440952 88338 441008
rect 88394 440952 113270 441008
rect 113326 440952 113331 441008
rect 88333 440950 113331 440952
rect 88333 440947 88399 440950
rect 113265 440947 113331 440950
rect 98637 439514 98703 439517
rect 117497 439514 117563 439517
rect 98637 439512 117563 439514
rect 98637 439456 98642 439512
rect 98698 439456 117502 439512
rect 117558 439456 117563 439512
rect 98637 439454 117563 439456
rect 98637 439451 98703 439454
rect 117497 439451 117563 439454
rect 85757 437610 85823 437613
rect 86861 437610 86927 437613
rect 120073 437610 120139 437613
rect 85757 437608 120139 437610
rect 85757 437552 85762 437608
rect 85818 437552 86866 437608
rect 86922 437552 120078 437608
rect 120134 437552 120139 437608
rect 85757 437550 120139 437552
rect 85757 437547 85823 437550
rect 86861 437547 86927 437550
rect 120073 437547 120139 437550
rect -960 436508 480 436748
rect 106733 436386 106799 436389
rect 103286 436384 106799 436386
rect 103286 436328 106738 436384
rect 106794 436328 106799 436384
rect 103286 436326 106799 436328
rect 52177 436250 52243 436253
rect 68461 436250 68527 436253
rect 52177 436248 68527 436250
rect 52177 436192 52182 436248
rect 52238 436192 68466 436248
rect 68522 436192 68527 436248
rect 52177 436190 68527 436192
rect 52177 436187 52243 436190
rect 68461 436187 68527 436190
rect 72734 436188 72740 436252
rect 72804 436250 72810 436252
rect 77385 436250 77451 436253
rect 72804 436248 77451 436250
rect 72804 436192 77390 436248
rect 77446 436192 77451 436248
rect 72804 436190 77451 436192
rect 72804 436188 72810 436190
rect 77385 436187 77451 436190
rect 86166 436188 86172 436252
rect 86236 436250 86242 436252
rect 91093 436250 91159 436253
rect 103286 436252 103346 436326
rect 106733 436323 106799 436326
rect 86236 436248 91159 436250
rect 86236 436192 91098 436248
rect 91154 436192 91159 436248
rect 86236 436190 91159 436192
rect 86236 436188 86242 436190
rect 91093 436187 91159 436190
rect 103278 436188 103284 436252
rect 103348 436188 103354 436252
rect 109125 436250 109191 436253
rect 103470 436248 109191 436250
rect 103470 436192 109130 436248
rect 109186 436192 109191 436248
rect 103470 436190 109191 436192
rect 78254 436052 78260 436116
rect 78324 436114 78330 436116
rect 83181 436114 83247 436117
rect 78324 436112 83247 436114
rect 78324 436056 83186 436112
rect 83242 436056 83247 436112
rect 78324 436054 83247 436056
rect 78324 436052 78330 436054
rect 83181 436051 83247 436054
rect 87321 436114 87387 436117
rect 88241 436114 88307 436117
rect 87321 436112 88307 436114
rect 87321 436056 87326 436112
rect 87382 436056 88246 436112
rect 88302 436056 88307 436112
rect 87321 436054 88307 436056
rect 87321 436051 87387 436054
rect 88241 436051 88307 436054
rect 100518 436052 100524 436116
rect 100588 436114 100594 436116
rect 103470 436114 103530 436190
rect 109125 436187 109191 436190
rect 100588 436054 103530 436114
rect 107653 436114 107719 436117
rect 108205 436114 108271 436117
rect 107653 436112 108271 436114
rect 107653 436056 107658 436112
rect 107714 436056 108210 436112
rect 108266 436056 108271 436112
rect 107653 436054 108271 436056
rect 100588 436052 100594 436054
rect 107653 436051 107719 436054
rect 108205 436051 108271 436054
rect 110413 436114 110479 436117
rect 110965 436114 111031 436117
rect 110413 436112 111031 436114
rect 110413 436056 110418 436112
rect 110474 436056 110970 436112
rect 111026 436056 111031 436112
rect 110413 436054 111031 436056
rect 110413 436051 110479 436054
rect 110965 436051 111031 436054
rect 82118 435916 82124 435980
rect 82188 435978 82194 435980
rect 83958 435978 83964 435980
rect 82188 435918 83964 435978
rect 82188 435916 82194 435918
rect 83958 435916 83964 435918
rect 84028 435916 84034 435980
rect 71630 435372 71636 435436
rect 71700 435434 71706 435436
rect 77477 435434 77543 435437
rect 71700 435432 77543 435434
rect 71700 435376 77482 435432
rect 77538 435376 77543 435432
rect 71700 435374 77543 435376
rect 71700 435372 71706 435374
rect 77477 435371 77543 435374
rect 104157 435298 104223 435301
rect 115197 435298 115263 435301
rect 104157 435296 115263 435298
rect 104157 435240 104162 435296
rect 104218 435240 115202 435296
rect 115258 435240 115263 435296
rect 104157 435238 115263 435240
rect 104157 435235 104223 435238
rect 115197 435235 115263 435238
rect 100017 435026 100083 435029
rect 100017 435024 103530 435026
rect 100017 434968 100022 435024
rect 100078 434968 103530 435024
rect 100017 434966 103530 434968
rect 100017 434963 100083 434966
rect 73470 434828 73476 434892
rect 73540 434890 73546 434892
rect 80421 434890 80487 434893
rect 73540 434888 80487 434890
rect 73540 434832 80426 434888
rect 80482 434832 80487 434888
rect 73540 434830 80487 434832
rect 73540 434828 73546 434830
rect 80421 434827 80487 434830
rect 90950 434828 90956 434892
rect 91020 434890 91026 434892
rect 101213 434890 101279 434893
rect 91020 434888 101279 434890
rect 91020 434832 101218 434888
rect 101274 434832 101279 434888
rect 91020 434830 101279 434832
rect 91020 434828 91026 434830
rect 101213 434827 101279 434830
rect 70158 434692 70164 434756
rect 70228 434754 70234 434756
rect 70228 434694 74550 434754
rect 70228 434692 70234 434694
rect 74490 434482 74550 434694
rect 75678 434692 75684 434756
rect 75748 434754 75754 434756
rect 77937 434754 78003 434757
rect 82905 434754 82971 434757
rect 75748 434752 82971 434754
rect 75748 434696 77942 434752
rect 77998 434696 82910 434752
rect 82966 434696 82971 434752
rect 75748 434694 82971 434696
rect 75748 434692 75754 434694
rect 77937 434691 78003 434694
rect 82905 434691 82971 434694
rect 85430 434692 85436 434756
rect 85500 434754 85506 434756
rect 92657 434754 92723 434757
rect 85500 434752 92723 434754
rect 85500 434696 92662 434752
rect 92718 434696 92723 434752
rect 85500 434694 92723 434696
rect 103470 434754 103530 434966
rect 124397 434754 124463 434757
rect 103470 434752 124463 434754
rect 103470 434696 124402 434752
rect 124458 434696 124463 434752
rect 103470 434694 124463 434696
rect 85500 434692 85506 434694
rect 92657 434691 92723 434694
rect 124397 434691 124463 434694
rect 83406 434556 83412 434620
rect 83476 434618 83482 434620
rect 84469 434618 84535 434621
rect 83476 434616 84535 434618
rect 83476 434560 84474 434616
rect 84530 434560 84535 434616
rect 83476 434558 84535 434560
rect 83476 434556 83482 434558
rect 84469 434555 84535 434558
rect 75453 434482 75519 434485
rect 74490 434480 75519 434482
rect 74490 434424 75458 434480
rect 75514 434424 75519 434480
rect 74490 434422 75519 434424
rect 75453 434419 75519 434422
rect 83590 434420 83596 434484
rect 83660 434482 83666 434484
rect 83733 434482 83799 434485
rect 83660 434480 83799 434482
rect 83660 434424 83738 434480
rect 83794 434424 83799 434480
rect 83660 434422 83799 434424
rect 83660 434420 83666 434422
rect 83733 434419 83799 434422
rect 74574 434284 74580 434348
rect 74644 434346 74650 434348
rect 74717 434346 74783 434349
rect 74644 434344 74783 434346
rect 74644 434288 74722 434344
rect 74778 434288 74783 434344
rect 74644 434286 74783 434288
rect 74644 434284 74650 434286
rect 74717 434283 74783 434286
rect 75862 434284 75868 434348
rect 75932 434346 75938 434348
rect 76189 434346 76255 434349
rect 75932 434344 76255 434346
rect 75932 434288 76194 434344
rect 76250 434288 76255 434344
rect 75932 434286 76255 434288
rect 75932 434284 75938 434286
rect 76189 434283 76255 434286
rect 80237 434348 80303 434349
rect 80237 434344 80284 434348
rect 80348 434346 80354 434348
rect 80237 434288 80242 434344
rect 80237 434284 80284 434288
rect 80348 434286 80394 434346
rect 80348 434284 80354 434286
rect 80646 434284 80652 434348
rect 80716 434346 80722 434348
rect 80973 434346 81039 434349
rect 80716 434344 81039 434346
rect 80716 434288 80978 434344
rect 81034 434288 81039 434344
rect 80716 434286 81039 434288
rect 80716 434284 80722 434286
rect 80237 434283 80303 434284
rect 80973 434283 81039 434286
rect 81893 434348 81959 434349
rect 85849 434348 85915 434349
rect 87137 434348 87203 434349
rect 81893 434344 81940 434348
rect 82004 434346 82010 434348
rect 85798 434346 85804 434348
rect 81893 434288 81898 434344
rect 81893 434284 81940 434288
rect 82004 434286 82050 434346
rect 85758 434286 85804 434346
rect 85868 434344 85915 434348
rect 87086 434346 87092 434348
rect 85910 434288 85915 434344
rect 82004 434284 82010 434286
rect 85798 434284 85804 434286
rect 85868 434284 85915 434288
rect 87046 434286 87092 434346
rect 87156 434344 87203 434348
rect 87198 434288 87203 434344
rect 87086 434284 87092 434286
rect 87156 434284 87203 434288
rect 93894 434284 93900 434348
rect 93964 434346 93970 434348
rect 94221 434346 94287 434349
rect 93964 434344 94287 434346
rect 93964 434288 94226 434344
rect 94282 434288 94287 434344
rect 93964 434286 94287 434288
rect 93964 434284 93970 434286
rect 81893 434283 81959 434284
rect 85849 434283 85915 434284
rect 87137 434283 87203 434284
rect 94221 434283 94287 434286
rect 97165 434348 97231 434349
rect 97165 434344 97212 434348
rect 97276 434346 97282 434348
rect 97165 434288 97170 434344
rect 97165 434284 97212 434288
rect 97276 434286 97322 434346
rect 97276 434284 97282 434286
rect 102174 434284 102180 434348
rect 102244 434346 102250 434348
rect 102593 434346 102659 434349
rect 102244 434344 102659 434346
rect 102244 434288 102598 434344
rect 102654 434288 102659 434344
rect 102244 434286 102659 434288
rect 102244 434284 102250 434286
rect 97165 434283 97231 434284
rect 102593 434283 102659 434286
rect 104157 434348 104223 434349
rect 108205 434348 108271 434349
rect 104157 434344 104204 434348
rect 104268 434346 104274 434348
rect 104157 434288 104162 434344
rect 104157 434284 104204 434288
rect 104268 434286 104314 434346
rect 108205 434344 108252 434348
rect 108316 434346 108322 434348
rect 108205 434288 108210 434344
rect 104268 434284 104274 434286
rect 108205 434284 108252 434288
rect 108316 434286 108362 434346
rect 108316 434284 108322 434286
rect 104157 434283 104223 434284
rect 108205 434283 108271 434284
rect 66069 433938 66135 433941
rect 71221 433938 71287 433941
rect 66069 433936 71287 433938
rect 66069 433880 66074 433936
rect 66130 433880 71226 433936
rect 71282 433880 71287 433936
rect 66069 433878 71287 433880
rect 66069 433875 66135 433878
rect 71221 433875 71287 433878
rect 97390 433876 97396 433940
rect 97460 433938 97466 433940
rect 100569 433938 100635 433941
rect 97460 433936 100635 433938
rect 97460 433880 100574 433936
rect 100630 433880 100635 433936
rect 97460 433878 100635 433880
rect 97460 433876 97466 433878
rect 100569 433875 100635 433878
rect 109166 433876 109172 433940
rect 109236 433938 109242 433940
rect 109585 433938 109651 433941
rect 109236 433936 109651 433938
rect 109236 433880 109590 433936
rect 109646 433880 109651 433936
rect 109236 433878 109651 433880
rect 109236 433876 109242 433878
rect 109585 433875 109651 433878
rect 70853 433804 70919 433805
rect 70853 433802 70900 433804
rect 70808 433800 70900 433802
rect 70808 433744 70858 433800
rect 70808 433742 70900 433744
rect 70853 433740 70900 433742
rect 70964 433740 70970 433804
rect 84694 433740 84700 433804
rect 84764 433802 84770 433804
rect 87965 433802 88031 433805
rect 84764 433800 88031 433802
rect 84764 433744 87970 433800
rect 88026 433744 88031 433800
rect 84764 433742 88031 433744
rect 84764 433740 84770 433742
rect 70853 433739 70919 433740
rect 87965 433739 88031 433742
rect 98126 433740 98132 433804
rect 98196 433802 98202 433804
rect 98453 433802 98519 433805
rect 98196 433800 98519 433802
rect 98196 433744 98458 433800
rect 98514 433744 98519 433800
rect 98196 433742 98519 433744
rect 98196 433740 98202 433742
rect 98453 433739 98519 433742
rect 101990 433740 101996 433804
rect 102060 433802 102066 433804
rect 102060 433742 112178 433802
rect 102060 433740 102066 433742
rect 53557 433666 53623 433669
rect 73429 433666 73495 433669
rect 53557 433664 73495 433666
rect 53557 433608 53562 433664
rect 53618 433608 73434 433664
rect 73490 433608 73495 433664
rect 53557 433606 73495 433608
rect 53557 433603 53623 433606
rect 73429 433603 73495 433606
rect 78397 433668 78463 433669
rect 78397 433664 78444 433668
rect 78508 433666 78514 433668
rect 79593 433666 79659 433669
rect 87321 433668 87387 433669
rect 79726 433666 79732 433668
rect 78397 433608 78402 433664
rect 78397 433604 78444 433608
rect 78508 433606 78554 433666
rect 79593 433664 79732 433666
rect 79593 433608 79598 433664
rect 79654 433608 79732 433664
rect 79593 433606 79732 433608
rect 78508 433604 78514 433606
rect 78397 433603 78463 433604
rect 79593 433603 79659 433606
rect 79726 433604 79732 433606
rect 79796 433604 79802 433668
rect 87270 433666 87276 433668
rect 87230 433606 87276 433666
rect 87340 433664 87387 433668
rect 87382 433608 87387 433664
rect 87270 433604 87276 433606
rect 87340 433604 87387 433608
rect 89662 433604 89668 433668
rect 89732 433666 89738 433668
rect 89989 433666 90055 433669
rect 89732 433664 90055 433666
rect 89732 433608 89994 433664
rect 90050 433608 90055 433664
rect 89732 433606 90055 433608
rect 89732 433604 89738 433606
rect 87321 433603 87387 433604
rect 89989 433603 90055 433606
rect 91318 433604 91324 433668
rect 91388 433666 91394 433668
rect 91461 433666 91527 433669
rect 91388 433664 91527 433666
rect 91388 433608 91466 433664
rect 91522 433608 91527 433664
rect 91388 433606 91527 433608
rect 91388 433604 91394 433606
rect 91461 433603 91527 433606
rect 93485 433666 93551 433669
rect 95141 433668 95207 433669
rect 93710 433666 93716 433668
rect 93485 433664 93716 433666
rect 93485 433608 93490 433664
rect 93546 433608 93716 433664
rect 93485 433606 93716 433608
rect 93485 433603 93551 433606
rect 93710 433604 93716 433606
rect 93780 433604 93786 433668
rect 95141 433664 95188 433668
rect 95252 433666 95258 433668
rect 98361 433666 98427 433669
rect 98494 433666 98500 433668
rect 95141 433608 95146 433664
rect 95141 433604 95188 433608
rect 95252 433606 95298 433666
rect 98361 433664 98500 433666
rect 98361 433608 98366 433664
rect 98422 433608 98500 433664
rect 98361 433606 98500 433608
rect 95252 433604 95258 433606
rect 95141 433603 95207 433604
rect 98361 433603 98427 433606
rect 98494 433604 98500 433606
rect 98564 433604 98570 433668
rect 99833 433666 99899 433669
rect 105169 433668 105235 433669
rect 99966 433666 99972 433668
rect 99833 433664 99972 433666
rect 99833 433608 99838 433664
rect 99894 433608 99972 433664
rect 99833 433606 99972 433608
rect 99833 433603 99899 433606
rect 99966 433604 99972 433606
rect 100036 433604 100042 433668
rect 105118 433666 105124 433668
rect 105078 433606 105124 433666
rect 105188 433664 105235 433668
rect 105230 433608 105235 433664
rect 105118 433604 105124 433606
rect 105188 433604 105235 433608
rect 106774 433604 106780 433668
rect 106844 433666 106850 433668
rect 110413 433666 110479 433669
rect 106844 433664 110479 433666
rect 106844 433608 110418 433664
rect 110474 433608 110479 433664
rect 106844 433606 110479 433608
rect 106844 433604 106850 433606
rect 105169 433603 105235 433604
rect 110413 433603 110479 433606
rect 111190 433604 111196 433668
rect 111260 433666 111266 433668
rect 111701 433666 111767 433669
rect 111260 433664 111767 433666
rect 111260 433608 111706 433664
rect 111762 433608 111767 433664
rect 111260 433606 111767 433608
rect 111260 433604 111266 433606
rect 111701 433603 111767 433606
rect 66345 433394 66411 433397
rect 66345 433392 68908 433394
rect 66345 433336 66350 433392
rect 66406 433336 68908 433392
rect 112118 433364 112178 433742
rect 66345 433334 68908 433336
rect 66345 433331 66411 433334
rect 67449 433260 67515 433261
rect 67398 433258 67404 433260
rect 67358 433198 67404 433258
rect 67468 433256 67515 433260
rect 67510 433200 67515 433256
rect 67398 433196 67404 433198
rect 67468 433196 67515 433200
rect 67449 433195 67515 433196
rect 112110 432788 112116 432852
rect 112180 432788 112186 432852
rect 66805 432578 66871 432581
rect 66805 432576 68908 432578
rect 66805 432520 66810 432576
rect 66866 432520 68908 432576
rect 66805 432518 68908 432520
rect 66805 432515 66871 432518
rect 112118 432306 112178 432788
rect 114737 432306 114803 432309
rect 112118 432304 114803 432306
rect 112118 432276 114742 432304
rect 112148 432248 114742 432276
rect 114798 432248 114803 432304
rect 112148 432246 114803 432248
rect 114737 432243 114803 432246
rect 583109 431626 583175 431629
rect 583520 431626 584960 431716
rect 583109 431624 584960 431626
rect 583109 431568 583114 431624
rect 583170 431568 584960 431624
rect 583109 431566 584960 431568
rect 583109 431563 583175 431566
rect 66805 431490 66871 431493
rect 66805 431488 68908 431490
rect 66805 431432 66810 431488
rect 66866 431432 68908 431488
rect 583520 431476 584960 431566
rect 66805 431430 68908 431432
rect 66805 431427 66871 431430
rect 113265 431218 113331 431221
rect 114737 431218 114803 431221
rect 112700 431216 114803 431218
rect 112700 431160 113270 431216
rect 113326 431160 114742 431216
rect 114798 431160 114803 431216
rect 112700 431158 114803 431160
rect 113265 431155 113331 431158
rect 114737 431155 114803 431158
rect 66805 430402 66871 430405
rect 66805 430400 68908 430402
rect 66805 430344 66810 430400
rect 66866 430344 68908 430400
rect 66805 430342 68908 430344
rect 66805 430339 66871 430342
rect 113449 430130 113515 430133
rect 112700 430128 113515 430130
rect 112700 430072 113454 430128
rect 113510 430072 113515 430128
rect 112700 430070 113515 430072
rect 113449 430067 113515 430070
rect 66253 429314 66319 429317
rect 113173 429314 113239 429317
rect 113817 429314 113883 429317
rect 66253 429312 68908 429314
rect 66253 429256 66258 429312
rect 66314 429256 68908 429312
rect 66253 429254 68908 429256
rect 112700 429312 113883 429314
rect 112700 429256 113178 429312
rect 113234 429256 113822 429312
rect 113878 429256 113883 429312
rect 112700 429254 113883 429256
rect 66253 429251 66319 429254
rect 113173 429251 113239 429254
rect 113817 429251 113883 429254
rect 66161 428226 66227 428229
rect 115381 428226 115447 428229
rect 66161 428224 68908 428226
rect 66161 428168 66166 428224
rect 66222 428168 68908 428224
rect 66161 428166 68908 428168
rect 112700 428224 115447 428226
rect 112700 428168 115386 428224
rect 115442 428168 115447 428224
rect 112700 428166 115447 428168
rect 66161 428163 66227 428166
rect 115381 428163 115447 428166
rect 66805 427410 66871 427413
rect 66805 427408 68908 427410
rect 66805 427352 66810 427408
rect 66866 427352 68908 427408
rect 66805 427350 68908 427352
rect 66805 427347 66871 427350
rect 112118 426596 112178 427108
rect 112110 426532 112116 426596
rect 112180 426532 112186 426596
rect 68878 425642 68938 426292
rect 115841 426050 115907 426053
rect 112700 426048 115907 426050
rect 112700 425992 115846 426048
rect 115902 425992 115907 426048
rect 112700 425990 115907 425992
rect 115841 425987 115907 425990
rect 64830 425582 68938 425642
rect 61878 425172 61884 425236
rect 61948 425234 61954 425236
rect 64830 425234 64890 425582
rect 61948 425174 64890 425234
rect 66529 425234 66595 425237
rect 66529 425232 68908 425234
rect 66529 425176 66534 425232
rect 66590 425176 68908 425232
rect 66529 425174 68908 425176
rect 61948 425172 61954 425174
rect 66529 425171 66595 425174
rect 114093 424962 114159 424965
rect 112700 424960 114159 424962
rect 112700 424904 114098 424960
rect 114154 424904 114159 424960
rect 112700 424902 114159 424904
rect 114093 424899 114159 424902
rect 66621 424146 66687 424149
rect 114645 424146 114711 424149
rect 115841 424146 115907 424149
rect 66621 424144 68908 424146
rect 66621 424088 66626 424144
rect 66682 424088 68908 424144
rect 66621 424086 68908 424088
rect 112700 424144 115907 424146
rect 112700 424088 114650 424144
rect 114706 424088 115846 424144
rect 115902 424088 115907 424144
rect 112700 424086 115907 424088
rect 66621 424083 66687 424086
rect 114645 424083 114711 424086
rect 115841 424083 115907 424086
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 66805 423330 66871 423333
rect 66805 423328 68908 423330
rect 66805 423272 66810 423328
rect 66866 423272 68908 423328
rect 66805 423270 68908 423272
rect 66805 423267 66871 423270
rect 115841 423058 115907 423061
rect 112700 423056 115907 423058
rect 112700 423000 115846 423056
rect 115902 423000 115907 423056
rect 112700 422998 115907 423000
rect 115841 422995 115907 422998
rect 66846 422180 66852 422244
rect 66916 422242 66922 422244
rect 66916 422182 68908 422242
rect 66916 422180 66922 422182
rect 115841 421970 115907 421973
rect 112700 421968 115907 421970
rect 112700 421912 115846 421968
rect 115902 421912 115907 421968
rect 112700 421910 115907 421912
rect 115841 421907 115907 421910
rect 66805 421154 66871 421157
rect 66805 421152 68908 421154
rect 66805 421096 66810 421152
rect 66866 421096 68908 421152
rect 66805 421094 68908 421096
rect 66805 421091 66871 421094
rect 112302 420340 112362 420852
rect 112294 420276 112300 420340
rect 112364 420276 112370 420340
rect 53741 420202 53807 420205
rect 66846 420202 66852 420204
rect 53741 420200 66852 420202
rect 53741 420144 53746 420200
rect 53802 420144 66852 420200
rect 53741 420142 66852 420144
rect 53741 420139 53807 420142
rect 66846 420140 66852 420142
rect 66916 420140 66922 420204
rect 66805 420066 66871 420069
rect 113173 420066 113239 420069
rect 66805 420064 68908 420066
rect 66805 420008 66810 420064
rect 66866 420008 68908 420064
rect 66805 420006 68908 420008
rect 112700 420064 113239 420066
rect 112700 420008 113178 420064
rect 113234 420008 113239 420064
rect 112700 420006 113239 420008
rect 66805 420003 66871 420006
rect 113173 420003 113239 420006
rect 114737 418978 114803 418981
rect 112700 418976 114803 418978
rect 68878 418434 68938 418948
rect 112700 418920 114742 418976
rect 114798 418920 114803 418976
rect 112700 418918 114803 418920
rect 114737 418915 114803 418918
rect 64830 418374 68938 418434
rect 61929 418298 61995 418301
rect 64830 418298 64890 418374
rect 61929 418296 64890 418298
rect 61929 418240 61934 418296
rect 61990 418240 64890 418296
rect 61929 418238 64890 418240
rect 583201 418298 583267 418301
rect 583520 418298 584960 418388
rect 583201 418296 584960 418298
rect 583201 418240 583206 418296
rect 583262 418240 584960 418296
rect 583201 418238 584960 418240
rect 61929 418235 61995 418238
rect 583201 418235 583267 418238
rect 66989 418162 67055 418165
rect 66989 418160 68908 418162
rect 66989 418104 66994 418160
rect 67050 418104 68908 418160
rect 583520 418148 584960 418238
rect 66989 418102 68908 418104
rect 66989 418099 67055 418102
rect 114645 417890 114711 417893
rect 112700 417888 114711 417890
rect 112700 417832 114650 417888
rect 114706 417832 114711 417888
rect 112700 417830 114711 417832
rect 114645 417827 114711 417830
rect 66805 417074 66871 417077
rect 66805 417072 68908 417074
rect 66805 417016 66810 417072
rect 66866 417016 68908 417072
rect 66805 417014 68908 417016
rect 66805 417011 66871 417014
rect 113357 416802 113423 416805
rect 115841 416802 115907 416805
rect 112700 416800 115907 416802
rect 112700 416744 113362 416800
rect 113418 416744 115846 416800
rect 115902 416744 115907 416800
rect 112700 416742 115907 416744
rect 113357 416739 113423 416742
rect 115841 416739 115907 416742
rect 66713 415986 66779 415989
rect 66713 415984 68908 415986
rect 66713 415928 66718 415984
rect 66774 415928 68908 415984
rect 66713 415926 68908 415928
rect 66713 415923 66779 415926
rect 115197 415714 115263 415717
rect 112700 415712 115263 415714
rect 112700 415656 115202 415712
rect 115258 415656 115263 415712
rect 112700 415654 115263 415656
rect 115197 415651 115263 415654
rect 66713 414898 66779 414901
rect 115841 414898 115907 414901
rect 66713 414896 68908 414898
rect 66713 414840 66718 414896
rect 66774 414840 68908 414896
rect 66713 414838 68908 414840
rect 112700 414896 115907 414898
rect 112700 414840 115846 414896
rect 115902 414840 115907 414896
rect 112700 414838 115907 414840
rect 66713 414835 66779 414838
rect 115841 414835 115907 414838
rect 67725 414082 67791 414085
rect 67725 414080 68908 414082
rect 67725 414024 67730 414080
rect 67786 414024 68908 414080
rect 67725 414022 68908 414024
rect 67725 414019 67791 414022
rect 115841 413810 115907 413813
rect 112700 413808 115907 413810
rect 112700 413752 115846 413808
rect 115902 413752 115907 413808
rect 112700 413750 115907 413752
rect 115841 413747 115907 413750
rect 66253 412994 66319 412997
rect 66253 412992 68908 412994
rect 66253 412936 66258 412992
rect 66314 412936 68908 412992
rect 66253 412934 68908 412936
rect 66253 412931 66319 412934
rect 115197 412722 115263 412725
rect 112700 412720 115263 412722
rect 112700 412664 115202 412720
rect 115258 412664 115263 412720
rect 112700 412662 115263 412664
rect 115197 412659 115263 412662
rect 59118 411300 59124 411364
rect 59188 411362 59194 411364
rect 64781 411362 64847 411365
rect 68878 411362 68938 411876
rect 115841 411634 115907 411637
rect 112700 411632 115907 411634
rect 112700 411576 115846 411632
rect 115902 411576 115907 411632
rect 112700 411574 115907 411576
rect 115841 411571 115907 411574
rect 59188 411360 68938 411362
rect 59188 411304 64786 411360
rect 64842 411304 68938 411360
rect 59188 411302 68938 411304
rect 59188 411300 59194 411302
rect 64781 411299 64847 411302
rect 66805 410818 66871 410821
rect 66805 410816 68908 410818
rect 66805 410760 66810 410816
rect 66866 410760 68908 410816
rect 66805 410758 68908 410760
rect 66805 410755 66871 410758
rect -960 410546 480 410636
rect 2865 410546 2931 410549
rect 115841 410546 115907 410549
rect -960 410544 2931 410546
rect -960 410488 2870 410544
rect 2926 410488 2931 410544
rect -960 410486 2931 410488
rect 112700 410544 115907 410546
rect 112700 410488 115846 410544
rect 115902 410488 115907 410544
rect 112700 410486 115907 410488
rect -960 410396 480 410486
rect 2865 410483 2931 410486
rect 115841 410483 115907 410486
rect 67449 409732 67515 409733
rect 67398 409730 67404 409732
rect 67322 409670 67404 409730
rect 67468 409730 67515 409732
rect 114502 409730 114508 409732
rect 67468 409728 68908 409730
rect 67510 409672 68908 409728
rect 67398 409668 67404 409670
rect 67468 409670 68908 409672
rect 112700 409670 114508 409730
rect 67468 409668 67515 409670
rect 114502 409668 114508 409670
rect 114572 409730 114578 409732
rect 115841 409730 115907 409733
rect 114572 409728 115907 409730
rect 114572 409672 115846 409728
rect 115902 409672 115907 409728
rect 114572 409670 115907 409672
rect 114572 409668 114578 409670
rect 67449 409667 67515 409668
rect 115841 409667 115907 409670
rect 66110 408852 66116 408916
rect 66180 408914 66186 408916
rect 66621 408914 66687 408917
rect 66180 408912 68908 408914
rect 66180 408856 66626 408912
rect 66682 408856 68908 408912
rect 66180 408854 68908 408856
rect 66180 408852 66186 408854
rect 66621 408851 66687 408854
rect 115054 408642 115060 408644
rect 112700 408582 115060 408642
rect 115054 408580 115060 408582
rect 115124 408580 115130 408644
rect 66805 407826 66871 407829
rect 66805 407824 68908 407826
rect 66805 407768 66810 407824
rect 66866 407768 68908 407824
rect 66805 407766 68908 407768
rect 66805 407763 66871 407766
rect 115841 407554 115907 407557
rect 112700 407552 115907 407554
rect 112700 407496 115846 407552
rect 115902 407496 115907 407552
rect 112700 407494 115907 407496
rect 115841 407491 115907 407494
rect 41229 407012 41295 407013
rect 41229 407008 41276 407012
rect 41340 407010 41346 407012
rect 56593 407010 56659 407013
rect 57830 407010 57836 407012
rect 41229 406952 41234 407008
rect 41229 406948 41276 406952
rect 41340 406950 41386 407010
rect 56593 407008 57836 407010
rect 56593 406952 56598 407008
rect 56654 406952 57836 407008
rect 56593 406950 57836 406952
rect 41340 406948 41346 406950
rect 41229 406947 41295 406948
rect 56593 406947 56659 406950
rect 57830 406948 57836 406950
rect 57900 406948 57906 407012
rect 68878 406058 68938 406708
rect 114553 406466 114619 406469
rect 114921 406466 114987 406469
rect 112700 406464 114987 406466
rect 112700 406408 114558 406464
rect 114614 406408 114926 406464
rect 114982 406408 114987 406464
rect 112700 406406 114987 406408
rect 114553 406403 114619 406406
rect 114921 406403 114987 406406
rect 64830 405998 68938 406058
rect 57830 405724 57836 405788
rect 57900 405786 57906 405788
rect 64830 405786 64890 405998
rect 57900 405726 64890 405786
rect 57900 405724 57906 405726
rect 66437 405650 66503 405653
rect 67541 405650 67607 405653
rect 115841 405650 115907 405653
rect 66437 405648 68908 405650
rect 66437 405592 66442 405648
rect 66498 405592 67546 405648
rect 67602 405592 68908 405648
rect 66437 405590 68908 405592
rect 112700 405648 115907 405650
rect 112700 405592 115846 405648
rect 115902 405592 115907 405648
rect 112700 405590 115907 405592
rect 66437 405587 66503 405590
rect 67541 405587 67607 405590
rect 115841 405587 115907 405590
rect 583293 404970 583359 404973
rect 583520 404970 584960 405060
rect 583293 404968 584960 404970
rect 583293 404912 583298 404968
rect 583354 404912 584960 404968
rect 583293 404910 584960 404912
rect 583293 404907 583359 404910
rect 583520 404820 584960 404910
rect 66805 404562 66871 404565
rect 115565 404562 115631 404565
rect 66805 404560 68908 404562
rect 66805 404504 66810 404560
rect 66866 404504 68908 404560
rect 66805 404502 68908 404504
rect 112700 404560 115631 404562
rect 112700 404504 115570 404560
rect 115626 404504 115631 404560
rect 112700 404502 115631 404504
rect 66805 404499 66871 404502
rect 115565 404499 115631 404502
rect 66805 403746 66871 403749
rect 66805 403744 68908 403746
rect 66805 403688 66810 403744
rect 66866 403688 68908 403744
rect 66805 403686 68908 403688
rect 66805 403683 66871 403686
rect 115841 403474 115907 403477
rect 112700 403472 115907 403474
rect 112700 403416 115846 403472
rect 115902 403416 115907 403472
rect 112700 403414 115907 403416
rect 115841 403411 115907 403414
rect 66345 402658 66411 402661
rect 66345 402656 68908 402658
rect 66345 402600 66350 402656
rect 66406 402600 68908 402656
rect 66345 402598 68908 402600
rect 66345 402595 66411 402598
rect 116117 402386 116183 402389
rect 112700 402384 116183 402386
rect 112700 402328 116122 402384
rect 116178 402328 116183 402384
rect 112700 402326 116183 402328
rect 116117 402323 116183 402326
rect 65885 401570 65951 401573
rect 65885 401568 68908 401570
rect 65885 401512 65890 401568
rect 65946 401512 68908 401568
rect 65885 401510 68908 401512
rect 65885 401507 65951 401510
rect 115657 401298 115723 401301
rect 112700 401296 115723 401298
rect 112700 401240 115662 401296
rect 115718 401240 115723 401296
rect 112700 401238 115723 401240
rect 115657 401235 115723 401238
rect 66805 400482 66871 400485
rect 115013 400482 115079 400485
rect 66805 400480 68908 400482
rect 66805 400424 66810 400480
rect 66866 400424 68908 400480
rect 66805 400422 68908 400424
rect 112700 400480 115079 400482
rect 112700 400424 115018 400480
rect 115074 400424 115079 400480
rect 112700 400422 115079 400424
rect 66805 400419 66871 400422
rect 115013 400419 115079 400422
rect 66805 399666 66871 399669
rect 66805 399664 68908 399666
rect 66805 399608 66810 399664
rect 66866 399608 68908 399664
rect 66805 399606 68908 399608
rect 66805 399603 66871 399606
rect 115197 399394 115263 399397
rect 112700 399392 115263 399394
rect 112700 399336 115202 399392
rect 115258 399336 115263 399392
rect 112700 399334 115263 399336
rect 115197 399331 115263 399334
rect 66805 398578 66871 398581
rect 66805 398576 68908 398578
rect 66805 398520 66810 398576
rect 66866 398520 68908 398576
rect 66805 398518 68908 398520
rect 66805 398515 66871 398518
rect 115841 398306 115907 398309
rect 112700 398304 115907 398306
rect 112700 398248 115846 398304
rect 115902 398248 115907 398304
rect 112700 398246 115907 398248
rect 115841 398243 115907 398246
rect 69422 397700 69428 397764
rect 69492 397700 69498 397764
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 17217 397490 17283 397493
rect 66897 397490 66963 397493
rect 69430 397490 69490 397700
rect 17217 397488 69490 397490
rect 17217 397432 17222 397488
rect 17278 397432 66902 397488
rect 66958 397460 69490 397488
rect 66958 397432 69460 397460
rect 17217 397430 69460 397432
rect 17217 397427 17283 397430
rect 66897 397427 66963 397430
rect 115841 397218 115907 397221
rect 112700 397216 115907 397218
rect 112700 397160 115846 397216
rect 115902 397160 115907 397216
rect 112700 397158 115907 397160
rect 115841 397155 115907 397158
rect 123334 396612 123340 396676
rect 123404 396674 123410 396676
rect 124121 396674 124187 396677
rect 132585 396674 132651 396677
rect 123404 396672 132651 396674
rect 123404 396616 124126 396672
rect 124182 396616 132590 396672
rect 132646 396616 132651 396672
rect 123404 396614 132651 396616
rect 123404 396612 123410 396614
rect 124121 396611 124187 396614
rect 132585 396611 132651 396614
rect 66805 396402 66871 396405
rect 113214 396402 113220 396404
rect 66805 396400 68908 396402
rect 66805 396344 66810 396400
rect 66866 396344 68908 396400
rect 66805 396342 68908 396344
rect 112700 396342 113220 396402
rect 66805 396339 66871 396342
rect 113214 396340 113220 396342
rect 113284 396402 113290 396404
rect 115841 396402 115907 396405
rect 113284 396400 115907 396402
rect 113284 396344 115846 396400
rect 115902 396344 115907 396400
rect 113284 396342 115907 396344
rect 113284 396340 113290 396342
rect 115841 396339 115907 396342
rect 66805 395314 66871 395317
rect 115841 395314 115907 395317
rect 66805 395312 68908 395314
rect 66805 395256 66810 395312
rect 66866 395256 68908 395312
rect 66805 395254 68908 395256
rect 112700 395312 115907 395314
rect 112700 395256 115846 395312
rect 115902 395256 115907 395312
rect 112700 395254 115907 395256
rect 66805 395251 66871 395254
rect 115841 395251 115907 395254
rect 66805 394498 66871 394501
rect 66805 394496 68908 394498
rect 66805 394440 66810 394496
rect 66866 394440 68908 394496
rect 66805 394438 68908 394440
rect 66805 394435 66871 394438
rect 115565 394226 115631 394229
rect 112700 394224 115631 394226
rect 112700 394168 115570 394224
rect 115626 394168 115631 394224
rect 112700 394166 115631 394168
rect 115565 394163 115631 394166
rect 49601 393546 49667 393549
rect 58985 393546 59051 393549
rect 49601 393544 64890 393546
rect 49601 393488 49606 393544
rect 49662 393488 58990 393544
rect 59046 393488 64890 393544
rect 49601 393486 64890 393488
rect 49601 393483 49667 393486
rect 58985 393483 59051 393486
rect 64830 393410 64890 393486
rect 64830 393350 68908 393410
rect 115841 393138 115907 393141
rect 112700 393136 115907 393138
rect 112700 393080 115846 393136
rect 115902 393080 115907 393136
rect 112700 393078 115907 393080
rect 115841 393075 115907 393078
rect 66805 392322 66871 392325
rect 66805 392320 68908 392322
rect 66805 392264 66810 392320
rect 66866 392264 68908 392320
rect 66805 392262 68908 392264
rect 66805 392259 66871 392262
rect 4061 392186 4127 392189
rect 69606 392186 69612 392188
rect 4061 392184 69612 392186
rect 4061 392128 4066 392184
rect 4122 392128 69612 392184
rect 4061 392126 69612 392128
rect 4061 392123 4127 392126
rect 69606 392124 69612 392126
rect 69676 392124 69682 392188
rect 115841 392050 115907 392053
rect 112700 392048 115907 392050
rect 112700 391992 115846 392048
rect 115902 391992 115907 392048
rect 112700 391990 115907 391992
rect 115841 391987 115907 391990
rect 7557 391914 7623 391917
rect 107694 391914 107700 391916
rect 7557 391912 107700 391914
rect 7557 391856 7562 391912
rect 7618 391856 107700 391912
rect 7557 391854 107700 391856
rect 7557 391851 7623 391854
rect 107694 391852 107700 391854
rect 107764 391852 107770 391916
rect 583520 391628 584960 391868
rect 66805 391234 66871 391237
rect 66805 391232 68908 391234
rect 66805 391176 66810 391232
rect 66866 391176 68908 391232
rect 66805 391174 68908 391176
rect 66805 391171 66871 391174
rect 82077 391100 82143 391101
rect 85481 391100 85547 391101
rect 82077 391098 82124 391100
rect 82032 391096 82124 391098
rect 82032 391040 82082 391096
rect 82032 391038 82124 391040
rect 82077 391036 82124 391038
rect 82188 391036 82194 391100
rect 85430 391098 85436 391100
rect 85390 391038 85436 391098
rect 85500 391096 85547 391100
rect 85542 391040 85547 391096
rect 85430 391036 85436 391038
rect 85500 391036 85547 391040
rect 88742 391036 88748 391100
rect 88812 391098 88818 391100
rect 89667 391098 89733 391101
rect 88812 391096 89733 391098
rect 88812 391040 89672 391096
rect 89728 391040 89733 391096
rect 88812 391038 89733 391040
rect 88812 391036 88818 391038
rect 82077 391035 82143 391036
rect 85481 391035 85547 391036
rect 89667 391035 89733 391038
rect 92606 391036 92612 391100
rect 92676 391098 92682 391100
rect 92749 391098 92815 391101
rect 92676 391096 92815 391098
rect 92676 391040 92754 391096
rect 92810 391040 92815 391096
rect 92676 391038 92815 391040
rect 92676 391036 92682 391038
rect 92749 391035 92815 391038
rect 100661 390964 100727 390965
rect 100661 390962 100708 390964
rect 100616 390960 100708 390962
rect 100616 390904 100666 390960
rect 100616 390902 100708 390904
rect 100661 390900 100708 390902
rect 100772 390900 100778 390964
rect 100661 390899 100727 390900
rect 77477 390690 77543 390693
rect 107745 390692 107811 390693
rect 78438 390690 78444 390692
rect 77477 390688 78444 390690
rect 77477 390632 77482 390688
rect 77538 390632 78444 390688
rect 77477 390630 78444 390632
rect 77477 390627 77543 390630
rect 78438 390628 78444 390630
rect 78508 390628 78514 390692
rect 107694 390690 107700 390692
rect 107654 390630 107700 390690
rect 107764 390688 107811 390692
rect 107806 390632 107811 390688
rect 107694 390628 107700 390630
rect 107764 390628 107811 390632
rect 108246 390628 108252 390692
rect 108316 390690 108322 390692
rect 108757 390690 108823 390693
rect 108316 390688 108823 390690
rect 108316 390632 108762 390688
rect 108818 390632 108823 390688
rect 108316 390630 108823 390632
rect 108316 390628 108322 390630
rect 107745 390627 107811 390628
rect 108757 390627 108823 390630
rect 111701 390690 111767 390693
rect 112118 390690 112178 391204
rect 111701 390688 112178 390690
rect 111701 390632 111706 390688
rect 111762 390632 112178 390688
rect 111701 390630 112178 390632
rect 111701 390627 111767 390630
rect 72417 390418 72483 390421
rect 77201 390420 77267 390421
rect 72550 390418 72556 390420
rect 72417 390416 72556 390418
rect 72417 390360 72422 390416
rect 72478 390360 72556 390416
rect 72417 390358 72556 390360
rect 72417 390355 72483 390358
rect 72550 390356 72556 390358
rect 72620 390356 72626 390420
rect 77150 390418 77156 390420
rect 77110 390358 77156 390418
rect 77220 390416 77267 390420
rect 77262 390360 77267 390416
rect 77150 390356 77156 390358
rect 77220 390356 77267 390360
rect 104934 390356 104940 390420
rect 105004 390418 105010 390420
rect 105261 390418 105327 390421
rect 105004 390416 105327 390418
rect 105004 390360 105266 390416
rect 105322 390360 105327 390416
rect 105004 390358 105327 390360
rect 105004 390356 105010 390358
rect 77201 390355 77267 390356
rect 105261 390355 105327 390358
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106733 390418 106799 390421
rect 106476 390416 106799 390418
rect 106476 390360 106738 390416
rect 106794 390360 106799 390416
rect 106476 390358 106799 390360
rect 106476 390356 106482 390358
rect 106733 390355 106799 390358
rect 62021 389330 62087 389333
rect 98453 389330 98519 389333
rect 128670 389330 128676 389332
rect 62021 389328 128676 389330
rect 62021 389272 62026 389328
rect 62082 389272 98458 389328
rect 98514 389272 128676 389328
rect 62021 389270 128676 389272
rect 62021 389267 62087 389270
rect 98453 389267 98519 389270
rect 128670 389268 128676 389270
rect 128740 389268 128746 389332
rect 50889 389194 50955 389197
rect 103513 389194 103579 389197
rect 103789 389194 103855 389197
rect 50889 389192 103855 389194
rect 50889 389136 50894 389192
rect 50950 389136 103518 389192
rect 103574 389136 103794 389192
rect 103850 389136 103855 389192
rect 50889 389134 103855 389136
rect 50889 389131 50955 389134
rect 103513 389131 103579 389134
rect 103789 389131 103855 389134
rect 71865 389060 71931 389061
rect 71814 388996 71820 389060
rect 71884 389058 71931 389060
rect 76005 389058 76071 389061
rect 76741 389058 76807 389061
rect 71884 389056 71976 389058
rect 71926 389000 71976 389056
rect 71884 388998 71976 389000
rect 76005 389056 76807 389058
rect 76005 389000 76010 389056
rect 76066 389000 76746 389056
rect 76802 389000 76807 389056
rect 76005 388998 76807 389000
rect 71884 388996 71931 388998
rect 71865 388995 71931 388996
rect 76005 388995 76071 388998
rect 76741 388995 76807 388998
rect 78949 389058 79015 389061
rect 79910 389058 79916 389060
rect 78949 389056 79916 389058
rect 78949 389000 78954 389056
rect 79010 389000 79916 389056
rect 78949 388998 79916 389000
rect 78949 388995 79015 388998
rect 79910 388996 79916 388998
rect 79980 389058 79986 389060
rect 86217 389058 86283 389061
rect 79980 389056 86283 389058
rect 79980 389000 86222 389056
rect 86278 389000 86283 389056
rect 79980 388998 86283 389000
rect 79980 388996 79986 388998
rect 86217 388995 86283 388998
rect 89161 389058 89227 389061
rect 91502 389058 91508 389060
rect 89161 389056 91508 389058
rect 89161 389000 89166 389056
rect 89222 389000 91508 389056
rect 89161 388998 91508 389000
rect 89161 388995 89227 388998
rect 91502 388996 91508 388998
rect 91572 389058 91578 389060
rect 93209 389058 93275 389061
rect 91572 389056 93275 389058
rect 91572 389000 93214 389056
rect 93270 389000 93275 389056
rect 91572 388998 93275 389000
rect 91572 388996 91578 388998
rect 93209 388995 93275 388998
rect 94446 388996 94452 389060
rect 94516 389058 94522 389060
rect 99741 389058 99807 389061
rect 100109 389058 100175 389061
rect 94516 389056 100175 389058
rect 94516 389000 99746 389056
rect 99802 389000 100114 389056
rect 100170 389000 100175 389056
rect 94516 388998 100175 389000
rect 94516 388996 94522 388998
rect 99741 388995 99807 388998
rect 100109 388995 100175 388998
rect 107745 389058 107811 389061
rect 108941 389058 109007 389061
rect 107745 389056 109007 389058
rect 107745 389000 107750 389056
rect 107806 389000 108946 389056
rect 109002 389000 109007 389056
rect 107745 388998 109007 389000
rect 107745 388995 107811 388998
rect 108941 388995 109007 388998
rect 121453 389058 121519 389061
rect 124254 389058 124260 389060
rect 121453 389056 124260 389058
rect 121453 389000 121458 389056
rect 121514 389000 124260 389056
rect 121453 388998 124260 389000
rect 121453 388995 121519 388998
rect 124254 388996 124260 388998
rect 124324 388996 124330 389060
rect 69606 388860 69612 388924
rect 69676 388922 69682 388924
rect 93853 388922 93919 388925
rect 94589 388922 94655 388925
rect 69676 388920 94655 388922
rect 69676 388864 93858 388920
rect 93914 388864 94594 388920
rect 94650 388864 94655 388920
rect 69676 388862 94655 388864
rect 69676 388860 69682 388862
rect 93853 388859 93919 388862
rect 94589 388859 94655 388862
rect 29637 388786 29703 388789
rect 81525 388786 81591 388789
rect 29637 388784 81591 388786
rect 29637 388728 29642 388784
rect 29698 388728 81530 388784
rect 81586 388728 81591 388784
rect 29637 388726 81591 388728
rect 29637 388723 29703 388726
rect 81525 388723 81591 388726
rect 100518 388452 100524 388516
rect 100588 388514 100594 388516
rect 100661 388514 100727 388517
rect 100588 388512 100727 388514
rect 100588 388456 100666 388512
rect 100722 388456 100727 388512
rect 100588 388454 100727 388456
rect 100588 388452 100594 388454
rect 100661 388451 100727 388454
rect 102317 388514 102383 388517
rect 103278 388514 103284 388516
rect 102317 388512 103284 388514
rect 102317 388456 102322 388512
rect 102378 388456 103284 388512
rect 102317 388454 103284 388456
rect 102317 388451 102383 388454
rect 103278 388452 103284 388454
rect 103348 388452 103354 388516
rect 99465 388378 99531 388381
rect 106406 388378 106412 388380
rect 99465 388376 106412 388378
rect 99465 388320 99470 388376
rect 99526 388320 106412 388376
rect 99465 388318 106412 388320
rect 99465 388315 99531 388318
rect 106406 388316 106412 388318
rect 106476 388316 106482 388380
rect 55121 387970 55187 387973
rect 55078 387968 55187 387970
rect 55078 387912 55126 387968
rect 55182 387912 55187 387968
rect 55078 387907 55187 387912
rect 80053 387970 80119 387973
rect 80646 387970 80652 387972
rect 80053 387968 80652 387970
rect 80053 387912 80058 387968
rect 80114 387912 80652 387968
rect 80053 387910 80652 387912
rect 80053 387907 80119 387910
rect 80646 387908 80652 387910
rect 80716 387908 80722 387972
rect 50889 387698 50955 387701
rect 55078 387698 55138 387907
rect 110689 387834 110755 387837
rect 111006 387834 111012 387836
rect 110689 387832 111012 387834
rect 110689 387776 110694 387832
rect 110750 387776 111012 387832
rect 110689 387774 111012 387776
rect 110689 387771 110755 387774
rect 111006 387772 111012 387774
rect 111076 387772 111082 387836
rect 80973 387698 81039 387701
rect 50889 387696 81039 387698
rect 50889 387640 50894 387696
rect 50950 387640 80978 387696
rect 81034 387640 81039 387696
rect 50889 387638 81039 387640
rect 50889 387635 50955 387638
rect 80973 387635 81039 387638
rect 82721 387698 82787 387701
rect 86166 387698 86172 387700
rect 82721 387696 86172 387698
rect 82721 387640 82726 387696
rect 82782 387640 86172 387696
rect 82721 387638 86172 387640
rect 82721 387635 82787 387638
rect 86166 387636 86172 387638
rect 86236 387636 86242 387700
rect 61694 387500 61700 387564
rect 61764 387562 61770 387564
rect 66805 387562 66871 387565
rect 61764 387560 66871 387562
rect 61764 387504 66810 387560
rect 66866 387504 66871 387560
rect 61764 387502 66871 387504
rect 61764 387500 61770 387502
rect 66805 387499 66871 387502
rect 89621 387154 89687 387157
rect 99966 387154 99972 387156
rect 89621 387152 99972 387154
rect 89621 387096 89626 387152
rect 89682 387096 99972 387152
rect 89621 387094 99972 387096
rect 89621 387091 89687 387094
rect 99966 387092 99972 387094
rect 100036 387092 100042 387156
rect 102041 387154 102107 387157
rect 111742 387154 111748 387156
rect 102041 387152 111748 387154
rect 102041 387096 102046 387152
rect 102102 387096 111748 387152
rect 102041 387094 111748 387096
rect 102041 387091 102107 387094
rect 111742 387092 111748 387094
rect 111812 387092 111818 387156
rect 93761 387018 93827 387021
rect 105118 387018 105124 387020
rect 93761 387016 105124 387018
rect 93761 386960 93766 387016
rect 93822 386960 105124 387016
rect 93761 386958 105124 386960
rect 93761 386955 93827 386958
rect 105118 386956 105124 386958
rect 105188 386956 105194 387020
rect 55121 386476 55187 386477
rect 55070 386474 55076 386476
rect 55030 386414 55076 386474
rect 55140 386472 55187 386476
rect 55182 386416 55187 386472
rect 55070 386412 55076 386414
rect 55140 386412 55187 386416
rect 55121 386411 55187 386412
rect 75821 386338 75887 386341
rect 78254 386338 78260 386340
rect 75821 386336 78260 386338
rect 75821 386280 75826 386336
rect 75882 386280 78260 386336
rect 75821 386278 78260 386280
rect 75821 386275 75887 386278
rect 78254 386276 78260 386278
rect 78324 386276 78330 386340
rect 89529 385658 89595 385661
rect 97390 385658 97396 385660
rect 89529 385656 97396 385658
rect 89529 385600 89534 385656
rect 89590 385600 97396 385656
rect 89529 385598 97396 385600
rect 89529 385595 89595 385598
rect 97390 385596 97396 385598
rect 97460 385596 97466 385660
rect 97809 385658 97875 385661
rect 106774 385658 106780 385660
rect 97809 385656 106780 385658
rect 97809 385600 97814 385656
rect 97870 385600 106780 385656
rect 97809 385598 106780 385600
rect 97809 385595 97875 385598
rect 106774 385596 106780 385598
rect 106844 385596 106850 385660
rect 70301 385114 70367 385117
rect 75862 385114 75868 385116
rect 70301 385112 75868 385114
rect 70301 385056 70306 385112
rect 70362 385056 75868 385112
rect 70301 385054 75868 385056
rect 70301 385051 70367 385054
rect 75862 385052 75868 385054
rect 75932 385052 75938 385116
rect 79961 385114 80027 385117
rect 84694 385114 84700 385116
rect 79961 385112 84700 385114
rect 79961 385056 79966 385112
rect 80022 385056 84700 385112
rect 79961 385054 84700 385056
rect 79961 385051 80027 385054
rect 84694 385052 84700 385054
rect 84764 385052 84770 385116
rect -960 384284 480 384524
rect 72969 384434 73035 384437
rect 80278 384434 80284 384436
rect 72969 384432 80284 384434
rect 72969 384376 72974 384432
rect 73030 384376 80284 384432
rect 72969 384374 80284 384376
rect 72969 384371 73035 384374
rect 80278 384372 80284 384374
rect 80348 384372 80354 384436
rect 43989 384298 44055 384301
rect 71814 384298 71820 384300
rect 43989 384296 71820 384298
rect 43989 384240 43994 384296
rect 44050 384240 71820 384296
rect 43989 384238 71820 384240
rect 43989 384235 44055 384238
rect 71814 384236 71820 384238
rect 71884 384236 71890 384300
rect 78581 383754 78647 383757
rect 85798 383754 85804 383756
rect 78581 383752 85804 383754
rect 78581 383696 78586 383752
rect 78642 383696 85804 383752
rect 78581 383694 85804 383696
rect 78581 383691 78647 383694
rect 85798 383692 85804 383694
rect 85868 383692 85874 383756
rect 126881 383754 126947 383757
rect 133822 383754 133828 383756
rect 126881 383752 133828 383754
rect 126881 383696 126886 383752
rect 126942 383696 133828 383752
rect 126881 383694 133828 383696
rect 126881 383691 126947 383694
rect 133822 383692 133828 383694
rect 133892 383692 133898 383756
rect 104893 383618 104959 383621
rect 117497 383618 117563 383621
rect 104893 383616 117563 383618
rect 104893 383560 104898 383616
rect 104954 383560 117502 383616
rect 117558 383560 117563 383616
rect 104893 383558 117563 383560
rect 104893 383555 104959 383558
rect 117497 383555 117563 383558
rect 86861 382394 86927 382397
rect 91093 382394 91159 382397
rect 86861 382392 91159 382394
rect 86861 382336 86866 382392
rect 86922 382336 91098 382392
rect 91154 382336 91159 382392
rect 86861 382334 91159 382336
rect 86861 382331 86927 382334
rect 91093 382331 91159 382334
rect 104893 382394 104959 382397
rect 106038 382394 106044 382396
rect 104893 382392 106044 382394
rect 104893 382336 104898 382392
rect 104954 382336 106044 382392
rect 104893 382334 106044 382336
rect 104893 382331 104959 382334
rect 106038 382332 106044 382334
rect 106108 382332 106114 382396
rect 97993 381578 98059 381581
rect 111190 381578 111196 381580
rect 97993 381576 111196 381578
rect 97993 381520 97998 381576
rect 98054 381520 111196 381576
rect 97993 381518 111196 381520
rect 97993 381515 98059 381518
rect 111190 381516 111196 381518
rect 111260 381516 111266 381580
rect 71681 380898 71747 380901
rect 74574 380898 74580 380900
rect 71681 380896 74580 380898
rect 71681 380840 71686 380896
rect 71742 380840 74580 380896
rect 71681 380838 74580 380840
rect 71681 380835 71747 380838
rect 74574 380836 74580 380838
rect 74644 380836 74650 380900
rect 85389 380218 85455 380221
rect 95182 380218 95188 380220
rect 85389 380216 95188 380218
rect 85389 380160 85394 380216
rect 85450 380160 95188 380216
rect 85389 380158 95188 380160
rect 85389 380155 85455 380158
rect 95182 380156 95188 380158
rect 95252 380156 95258 380220
rect 75177 379538 75243 379541
rect 81934 379538 81940 379540
rect 75177 379536 81940 379538
rect 75177 379480 75182 379536
rect 75238 379480 81940 379536
rect 75177 379478 81940 379480
rect 75177 379475 75243 379478
rect 81934 379476 81940 379478
rect 82004 379476 82010 379540
rect 85297 378722 85363 378725
rect 93894 378722 93900 378724
rect 85297 378720 93900 378722
rect 85297 378664 85302 378720
rect 85358 378664 93900 378720
rect 85297 378662 93900 378664
rect 85297 378659 85363 378662
rect 93894 378660 93900 378662
rect 93964 378660 93970 378724
rect 583385 378450 583451 378453
rect 583520 378450 584960 378540
rect 583385 378448 584960 378450
rect 583385 378392 583390 378448
rect 583446 378392 584960 378448
rect 583385 378390 584960 378392
rect 583385 378387 583451 378390
rect 583520 378300 584960 378390
rect 81249 377362 81315 377365
rect 89662 377362 89668 377364
rect 81249 377360 89668 377362
rect 81249 377304 81254 377360
rect 81310 377304 89668 377360
rect 81249 377302 89668 377304
rect 81249 377299 81315 377302
rect 89662 377300 89668 377302
rect 89732 377300 89738 377364
rect 88241 373282 88307 373285
rect 98126 373282 98132 373284
rect 88241 373280 98132 373282
rect 88241 373224 88246 373280
rect 88302 373224 98132 373280
rect 88241 373222 98132 373224
rect 88241 373219 88307 373222
rect 98126 373220 98132 373222
rect 98196 373220 98202 373284
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 86217 369066 86283 369069
rect 107694 369066 107700 369068
rect 86217 369064 107700 369066
rect 86217 369008 86222 369064
rect 86278 369008 107700 369064
rect 86217 369006 107700 369008
rect 86217 369003 86283 369006
rect 107694 369004 107700 369006
rect 107764 369004 107770 369068
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 93669 364986 93735 364989
rect 102174 364986 102180 364988
rect 93669 364984 102180 364986
rect 93669 364928 93674 364984
rect 93730 364928 102180 364984
rect 93669 364926 102180 364928
rect 93669 364923 93735 364926
rect 102174 364924 102180 364926
rect 102244 364924 102250 364988
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 583520 351930 584960 352020
rect 583342 351870 584960 351930
rect 583342 351794 583402 351870
rect 583520 351794 584960 351870
rect 583342 351780 584960 351794
rect 583342 351734 583586 351780
rect 583526 351661 583586 351734
rect 583477 351656 583586 351661
rect 583477 351600 583482 351656
rect 583538 351600 583586 351656
rect 583477 351598 583586 351600
rect 583477 351595 583543 351598
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 73470 343708 73476 343772
rect 73540 343770 73546 343772
rect 73797 343770 73863 343773
rect 73540 343768 73863 343770
rect 73540 343712 73802 343768
rect 73858 343712 73863 343768
rect 73540 343710 73863 343712
rect 73540 343708 73546 343710
rect 73797 343707 73863 343710
rect 75269 340914 75335 340917
rect 75678 340914 75684 340916
rect 75269 340912 75684 340914
rect 75269 340856 75274 340912
rect 75330 340856 75684 340912
rect 75269 340854 75684 340856
rect 75269 340851 75335 340854
rect 75678 340852 75684 340854
rect 75748 340852 75754 340916
rect 83549 339556 83615 339557
rect 82854 339492 82860 339556
rect 82924 339554 82930 339556
rect 83549 339554 83596 339556
rect 82924 339552 83596 339554
rect 83660 339554 83666 339556
rect 82924 339496 83554 339552
rect 82924 339494 83596 339496
rect 82924 339492 82930 339494
rect 83549 339492 83596 339494
rect 83660 339494 83742 339554
rect 83660 339492 83666 339494
rect 83549 339491 83615 339492
rect 43805 338738 43871 338741
rect 77293 338738 77359 338741
rect 248413 338738 248479 338741
rect 43805 338736 248479 338738
rect 43805 338680 43810 338736
rect 43866 338680 77298 338736
rect 77354 338680 248418 338736
rect 248474 338680 248479 338736
rect 43805 338678 248479 338680
rect 43805 338675 43871 338678
rect 77293 338675 77359 338678
rect 248413 338675 248479 338678
rect 583520 338452 584960 338692
rect 69657 338058 69723 338061
rect 70158 338058 70164 338060
rect 69657 338056 70164 338058
rect 69657 338000 69662 338056
rect 69718 338000 70164 338056
rect 69657 337998 70164 338000
rect 69657 337995 69723 337998
rect 70158 337996 70164 337998
rect 70228 337996 70234 338060
rect 102225 335474 102291 335477
rect 102726 335474 102732 335476
rect 102225 335472 102732 335474
rect 102225 335416 102230 335472
rect 102286 335416 102732 335472
rect 102225 335414 102732 335416
rect 102225 335411 102291 335414
rect 102726 335412 102732 335414
rect 102796 335474 102802 335476
rect 246297 335474 246363 335477
rect 102796 335472 246363 335474
rect 102796 335416 246302 335472
rect 246358 335416 246363 335472
rect 102796 335414 246363 335416
rect 102796 335412 102802 335414
rect 246297 335411 246363 335414
rect 65885 334114 65951 334117
rect 66110 334114 66116 334116
rect 65885 334112 66116 334114
rect 65885 334056 65890 334112
rect 65946 334056 66116 334112
rect 65885 334054 66116 334056
rect 65885 334051 65951 334054
rect 66110 334052 66116 334054
rect 66180 334114 66186 334116
rect 244917 334114 244983 334117
rect 66180 334112 244983 334114
rect 66180 334056 244922 334112
rect 244978 334056 244983 334112
rect 66180 334054 244983 334056
rect 66180 334052 66186 334054
rect 244917 334051 244983 334054
rect 82629 333298 82695 333301
rect 91318 333298 91324 333300
rect 82629 333296 91324 333298
rect 82629 333240 82634 333296
rect 82690 333240 91324 333296
rect 82629 333238 91324 333240
rect 82629 333235 82695 333238
rect 91318 333236 91324 333238
rect 91388 333236 91394 333300
rect 91502 332692 91508 332756
rect 91572 332754 91578 332756
rect 92381 332754 92447 332757
rect 91572 332752 92447 332754
rect 91572 332696 92386 332752
rect 92442 332696 92447 332752
rect 91572 332694 92447 332696
rect 91572 332692 91578 332694
rect 92381 332691 92447 332694
rect 92974 332692 92980 332756
rect 93044 332754 93050 332756
rect 93710 332754 93716 332756
rect 93044 332694 93716 332754
rect 93044 332692 93050 332694
rect 93710 332692 93716 332694
rect 93780 332754 93786 332756
rect 263685 332754 263751 332757
rect 93780 332752 263751 332754
rect 93780 332696 263690 332752
rect 263746 332696 263751 332752
rect 93780 332694 263751 332696
rect 93780 332692 93786 332694
rect 263685 332691 263751 332694
rect 79174 332556 79180 332620
rect 79244 332618 79250 332620
rect 258257 332618 258323 332621
rect 79244 332616 258323 332618
rect 79244 332560 258262 332616
rect 258318 332560 258323 332616
rect 79244 332558 258323 332560
rect 79244 332556 79250 332558
rect 258257 332555 258323 332558
rect -960 332196 480 332436
rect 57697 331258 57763 331261
rect 262397 331258 262463 331261
rect 57697 331256 262463 331258
rect 57697 331200 57702 331256
rect 57758 331200 262402 331256
rect 262458 331200 262463 331256
rect 57697 331198 262463 331200
rect 57697 331195 57763 331198
rect 262397 331195 262463 331198
rect 108246 330380 108252 330444
rect 108316 330442 108322 330444
rect 111701 330442 111767 330445
rect 255446 330442 255452 330444
rect 108316 330440 255452 330442
rect 108316 330384 111706 330440
rect 111762 330384 255452 330440
rect 108316 330382 255452 330384
rect 108316 330380 108322 330382
rect 111701 330379 111767 330382
rect 255446 330380 255452 330382
rect 255516 330380 255522 330444
rect 97942 329836 97948 329900
rect 98012 329898 98018 329900
rect 99281 329898 99347 329901
rect 98012 329896 99347 329898
rect 98012 329840 99286 329896
rect 99342 329840 99347 329896
rect 98012 329838 99347 329840
rect 98012 329836 98018 329838
rect 99281 329835 99347 329838
rect 84101 329082 84167 329085
rect 87086 329082 87092 329084
rect 84101 329080 87092 329082
rect 84101 329024 84106 329080
rect 84162 329024 87092 329080
rect 84101 329022 87092 329024
rect 84101 329019 84167 329022
rect 87086 329020 87092 329022
rect 87156 329020 87162 329084
rect 70485 328538 70551 328541
rect 71446 328538 71452 328540
rect 70485 328536 71452 328538
rect 70485 328480 70490 328536
rect 70546 328480 71452 328536
rect 70485 328478 71452 328480
rect 70485 328475 70551 328478
rect 71446 328476 71452 328478
rect 71516 328538 71522 328540
rect 256785 328538 256851 328541
rect 71516 328536 256851 328538
rect 71516 328480 256790 328536
rect 256846 328480 256851 328536
rect 71516 328478 256851 328480
rect 71516 328476 71522 328478
rect 256785 328475 256851 328478
rect 94998 326980 95004 327044
rect 95068 327042 95074 327044
rect 102133 327042 102199 327045
rect 95068 327040 102199 327042
rect 95068 326984 102138 327040
rect 102194 326984 102199 327040
rect 95068 326982 102199 326984
rect 95068 326980 95074 326982
rect 102133 326979 102199 326982
rect 67541 326362 67607 326365
rect 245009 326362 245075 326365
rect 67541 326360 245075 326362
rect 67541 326304 67546 326360
rect 67602 326304 245014 326360
rect 245070 326304 245075 326360
rect 67541 326302 245075 326304
rect 67541 326299 67607 326302
rect 245009 326299 245075 326302
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 109677 325002 109743 325005
rect 119337 325002 119403 325005
rect 252502 325002 252508 325004
rect 109677 325000 252508 325002
rect 109677 324944 109682 325000
rect 109738 324944 119342 325000
rect 119398 324944 252508 325000
rect 109677 324942 252508 324944
rect 109677 324939 109743 324942
rect 119337 324939 119403 324942
rect 252502 324940 252508 324942
rect 252572 324940 252578 325004
rect 83457 323642 83523 323645
rect 92974 323642 92980 323644
rect 83457 323640 92980 323642
rect 83457 323584 83462 323640
rect 83518 323584 92980 323640
rect 83457 323582 92980 323584
rect 83457 323579 83523 323582
rect 92974 323580 92980 323582
rect 93044 323580 93050 323644
rect 102777 323642 102843 323645
rect 141417 323642 141483 323645
rect 102777 323640 141483 323642
rect 102777 323584 102782 323640
rect 102838 323584 141422 323640
rect 141478 323584 141483 323640
rect 102777 323582 141483 323584
rect 102777 323579 102843 323582
rect 141417 323579 141483 323582
rect 76741 322962 76807 322965
rect 82854 322962 82860 322964
rect 76741 322960 82860 322962
rect 76741 322904 76746 322960
rect 76802 322904 82860 322960
rect 76741 322902 82860 322904
rect 76741 322899 76807 322902
rect 82854 322900 82860 322902
rect 82924 322900 82930 322964
rect 92381 322146 92447 322149
rect 104198 322146 104204 322148
rect 92381 322144 104204 322146
rect 92381 322088 92386 322144
rect 92442 322088 104204 322144
rect 92381 322086 104204 322088
rect 92381 322083 92447 322086
rect 104198 322084 104204 322086
rect 104268 322084 104274 322148
rect 106181 322146 106247 322149
rect 124397 322146 124463 322149
rect 125501 322146 125567 322149
rect 106181 322144 125567 322146
rect 106181 322088 106186 322144
rect 106242 322088 124402 322144
rect 124458 322088 125506 322144
rect 125562 322088 125567 322144
rect 106181 322086 125567 322088
rect 106181 322083 106247 322086
rect 124397 322083 124463 322086
rect 125501 322083 125567 322086
rect 43897 321602 43963 321605
rect 265065 321602 265131 321605
rect 43897 321600 265131 321602
rect 43897 321544 43902 321600
rect 43958 321544 265070 321600
rect 265126 321544 265131 321600
rect 43897 321542 265131 321544
rect 43897 321539 43963 321542
rect 265065 321539 265131 321542
rect 97717 321058 97783 321061
rect 108982 321058 108988 321060
rect 97717 321056 108988 321058
rect 97717 321000 97722 321056
rect 97778 321000 108988 321056
rect 97717 320998 108988 321000
rect 97717 320995 97783 320998
rect 108982 320996 108988 320998
rect 109052 320996 109058 321060
rect 85665 320922 85731 320925
rect 97206 320922 97212 320924
rect 85665 320920 97212 320922
rect 85665 320864 85670 320920
rect 85726 320864 97212 320920
rect 85665 320862 97212 320864
rect 85665 320859 85731 320862
rect 97206 320860 97212 320862
rect 97276 320922 97282 320924
rect 118877 320922 118943 320925
rect 97276 320920 118943 320922
rect 97276 320864 118882 320920
rect 118938 320864 118943 320920
rect 97276 320862 118943 320864
rect 97276 320860 97282 320862
rect 118877 320859 118943 320862
rect 77937 320786 78003 320789
rect 120073 320786 120139 320789
rect 262305 320786 262371 320789
rect 77937 320784 262371 320786
rect 77937 320728 77942 320784
rect 77998 320728 120078 320784
rect 120134 320728 262310 320784
rect 262366 320728 262371 320784
rect 77937 320726 262371 320728
rect 77937 320723 78003 320726
rect 120073 320723 120139 320726
rect 262305 320723 262371 320726
rect 191046 320180 191052 320244
rect 191116 320242 191122 320244
rect 201585 320242 201651 320245
rect 191116 320240 201651 320242
rect 191116 320184 201590 320240
rect 201646 320184 201651 320240
rect 191116 320182 201651 320184
rect 191116 320180 191122 320182
rect 201585 320179 201651 320182
rect 81341 319562 81407 319565
rect 114502 319562 114508 319564
rect 81341 319560 114508 319562
rect 81341 319504 81346 319560
rect 81402 319504 114508 319560
rect 81341 319502 114508 319504
rect 81341 319499 81407 319502
rect 114502 319500 114508 319502
rect 114572 319500 114578 319564
rect 72417 319426 72483 319429
rect 79174 319426 79180 319428
rect 72417 319424 79180 319426
rect -960 319290 480 319380
rect 72417 319368 72422 319424
rect 72478 319368 79180 319424
rect 72417 319366 79180 319368
rect 72417 319363 72483 319366
rect 79174 319364 79180 319366
rect 79244 319364 79250 319428
rect 88149 319426 88215 319429
rect 256877 319426 256943 319429
rect 88149 319424 256943 319426
rect 88149 319368 88154 319424
rect 88210 319368 256882 319424
rect 256938 319368 256943 319424
rect 88149 319366 256943 319368
rect 88149 319363 88215 319366
rect 256877 319363 256943 319366
rect 3877 319290 3943 319293
rect -960 319288 3943 319290
rect -960 319232 3882 319288
rect 3938 319232 3943 319288
rect -960 319230 3943 319232
rect -960 319140 480 319230
rect 3877 319227 3943 319230
rect 72601 318882 72667 318885
rect 72734 318882 72740 318884
rect 72601 318880 72740 318882
rect 72601 318824 72606 318880
rect 72662 318824 72740 318880
rect 72601 318822 72740 318824
rect 72601 318819 72667 318822
rect 72734 318820 72740 318822
rect 72804 318882 72810 318884
rect 72969 318882 73035 318885
rect 72804 318880 73035 318882
rect 72804 318824 72974 318880
rect 73030 318824 73035 318880
rect 72804 318822 73035 318824
rect 72804 318820 72810 318822
rect 72969 318819 73035 318822
rect 76649 318746 76715 318749
rect 83406 318746 83412 318748
rect 76649 318744 83412 318746
rect 76649 318688 76654 318744
rect 76710 318688 83412 318744
rect 76649 318686 83412 318688
rect 76649 318683 76715 318686
rect 83406 318684 83412 318686
rect 83476 318684 83482 318748
rect 103421 318202 103487 318205
rect 114737 318202 114803 318205
rect 103421 318200 114803 318202
rect 103421 318144 103426 318200
rect 103482 318144 114742 318200
rect 114798 318144 114803 318200
rect 103421 318142 114803 318144
rect 103421 318139 103487 318142
rect 114737 318139 114803 318142
rect 61837 318066 61903 318069
rect 71681 318066 71747 318069
rect 258390 318066 258396 318068
rect 61837 318064 258396 318066
rect 61837 318008 61842 318064
rect 61898 318008 71686 318064
rect 71742 318008 258396 318064
rect 61837 318006 258396 318008
rect 61837 318003 61903 318006
rect 71681 318003 71747 318006
rect 258390 318004 258396 318006
rect 258460 318004 258466 318068
rect 188337 317522 188403 317525
rect 227713 317522 227779 317525
rect 188337 317520 227779 317522
rect 188337 317464 188342 317520
rect 188398 317464 227718 317520
rect 227774 317464 227779 317520
rect 188337 317462 227779 317464
rect 188337 317459 188403 317462
rect 227713 317459 227779 317462
rect 193765 316298 193831 316301
rect 252686 316298 252692 316300
rect 193765 316296 252692 316298
rect 193765 316240 193770 316296
rect 193826 316240 252692 316296
rect 193765 316238 252692 316240
rect 193765 316235 193831 316238
rect 252686 316236 252692 316238
rect 252756 316236 252762 316300
rect 35801 316162 35867 316165
rect 222193 316162 222259 316165
rect 35801 316160 222259 316162
rect 35801 316104 35806 316160
rect 35862 316104 222198 316160
rect 222254 316104 222259 316160
rect 35801 316102 222259 316104
rect 35801 316099 35867 316102
rect 222193 316099 222259 316102
rect 226977 315346 227043 315349
rect 254526 315346 254532 315348
rect 226977 315344 254532 315346
rect 226977 315288 226982 315344
rect 227038 315288 254532 315344
rect 226977 315286 254532 315288
rect 226977 315283 227043 315286
rect 254526 315284 254532 315286
rect 254596 315284 254602 315348
rect 69105 314938 69171 314941
rect 70301 314938 70367 314941
rect 214557 314938 214623 314941
rect 69105 314936 214623 314938
rect 69105 314880 69110 314936
rect 69166 314880 70306 314936
rect 70362 314880 214562 314936
rect 214618 314880 214623 314936
rect 69105 314878 214623 314880
rect 69105 314875 69171 314878
rect 70301 314875 70367 314878
rect 214557 314875 214623 314878
rect 17217 314802 17283 314805
rect 218513 314802 218579 314805
rect 17217 314800 218579 314802
rect 17217 314744 17222 314800
rect 17278 314744 218518 314800
rect 218574 314744 218579 314800
rect 17217 314742 218579 314744
rect 17217 314739 17283 314742
rect 218513 314739 218579 314742
rect 180149 313442 180215 313445
rect 213177 313442 213243 313445
rect 180149 313440 213243 313442
rect 180149 313384 180154 313440
rect 180210 313384 213182 313440
rect 213238 313384 213243 313440
rect 180149 313382 213243 313384
rect 180149 313379 180215 313382
rect 213177 313379 213243 313382
rect 34421 313306 34487 313309
rect 203241 313306 203307 313309
rect 34421 313304 203307 313306
rect 34421 313248 34426 313304
rect 34482 313248 203246 313304
rect 203302 313248 203307 313304
rect 34421 313246 203307 313248
rect 34421 313243 34487 313246
rect 203241 313243 203307 313246
rect 75821 312490 75887 312493
rect 253933 312490 253999 312493
rect 75821 312488 253999 312490
rect 75821 312432 75826 312488
rect 75882 312432 253938 312488
rect 253994 312432 253999 312488
rect 75821 312430 253999 312432
rect 75821 312427 75887 312430
rect 253933 312427 253999 312430
rect 91185 312082 91251 312085
rect 92381 312082 92447 312085
rect 125593 312082 125659 312085
rect 263777 312082 263843 312085
rect 91185 312080 263843 312082
rect 91185 312024 91190 312080
rect 91246 312024 92386 312080
rect 92442 312024 125598 312080
rect 125654 312024 263782 312080
rect 263838 312024 263843 312080
rect 91185 312022 263843 312024
rect 91185 312019 91251 312022
rect 92381 312019 92447 312022
rect 125593 312019 125659 312022
rect 263777 312019 263843 312022
rect 582373 312082 582439 312085
rect 583520 312082 584960 312172
rect 582373 312080 584960 312082
rect 582373 312024 582378 312080
rect 582434 312024 584960 312080
rect 582373 312022 584960 312024
rect 582373 312019 582439 312022
rect 22737 311946 22803 311949
rect 200297 311946 200363 311949
rect 22737 311944 200363 311946
rect 22737 311888 22742 311944
rect 22798 311888 200302 311944
rect 200358 311888 200363 311944
rect 583520 311932 584960 312022
rect 22737 311886 200363 311888
rect 22737 311883 22803 311886
rect 200297 311883 200363 311886
rect 188521 310858 188587 310861
rect 264094 310858 264100 310860
rect 188521 310856 264100 310858
rect 188521 310800 188526 310856
rect 188582 310800 264100 310856
rect 188521 310798 264100 310800
rect 188521 310795 188587 310798
rect 264094 310796 264100 310798
rect 264164 310796 264170 310860
rect 18597 310722 18663 310725
rect 200389 310722 200455 310725
rect 18597 310720 200455 310722
rect 18597 310664 18602 310720
rect 18658 310664 200394 310720
rect 200450 310664 200455 310720
rect 18597 310662 200455 310664
rect 18597 310659 18663 310662
rect 200389 310659 200455 310662
rect 16481 310586 16547 310589
rect 219617 310586 219683 310589
rect 16481 310584 219683 310586
rect 16481 310528 16486 310584
rect 16542 310528 219622 310584
rect 219678 310528 219683 310584
rect 16481 310526 219683 310528
rect 16481 310523 16547 310526
rect 219617 310523 219683 310526
rect 276013 310450 276079 310453
rect 276657 310450 276723 310453
rect 276013 310448 276723 310450
rect 276013 310392 276018 310448
rect 276074 310392 276662 310448
rect 276718 310392 276723 310448
rect 276013 310390 276723 310392
rect 276013 310387 276079 310390
rect 276657 310387 276723 310390
rect 188337 309498 188403 309501
rect 209773 309498 209839 309501
rect 188337 309496 209839 309498
rect 188337 309440 188342 309496
rect 188398 309440 209778 309496
rect 209834 309440 209839 309496
rect 188337 309438 209839 309440
rect 188337 309435 188403 309438
rect 209773 309435 209839 309438
rect 185669 309362 185735 309365
rect 276013 309362 276079 309365
rect 185669 309360 276079 309362
rect 185669 309304 185674 309360
rect 185730 309304 276018 309360
rect 276074 309304 276079 309360
rect 185669 309302 276079 309304
rect 185669 309299 185735 309302
rect 276013 309299 276079 309302
rect 29637 309226 29703 309229
rect 220813 309226 220879 309229
rect 29637 309224 220879 309226
rect 29637 309168 29642 309224
rect 29698 309168 220818 309224
rect 220874 309168 220879 309224
rect 29637 309166 220879 309168
rect 29637 309163 29703 309166
rect 220813 309163 220879 309166
rect 128445 309090 128511 309093
rect 285673 309090 285739 309093
rect 286317 309090 286383 309093
rect 128445 309088 286383 309090
rect 128445 309032 128450 309088
rect 128506 309032 285678 309088
rect 285734 309032 286322 309088
rect 286378 309032 286383 309088
rect 128445 309030 286383 309032
rect 128445 309027 128511 309030
rect 285673 309027 285739 309030
rect 286317 309027 286383 309030
rect 244917 308954 244983 308957
rect 246205 308954 246271 308957
rect 244917 308952 246271 308954
rect 244917 308896 244922 308952
rect 244978 308896 246210 308952
rect 246266 308896 246271 308952
rect 244917 308894 246271 308896
rect 244917 308891 244983 308894
rect 246205 308891 246271 308894
rect 91001 308410 91067 308413
rect 128445 308410 128511 308413
rect 91001 308408 128511 308410
rect 91001 308352 91006 308408
rect 91062 308352 128450 308408
rect 128506 308352 128511 308408
rect 91001 308350 128511 308352
rect 91001 308347 91067 308350
rect 128445 308347 128511 308350
rect 191373 308002 191439 308005
rect 207749 308002 207815 308005
rect 191373 308000 207815 308002
rect 191373 307944 191378 308000
rect 191434 307944 207754 308000
rect 207810 307944 207815 308000
rect 191373 307942 207815 307944
rect 191373 307939 191439 307942
rect 207749 307939 207815 307942
rect 106774 307804 106780 307868
rect 106844 307866 106850 307868
rect 114645 307866 114711 307869
rect 106844 307864 114711 307866
rect 106844 307808 114650 307864
rect 114706 307808 114711 307864
rect 106844 307806 114711 307808
rect 106844 307804 106850 307806
rect 114645 307803 114711 307806
rect 152457 307866 152523 307869
rect 234613 307866 234679 307869
rect 152457 307864 234679 307866
rect 152457 307808 152462 307864
rect 152518 307808 234618 307864
rect 234674 307808 234679 307864
rect 152457 307806 234679 307808
rect 152457 307803 152523 307806
rect 234613 307803 234679 307806
rect 246205 307866 246271 307869
rect 305637 307866 305703 307869
rect 246205 307864 305703 307866
rect 246205 307808 246210 307864
rect 246266 307808 305642 307864
rect 305698 307808 305703 307864
rect 246205 307806 305703 307808
rect 246205 307803 246271 307806
rect 305637 307803 305703 307806
rect 248413 307050 248479 307053
rect 321553 307050 321619 307053
rect 248413 307048 321619 307050
rect 248413 306992 248418 307048
rect 248474 306992 321558 307048
rect 321614 306992 321619 307048
rect 248413 306990 321619 306992
rect 248413 306987 248479 306990
rect 321553 306987 321619 306990
rect 187049 306778 187115 306781
rect 208393 306778 208459 306781
rect 187049 306776 208459 306778
rect 187049 306720 187054 306776
rect 187110 306720 208398 306776
rect 208454 306720 208459 306776
rect 187049 306718 208459 306720
rect 187049 306715 187115 306718
rect 208393 306715 208459 306718
rect 178769 306642 178835 306645
rect 204253 306642 204319 306645
rect 178769 306640 204319 306642
rect 178769 306584 178774 306640
rect 178830 306584 204258 306640
rect 204314 306584 204319 306640
rect 178769 306582 204319 306584
rect 178769 306579 178835 306582
rect 204253 306579 204319 306582
rect 26141 306506 26207 306509
rect 199653 306506 199719 306509
rect 26141 306504 199719 306506
rect 26141 306448 26146 306504
rect 26202 306448 199658 306504
rect 199714 306448 199719 306504
rect 26141 306446 199719 306448
rect 26141 306443 26207 306446
rect 199653 306443 199719 306446
rect 245653 306506 245719 306509
rect 276657 306506 276723 306509
rect 245653 306504 276723 306506
rect 245653 306448 245658 306504
rect 245714 306448 276662 306504
rect 276718 306448 276723 306504
rect 245653 306446 276723 306448
rect 245653 306443 245719 306446
rect 276657 306443 276723 306446
rect 52177 306370 52243 306373
rect 188521 306370 188587 306373
rect 52177 306368 188587 306370
rect -960 306234 480 306324
rect 52177 306312 52182 306368
rect 52238 306312 188526 306368
rect 188582 306312 188587 306368
rect 52177 306310 188587 306312
rect 52177 306307 52243 306310
rect 188521 306307 188587 306310
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 185577 305146 185643 305149
rect 206001 305146 206067 305149
rect 185577 305144 206067 305146
rect 185577 305088 185582 305144
rect 185638 305088 206006 305144
rect 206062 305088 206067 305144
rect 185577 305086 206067 305088
rect 185577 305083 185643 305086
rect 206001 305083 206067 305086
rect 52177 305010 52243 305013
rect 52310 305010 52316 305012
rect 52177 305008 52316 305010
rect 52177 304952 52182 305008
rect 52238 304952 52316 305008
rect 52177 304950 52316 304952
rect 52177 304947 52243 304950
rect 52310 304948 52316 304950
rect 52380 304948 52386 305012
rect 189809 305010 189875 305013
rect 211889 305010 211955 305013
rect 189809 305008 211955 305010
rect 189809 304952 189814 305008
rect 189870 304952 211894 305008
rect 211950 304952 211955 305008
rect 189809 304950 211955 304952
rect 189809 304947 189875 304950
rect 211889 304947 211955 304950
rect 218646 304948 218652 305012
rect 218716 305010 218722 305012
rect 226977 305010 227043 305013
rect 218716 305008 227043 305010
rect 218716 304952 226982 305008
rect 227038 304952 227043 305008
rect 218716 304950 227043 304952
rect 218716 304948 218722 304950
rect 226977 304947 227043 304950
rect 242157 305010 242223 305013
rect 277393 305010 277459 305013
rect 242157 305008 277459 305010
rect 242157 304952 242162 305008
rect 242218 304952 277398 305008
rect 277454 304952 277459 305008
rect 242157 304950 277459 304952
rect 242157 304947 242223 304950
rect 277393 304947 277459 304950
rect 79869 304194 79935 304197
rect 87270 304194 87276 304196
rect 79869 304192 87276 304194
rect 79869 304136 79874 304192
rect 79930 304136 87276 304192
rect 79869 304134 87276 304136
rect 79869 304131 79935 304134
rect 87270 304132 87276 304134
rect 87340 304132 87346 304196
rect 93669 304194 93735 304197
rect 104249 304194 104315 304197
rect 93669 304192 104315 304194
rect 93669 304136 93674 304192
rect 93730 304136 104254 304192
rect 104310 304136 104315 304192
rect 93669 304134 104315 304136
rect 93669 304131 93735 304134
rect 104249 304131 104315 304134
rect 104433 304194 104499 304197
rect 121637 304194 121703 304197
rect 104433 304192 121703 304194
rect 104433 304136 104438 304192
rect 104494 304136 121642 304192
rect 121698 304136 121703 304192
rect 104433 304134 121703 304136
rect 104433 304131 104499 304134
rect 121637 304131 121703 304134
rect 247677 304194 247743 304197
rect 253197 304194 253263 304197
rect 247677 304192 253263 304194
rect 247677 304136 247682 304192
rect 247738 304136 253202 304192
rect 253258 304136 253263 304192
rect 247677 304134 253263 304136
rect 247677 304131 247743 304134
rect 253197 304131 253263 304134
rect 186814 303860 186820 303924
rect 186884 303922 186890 303924
rect 195513 303922 195579 303925
rect 186884 303920 195579 303922
rect 186884 303864 195518 303920
rect 195574 303864 195579 303920
rect 186884 303862 195579 303864
rect 186884 303860 186890 303862
rect 195513 303859 195579 303862
rect 238661 303922 238727 303925
rect 242014 303922 242020 303924
rect 238661 303920 242020 303922
rect 238661 303864 238666 303920
rect 238722 303864 242020 303920
rect 238661 303862 242020 303864
rect 238661 303859 238727 303862
rect 242014 303860 242020 303862
rect 242084 303860 242090 303924
rect 215886 303724 215892 303788
rect 215956 303786 215962 303788
rect 229369 303786 229435 303789
rect 215956 303784 229435 303786
rect 215956 303728 229374 303784
rect 229430 303728 229435 303784
rect 215956 303726 229435 303728
rect 215956 303724 215962 303726
rect 229369 303723 229435 303726
rect 250897 303786 250963 303789
rect 260230 303786 260236 303788
rect 250897 303784 260236 303786
rect 250897 303728 250902 303784
rect 250958 303728 260236 303784
rect 250897 303726 260236 303728
rect 250897 303723 250963 303726
rect 260230 303724 260236 303726
rect 260300 303724 260306 303788
rect 192702 303588 192708 303652
rect 192772 303650 192778 303652
rect 197905 303650 197971 303653
rect 192772 303648 197971 303650
rect 192772 303592 197910 303648
rect 197966 303592 197971 303648
rect 192772 303590 197971 303592
rect 192772 303588 192778 303590
rect 197905 303587 197971 303590
rect 230473 303650 230539 303653
rect 237782 303650 237788 303652
rect 230473 303648 237788 303650
rect 230473 303592 230478 303648
rect 230534 303592 237788 303648
rect 230473 303590 237788 303592
rect 230473 303587 230539 303590
rect 237782 303588 237788 303590
rect 237852 303588 237858 303652
rect 249701 303650 249767 303653
rect 260046 303650 260052 303652
rect 249701 303648 260052 303650
rect 249701 303592 249706 303648
rect 249762 303592 260052 303648
rect 249701 303590 260052 303592
rect 249701 303587 249767 303590
rect 260046 303588 260052 303590
rect 260116 303588 260122 303652
rect 248873 302834 248939 302837
rect 249793 302834 249859 302837
rect 295977 302834 296043 302837
rect 248873 302832 296043 302834
rect 248873 302776 248878 302832
rect 248934 302776 249798 302832
rect 249854 302776 295982 302832
rect 296038 302776 296043 302832
rect 248873 302774 296043 302776
rect 248873 302771 248939 302774
rect 249793 302771 249859 302774
rect 295977 302771 296043 302774
rect 151077 302562 151143 302565
rect 246849 302562 246915 302565
rect 151077 302560 246915 302562
rect 151077 302504 151082 302560
rect 151138 302504 246854 302560
rect 246910 302504 246915 302560
rect 151077 302502 246915 302504
rect 151077 302499 151143 302502
rect 246849 302499 246915 302502
rect 191281 302426 191347 302429
rect 252645 302426 252711 302429
rect 191281 302424 252711 302426
rect 191281 302368 191286 302424
rect 191342 302368 252650 302424
rect 252706 302368 252711 302424
rect 191281 302366 252711 302368
rect 191281 302363 191347 302366
rect 252645 302363 252711 302366
rect 238017 302290 238083 302293
rect 240358 302290 240364 302292
rect 238017 302288 240364 302290
rect 238017 302232 238022 302288
rect 238078 302232 240364 302288
rect 238017 302230 240364 302232
rect 238017 302227 238083 302230
rect 240358 302228 240364 302230
rect 240428 302228 240434 302292
rect 246849 302290 246915 302293
rect 327073 302290 327139 302293
rect 246849 302288 327139 302290
rect 246849 302232 246854 302288
rect 246910 302232 327078 302288
rect 327134 302232 327139 302288
rect 246849 302230 327139 302232
rect 246849 302227 246915 302230
rect 327073 302227 327139 302230
rect 192569 301746 192635 301749
rect 197537 301746 197603 301749
rect 192569 301744 197603 301746
rect 192569 301688 192574 301744
rect 192630 301688 197542 301744
rect 197598 301688 197603 301744
rect 192569 301686 197603 301688
rect 192569 301683 192635 301686
rect 197537 301683 197603 301686
rect 250345 301746 250411 301749
rect 345013 301746 345079 301749
rect 250345 301744 345079 301746
rect 250345 301688 250350 301744
rect 250406 301688 345018 301744
rect 345074 301688 345079 301744
rect 250345 301686 345079 301688
rect 250345 301683 250411 301686
rect 345013 301683 345079 301686
rect 178677 301610 178743 301613
rect 247769 301610 247835 301613
rect 178677 301608 247835 301610
rect 178677 301552 178682 301608
rect 178738 301552 247774 301608
rect 247830 301552 247835 301608
rect 178677 301550 247835 301552
rect 178677 301547 178743 301550
rect 247769 301547 247835 301550
rect 253289 301610 253355 301613
rect 254158 301610 254164 301612
rect 253289 301608 254164 301610
rect 253289 301552 253294 301608
rect 253350 301552 254164 301608
rect 253289 301550 254164 301552
rect 253289 301547 253355 301550
rect 254158 301548 254164 301550
rect 254228 301548 254234 301612
rect 75821 301474 75887 301477
rect 186313 301474 186379 301477
rect 75821 301472 186379 301474
rect 75821 301416 75826 301472
rect 75882 301416 186318 301472
rect 186374 301416 186379 301472
rect 75821 301414 186379 301416
rect 75821 301411 75887 301414
rect 186313 301411 186379 301414
rect 193438 301412 193444 301476
rect 193508 301474 193514 301476
rect 194225 301474 194291 301477
rect 193508 301472 194291 301474
rect 193508 301416 194230 301472
rect 194286 301416 194291 301472
rect 193508 301414 194291 301416
rect 193508 301412 193514 301414
rect 194225 301411 194291 301414
rect 197537 301474 197603 301477
rect 244825 301474 244891 301477
rect 197537 301472 244891 301474
rect 197537 301416 197542 301472
rect 197598 301416 244830 301472
rect 244886 301416 244891 301472
rect 197537 301414 244891 301416
rect 197537 301411 197603 301414
rect 244825 301411 244891 301414
rect 246481 301474 246547 301477
rect 253473 301474 253539 301477
rect 246481 301472 253539 301474
rect 246481 301416 246486 301472
rect 246542 301416 253478 301472
rect 253534 301416 253539 301472
rect 246481 301414 253539 301416
rect 246481 301411 246547 301414
rect 253473 301411 253539 301414
rect 188429 301338 188495 301341
rect 251817 301338 251883 301341
rect 188429 301336 251883 301338
rect 188429 301280 188434 301336
rect 188490 301280 251822 301336
rect 251878 301280 251883 301336
rect 188429 301278 251883 301280
rect 188429 301275 188495 301278
rect 251817 301275 251883 301278
rect 193254 301140 193260 301204
rect 193324 301202 193330 301204
rect 194501 301202 194567 301205
rect 193324 301200 194567 301202
rect 193324 301144 194506 301200
rect 194562 301144 194567 301200
rect 193324 301142 194567 301144
rect 193324 301140 193330 301142
rect 194501 301139 194567 301142
rect 210366 301140 210372 301204
rect 210436 301202 210442 301204
rect 212809 301202 212875 301205
rect 210436 301200 212875 301202
rect 210436 301144 212814 301200
rect 212870 301144 212875 301200
rect 210436 301142 212875 301144
rect 210436 301140 210442 301142
rect 212809 301139 212875 301142
rect 222694 301140 222700 301204
rect 222764 301202 222770 301204
rect 224953 301202 225019 301205
rect 258574 301202 258580 301204
rect 222764 301200 225019 301202
rect 222764 301144 224958 301200
rect 225014 301144 225019 301200
rect 222764 301142 225019 301144
rect 253460 301142 258580 301202
rect 222764 301140 222770 301142
rect 224953 301139 225019 301142
rect 258574 301140 258580 301142
rect 258644 301140 258650 301204
rect 208894 301004 208900 301068
rect 208964 301066 208970 301068
rect 210417 301066 210483 301069
rect 208964 301064 210483 301066
rect 208964 301008 210422 301064
rect 210478 301008 210483 301064
rect 208964 301006 210483 301008
rect 208964 301004 208970 301006
rect 210417 301003 210483 301006
rect 213678 301004 213684 301068
rect 213748 301066 213754 301068
rect 216305 301066 216371 301069
rect 213748 301064 216371 301066
rect 213748 301008 216310 301064
rect 216366 301008 216371 301064
rect 213748 301006 216371 301008
rect 213748 301004 213754 301006
rect 216305 301003 216371 301006
rect 219382 301004 219388 301068
rect 219452 301066 219458 301068
rect 220353 301066 220419 301069
rect 219452 301064 220419 301066
rect 219452 301008 220358 301064
rect 220414 301008 220419 301064
rect 219452 301006 220419 301008
rect 219452 301004 219458 301006
rect 220353 301003 220419 301006
rect 221222 301004 221228 301068
rect 221292 301066 221298 301068
rect 222745 301066 222811 301069
rect 221292 301064 222811 301066
rect 221292 301008 222750 301064
rect 222806 301008 222811 301064
rect 221292 301006 222811 301008
rect 221292 301004 221298 301006
rect 222745 301003 222811 301006
rect 223798 301004 223804 301068
rect 223868 301066 223874 301068
rect 224401 301066 224467 301069
rect 223868 301064 224467 301066
rect 223868 301008 224406 301064
rect 224462 301008 224467 301064
rect 223868 301006 224467 301008
rect 223868 301004 223874 301006
rect 224401 301003 224467 301006
rect 230422 301004 230428 301068
rect 230492 301066 230498 301068
rect 231393 301066 231459 301069
rect 230492 301064 231459 301066
rect 230492 301008 231398 301064
rect 231454 301008 231459 301064
rect 230492 301006 231459 301008
rect 230492 301004 230498 301006
rect 231393 301003 231459 301006
rect 232078 301004 232084 301068
rect 232148 301066 232154 301068
rect 232589 301066 232655 301069
rect 232148 301064 232655 301066
rect 232148 301008 232594 301064
rect 232650 301008 232655 301064
rect 232148 301006 232655 301008
rect 232148 301004 232154 301006
rect 232589 301003 232655 301006
rect 233182 301004 233188 301068
rect 233252 301066 233258 301068
rect 233785 301066 233851 301069
rect 233252 301064 233851 301066
rect 233252 301008 233790 301064
rect 233846 301008 233851 301064
rect 233252 301006 233851 301008
rect 233252 301004 233258 301006
rect 233785 301003 233851 301006
rect 234838 301004 234844 301068
rect 234908 301066 234914 301068
rect 235441 301066 235507 301069
rect 234908 301064 235507 301066
rect 234908 301008 235446 301064
rect 235502 301008 235507 301064
rect 234908 301006 235507 301008
rect 234908 301004 234914 301006
rect 235441 301003 235507 301006
rect 191189 300930 191255 300933
rect 196065 300932 196131 300933
rect 196014 300930 196020 300932
rect 191189 300928 193660 300930
rect 191189 300872 191194 300928
rect 191250 300872 193660 300928
rect 191189 300870 193660 300872
rect 195974 300870 196020 300930
rect 196084 300928 196131 300932
rect 196126 300872 196131 300928
rect 191189 300867 191255 300870
rect 196014 300868 196020 300870
rect 196084 300868 196131 300872
rect 197486 300868 197492 300932
rect 197556 300930 197562 300932
rect 198181 300930 198247 300933
rect 198825 300932 198891 300933
rect 198774 300930 198780 300932
rect 197556 300928 198247 300930
rect 197556 300872 198186 300928
rect 198242 300872 198247 300928
rect 197556 300870 198247 300872
rect 198734 300870 198780 300930
rect 198844 300928 198891 300932
rect 198886 300872 198891 300928
rect 197556 300868 197562 300870
rect 196065 300867 196131 300868
rect 198181 300867 198247 300870
rect 198774 300868 198780 300870
rect 198844 300868 198891 300872
rect 201534 300868 201540 300932
rect 201604 300930 201610 300932
rect 202321 300930 202387 300933
rect 203057 300932 203123 300933
rect 203006 300930 203012 300932
rect 201604 300928 202387 300930
rect 201604 300872 202326 300928
rect 202382 300872 202387 300928
rect 201604 300870 202387 300872
rect 202966 300870 203012 300930
rect 203076 300928 203123 300932
rect 203118 300872 203123 300928
rect 201604 300868 201610 300870
rect 198825 300867 198891 300868
rect 202321 300867 202387 300870
rect 203006 300868 203012 300870
rect 203076 300868 203123 300872
rect 204294 300868 204300 300932
rect 204364 300930 204370 300932
rect 204621 300930 204687 300933
rect 204364 300928 204687 300930
rect 204364 300872 204626 300928
rect 204682 300872 204687 300928
rect 204364 300870 204687 300872
rect 204364 300868 204370 300870
rect 203057 300867 203123 300868
rect 204621 300867 204687 300870
rect 205582 300868 205588 300932
rect 205652 300930 205658 300932
rect 206277 300930 206343 300933
rect 207105 300932 207171 300933
rect 207054 300930 207060 300932
rect 205652 300928 206343 300930
rect 205652 300872 206282 300928
rect 206338 300872 206343 300928
rect 205652 300870 206343 300872
rect 207014 300870 207060 300930
rect 207124 300928 207171 300932
rect 207166 300872 207171 300928
rect 205652 300868 205658 300870
rect 206277 300867 206343 300870
rect 207054 300868 207060 300870
rect 207124 300868 207171 300872
rect 208342 300868 208348 300932
rect 208412 300930 208418 300932
rect 209313 300930 209379 300933
rect 208412 300928 209379 300930
rect 208412 300872 209318 300928
rect 209374 300872 209379 300928
rect 208412 300870 209379 300872
rect 208412 300868 208418 300870
rect 207105 300867 207171 300868
rect 209313 300867 209379 300870
rect 211654 300868 211660 300932
rect 211724 300930 211730 300932
rect 212165 300930 212231 300933
rect 211724 300928 212231 300930
rect 211724 300872 212170 300928
rect 212226 300872 212231 300928
rect 211724 300870 212231 300872
rect 211724 300868 211730 300870
rect 212165 300867 212231 300870
rect 213862 300868 213868 300932
rect 213932 300930 213938 300932
rect 214281 300930 214347 300933
rect 213932 300928 214347 300930
rect 213932 300872 214286 300928
rect 214342 300872 214347 300928
rect 213932 300870 214347 300872
rect 213932 300868 213938 300870
rect 214281 300867 214347 300870
rect 214414 300868 214420 300932
rect 214484 300930 214490 300932
rect 215109 300930 215175 300933
rect 214484 300928 215175 300930
rect 214484 300872 215114 300928
rect 215170 300872 215175 300928
rect 214484 300870 215175 300872
rect 214484 300868 214490 300870
rect 215109 300867 215175 300870
rect 216070 300868 216076 300932
rect 216140 300930 216146 300932
rect 216673 300930 216739 300933
rect 216140 300928 216739 300930
rect 216140 300872 216678 300928
rect 216734 300872 216739 300928
rect 216140 300870 216739 300872
rect 216140 300868 216146 300870
rect 216673 300867 216739 300870
rect 216806 300868 216812 300932
rect 216876 300930 216882 300932
rect 217317 300930 217383 300933
rect 216876 300928 217383 300930
rect 216876 300872 217322 300928
rect 217378 300872 217383 300928
rect 216876 300870 217383 300872
rect 216876 300868 216882 300870
rect 217317 300867 217383 300870
rect 219525 300932 219591 300933
rect 219525 300928 219572 300932
rect 219636 300930 219642 300932
rect 219525 300872 219530 300928
rect 219525 300868 219572 300872
rect 219636 300870 219682 300930
rect 219636 300868 219642 300870
rect 220854 300868 220860 300932
rect 220924 300930 220930 300932
rect 221457 300930 221523 300933
rect 220924 300928 221523 300930
rect 220924 300872 221462 300928
rect 221518 300872 221523 300928
rect 220924 300870 221523 300872
rect 220924 300868 220930 300870
rect 219525 300867 219591 300868
rect 221457 300867 221523 300870
rect 222326 300868 222332 300932
rect 222396 300930 222402 300932
rect 223205 300930 223271 300933
rect 224033 300932 224099 300933
rect 223982 300930 223988 300932
rect 222396 300928 223271 300930
rect 222396 300872 223210 300928
rect 223266 300872 223271 300928
rect 222396 300870 223271 300872
rect 223942 300870 223988 300930
rect 224052 300928 224099 300932
rect 224094 300872 224099 300928
rect 222396 300868 222402 300870
rect 223205 300867 223271 300870
rect 223982 300868 223988 300870
rect 224052 300868 224099 300872
rect 225086 300868 225092 300932
rect 225156 300930 225162 300932
rect 225597 300930 225663 300933
rect 225156 300928 225663 300930
rect 225156 300872 225602 300928
rect 225658 300872 225663 300928
rect 225156 300870 225663 300872
rect 225156 300868 225162 300870
rect 224033 300867 224099 300868
rect 225597 300867 225663 300870
rect 226333 300932 226399 300933
rect 226333 300928 226380 300932
rect 226444 300930 226450 300932
rect 226333 300872 226338 300928
rect 226333 300868 226380 300872
rect 226444 300870 226490 300930
rect 226444 300868 226450 300870
rect 226558 300868 226564 300932
rect 226628 300930 226634 300932
rect 227253 300930 227319 300933
rect 226628 300928 227319 300930
rect 226628 300872 227258 300928
rect 227314 300872 227319 300928
rect 226628 300870 227319 300872
rect 226628 300868 226634 300870
rect 226333 300867 226399 300868
rect 227253 300867 227319 300870
rect 227662 300868 227668 300932
rect 227732 300930 227738 300932
rect 228449 300930 228515 300933
rect 229737 300932 229803 300933
rect 231025 300932 231091 300933
rect 232313 300932 232379 300933
rect 229686 300930 229692 300932
rect 227732 300928 228515 300930
rect 227732 300872 228454 300928
rect 228510 300872 228515 300928
rect 227732 300870 228515 300872
rect 229646 300870 229692 300930
rect 229756 300928 229803 300932
rect 230974 300930 230980 300932
rect 229798 300872 229803 300928
rect 227732 300868 227738 300870
rect 228449 300867 228515 300870
rect 229686 300868 229692 300870
rect 229756 300868 229803 300872
rect 230934 300870 230980 300930
rect 231044 300928 231091 300932
rect 232262 300930 232268 300932
rect 231086 300872 231091 300928
rect 230974 300868 230980 300870
rect 231044 300868 231091 300872
rect 232222 300870 232268 300930
rect 232332 300928 232379 300932
rect 232374 300872 232379 300928
rect 232262 300868 232268 300870
rect 232332 300868 232379 300872
rect 229737 300867 229803 300868
rect 231025 300867 231091 300868
rect 232313 300867 232379 300868
rect 233325 300932 233391 300933
rect 233325 300928 233372 300932
rect 233436 300930 233442 300932
rect 233325 300872 233330 300928
rect 233325 300868 233372 300872
rect 233436 300870 233482 300930
rect 233436 300868 233442 300870
rect 234654 300868 234660 300932
rect 234724 300930 234730 300932
rect 234889 300930 234955 300933
rect 234724 300928 234955 300930
rect 234724 300872 234894 300928
rect 234950 300872 234955 300928
rect 234724 300870 234955 300872
rect 234724 300868 234730 300870
rect 233325 300867 233391 300868
rect 234889 300867 234955 300870
rect 236494 300868 236500 300932
rect 236564 300930 236570 300932
rect 236729 300930 236795 300933
rect 236564 300928 236795 300930
rect 236564 300872 236734 300928
rect 236790 300872 236795 300928
rect 236564 300870 236795 300872
rect 236564 300868 236570 300870
rect 236729 300867 236795 300870
rect 237833 300930 237899 300933
rect 238150 300930 238156 300932
rect 237833 300928 238156 300930
rect 237833 300872 237838 300928
rect 237894 300872 238156 300928
rect 237833 300870 238156 300872
rect 237833 300867 237899 300870
rect 238150 300868 238156 300870
rect 238220 300868 238226 300932
rect 238702 300868 238708 300932
rect 238772 300930 238778 300932
rect 238845 300930 238911 300933
rect 238772 300928 238911 300930
rect 238772 300872 238850 300928
rect 238906 300872 238911 300928
rect 238772 300870 238911 300872
rect 238772 300868 238778 300870
rect 238845 300867 238911 300870
rect 240041 300930 240107 300933
rect 244406 300930 244412 300932
rect 240041 300928 244412 300930
rect 240041 300872 240046 300928
rect 240102 300872 244412 300928
rect 240041 300870 244412 300872
rect 240041 300867 240107 300870
rect 244406 300868 244412 300870
rect 244476 300868 244482 300932
rect 255681 300794 255747 300797
rect 253460 300792 255747 300794
rect 253460 300736 255686 300792
rect 255742 300736 255747 300792
rect 253460 300734 255747 300736
rect 255681 300731 255747 300734
rect 253197 300522 253263 300525
rect 324957 300522 325023 300525
rect 253197 300520 325023 300522
rect 253197 300464 253202 300520
rect 253258 300464 324962 300520
rect 325018 300464 325023 300520
rect 253197 300462 325023 300464
rect 253197 300459 253263 300462
rect 324957 300459 325023 300462
rect 73245 300250 73311 300253
rect 73797 300250 73863 300253
rect 193673 300250 193739 300253
rect 254526 300250 254532 300252
rect 73245 300248 193739 300250
rect 73245 300192 73250 300248
rect 73306 300192 73802 300248
rect 73858 300192 193678 300248
rect 193734 300192 193739 300248
rect 73245 300190 193739 300192
rect 253460 300190 254532 300250
rect 73245 300187 73311 300190
rect 73797 300187 73863 300190
rect 193673 300187 193739 300190
rect 254526 300188 254532 300190
rect 254596 300250 254602 300252
rect 255865 300250 255931 300253
rect 254596 300248 255931 300250
rect 254596 300192 255870 300248
rect 255926 300192 255931 300248
rect 254596 300190 255931 300192
rect 254596 300188 254602 300190
rect 255865 300187 255931 300190
rect 191097 299978 191163 299981
rect 191097 299976 193660 299978
rect 191097 299920 191102 299976
rect 191158 299920 193660 299976
rect 191097 299918 193660 299920
rect 191097 299915 191163 299918
rect 255446 299842 255452 299844
rect 253460 299782 255452 299842
rect 255446 299780 255452 299782
rect 255516 299780 255522 299844
rect 255681 299434 255747 299437
rect 253460 299432 255747 299434
rect 253460 299376 255686 299432
rect 255742 299376 255747 299432
rect 253460 299374 255747 299376
rect 255681 299371 255747 299374
rect 191741 299026 191807 299029
rect 191741 299024 193660 299026
rect 191741 298968 191746 299024
rect 191802 298968 193660 299024
rect 191741 298966 193660 298968
rect 191741 298963 191807 298966
rect 166349 298890 166415 298893
rect 193438 298890 193444 298892
rect 166349 298888 193444 298890
rect 166349 298832 166354 298888
rect 166410 298832 193444 298888
rect 166349 298830 193444 298832
rect 166349 298827 166415 298830
rect 193438 298828 193444 298830
rect 193508 298828 193514 298892
rect 255773 298890 255839 298893
rect 253460 298888 255839 298890
rect 253460 298832 255778 298888
rect 255834 298832 255839 298888
rect 253460 298830 255839 298832
rect 255773 298827 255839 298830
rect 22001 298754 22067 298757
rect 191046 298754 191052 298756
rect 22001 298752 191052 298754
rect 22001 298696 22006 298752
rect 22062 298696 191052 298752
rect 22001 298694 191052 298696
rect 22001 298691 22067 298694
rect 191046 298692 191052 298694
rect 191116 298692 191122 298756
rect 253473 298754 253539 298757
rect 253430 298752 253539 298754
rect 253430 298696 253478 298752
rect 253534 298696 253539 298752
rect 253430 298691 253539 298696
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 253430 298482 253490 298691
rect 583520 298604 584960 298694
rect 255262 298482 255268 298484
rect 253430 298452 255268 298482
rect 253460 298422 255268 298452
rect 255262 298420 255268 298422
rect 255332 298420 255338 298484
rect 255681 298074 255747 298077
rect 253460 298072 255747 298074
rect 191465 297530 191531 297533
rect 193630 297530 193690 298044
rect 253460 298016 255686 298072
rect 255742 298016 255747 298072
rect 253460 298014 255747 298016
rect 255681 298011 255747 298014
rect 252870 297876 252876 297940
rect 252940 297876 252946 297940
rect 191465 297528 193690 297530
rect 191465 297472 191470 297528
rect 191526 297472 193690 297528
rect 252878 297530 252938 297876
rect 284293 297530 284359 297533
rect 252878 297528 284359 297530
rect 252878 297500 284298 297528
rect 191465 297470 193690 297472
rect 252908 297472 284298 297500
rect 284354 297472 284359 297528
rect 252908 297470 284359 297472
rect 191465 297467 191531 297470
rect 284293 297467 284359 297470
rect 262121 297394 262187 297397
rect 262397 297394 262463 297397
rect 280797 297394 280863 297397
rect 262121 297392 280863 297394
rect 262121 297336 262126 297392
rect 262182 297336 262402 297392
rect 262458 297336 280802 297392
rect 280858 297336 280863 297392
rect 262121 297334 280863 297336
rect 262121 297331 262187 297334
rect 262397 297331 262463 297334
rect 280797 297331 280863 297334
rect 255773 297122 255839 297125
rect 253460 297120 255839 297122
rect 67766 296924 67772 296988
rect 67836 296986 67842 296988
rect 193630 296986 193690 297092
rect 253460 297064 255778 297120
rect 255834 297064 255839 297120
rect 253460 297062 255839 297064
rect 255773 297059 255839 297062
rect 67836 296926 193690 296986
rect 67836 296924 67842 296926
rect 61878 296788 61884 296852
rect 61948 296850 61954 296852
rect 191465 296850 191531 296853
rect 61948 296848 191531 296850
rect 61948 296792 191470 296848
rect 191526 296792 191531 296848
rect 61948 296790 191531 296792
rect 61948 296788 61954 296790
rect 191465 296787 191531 296790
rect 255681 296578 255747 296581
rect 253460 296576 255747 296578
rect 253460 296520 255686 296576
rect 255742 296520 255747 296576
rect 253460 296518 255747 296520
rect 255681 296515 255747 296518
rect 191741 296170 191807 296173
rect 191741 296168 193660 296170
rect 191741 296112 191746 296168
rect 191802 296112 193660 296168
rect 191741 296110 193660 296112
rect 191741 296107 191807 296110
rect 253430 296034 253490 296140
rect 261477 296034 261543 296037
rect 253430 296032 261543 296034
rect 253430 295976 261482 296032
rect 261538 295976 261543 296032
rect 253430 295974 261543 295976
rect 261477 295971 261543 295974
rect 255405 295762 255471 295765
rect 253460 295760 255471 295762
rect 253460 295704 255410 295760
rect 255466 295704 255471 295760
rect 253460 295702 255471 295704
rect 255405 295699 255471 295702
rect 61929 295354 61995 295357
rect 179413 295354 179479 295357
rect 61929 295352 179479 295354
rect 61929 295296 61934 295352
rect 61990 295296 179418 295352
rect 179474 295296 179479 295352
rect 61929 295294 179479 295296
rect 61929 295291 61995 295294
rect 179413 295291 179479 295294
rect 256785 295218 256851 295221
rect 253460 295216 256851 295218
rect 193630 294538 193690 295188
rect 253460 295160 256790 295216
rect 256846 295160 256851 295216
rect 253460 295158 256851 295160
rect 256785 295155 256851 295158
rect 255405 294810 255471 294813
rect 253460 294808 255471 294810
rect 253460 294752 255410 294808
rect 255466 294752 255471 294808
rect 253460 294750 255471 294752
rect 255405 294747 255471 294750
rect 180750 294478 193690 294538
rect 65885 294130 65951 294133
rect 180750 294130 180810 294478
rect 255262 294476 255268 294540
rect 255332 294538 255338 294540
rect 299473 294538 299539 294541
rect 255332 294536 299539 294538
rect 255332 294480 299478 294536
rect 299534 294480 299539 294536
rect 255332 294478 299539 294480
rect 255332 294476 255338 294478
rect 299473 294475 299539 294478
rect 255446 294402 255452 294404
rect 253460 294342 255452 294402
rect 255446 294340 255452 294342
rect 255516 294340 255522 294404
rect 191649 294266 191715 294269
rect 191649 294264 193660 294266
rect 191649 294208 191654 294264
rect 191710 294208 193660 294264
rect 191649 294206 193660 294208
rect 191649 294203 191715 294206
rect 65885 294128 180810 294130
rect 65885 294072 65890 294128
rect 65946 294072 180810 294128
rect 65885 294070 180810 294072
rect 65885 294067 65951 294070
rect 255814 293858 255820 293860
rect 253460 293798 255820 293858
rect 255814 293796 255820 293798
rect 255884 293796 255890 293860
rect 255405 293450 255471 293453
rect 253460 293448 255471 293450
rect 253460 293392 255410 293448
rect 255466 293392 255471 293448
rect 253460 293390 255471 293392
rect 255405 293387 255471 293390
rect -960 293178 480 293268
rect 3509 293178 3575 293181
rect -960 293176 3575 293178
rect -960 293120 3514 293176
rect 3570 293120 3575 293176
rect -960 293118 3575 293120
rect -960 293028 480 293118
rect 3509 293115 3575 293118
rect 191741 293178 191807 293181
rect 191741 293176 193660 293178
rect 191741 293120 191746 293176
rect 191802 293120 193660 293176
rect 191741 293118 193660 293120
rect 191741 293115 191807 293118
rect 255446 293116 255452 293180
rect 255516 293178 255522 293180
rect 582925 293178 582991 293181
rect 255516 293176 582991 293178
rect 255516 293120 582930 293176
rect 582986 293120 582991 293176
rect 255516 293118 582991 293120
rect 255516 293116 255522 293118
rect 582925 293115 582991 293118
rect 255681 293042 255747 293045
rect 253460 293040 255747 293042
rect 253460 292984 255686 293040
rect 255742 292984 255747 293040
rect 253460 292982 255747 292984
rect 255681 292979 255747 292982
rect 103830 292770 103836 292772
rect 84150 292710 103836 292770
rect 78765 292634 78831 292637
rect 79869 292634 79935 292637
rect 84150 292634 84210 292710
rect 103830 292708 103836 292710
rect 103900 292708 103906 292772
rect 78765 292632 84210 292634
rect 78765 292576 78770 292632
rect 78826 292576 79874 292632
rect 79930 292576 84210 292632
rect 78765 292574 84210 292576
rect 89713 292634 89779 292637
rect 90950 292634 90956 292636
rect 89713 292632 90956 292634
rect 89713 292576 89718 292632
rect 89774 292576 90956 292632
rect 89713 292574 90956 292576
rect 78765 292571 78831 292574
rect 79869 292571 79935 292574
rect 89713 292571 89779 292574
rect 90950 292572 90956 292574
rect 91020 292634 91026 292636
rect 122097 292634 122163 292637
rect 91020 292632 122163 292634
rect 91020 292576 122102 292632
rect 122158 292576 122163 292632
rect 91020 292574 122163 292576
rect 91020 292572 91026 292574
rect 122097 292571 122163 292574
rect 254025 292498 254091 292501
rect 253460 292496 254091 292498
rect 253460 292440 254030 292496
rect 254086 292440 254091 292496
rect 253460 292438 254091 292440
rect 254025 292435 254091 292438
rect 191189 292226 191255 292229
rect 191189 292224 193660 292226
rect 191189 292168 191194 292224
rect 191250 292168 193660 292224
rect 191189 292166 193660 292168
rect 191189 292163 191255 292166
rect 255405 292090 255471 292093
rect 253460 292088 255471 292090
rect 253460 292032 255410 292088
rect 255466 292032 255471 292088
rect 253460 292030 255471 292032
rect 255405 292027 255471 292030
rect 116025 291818 116091 291821
rect 116526 291818 116532 291820
rect 116025 291816 116532 291818
rect 116025 291760 116030 291816
rect 116086 291760 116532 291816
rect 116025 291758 116532 291760
rect 116025 291755 116091 291758
rect 116526 291756 116532 291758
rect 116596 291756 116602 291820
rect 166257 291818 166323 291821
rect 191373 291818 191439 291821
rect 166257 291816 191439 291818
rect 166257 291760 166262 291816
rect 166318 291760 191378 291816
rect 191434 291760 191439 291816
rect 166257 291758 191439 291760
rect 166257 291755 166323 291758
rect 191373 291755 191439 291758
rect 255773 291546 255839 291549
rect 253460 291544 255839 291546
rect 253460 291488 255778 291544
rect 255834 291488 255839 291544
rect 253460 291486 255839 291488
rect 255773 291483 255839 291486
rect 85481 291410 85547 291413
rect 100150 291410 100156 291412
rect 85481 291408 100156 291410
rect 85481 291352 85486 291408
rect 85542 291352 100156 291408
rect 85481 291350 100156 291352
rect 85481 291347 85547 291350
rect 100150 291348 100156 291350
rect 100220 291348 100226 291412
rect 252870 291348 252876 291412
rect 252940 291348 252946 291412
rect 88057 291274 88123 291277
rect 121637 291274 121703 291277
rect 88057 291272 121703 291274
rect 88057 291216 88062 291272
rect 88118 291216 121642 291272
rect 121698 291216 121703 291272
rect 88057 291214 121703 291216
rect 88057 291211 88123 291214
rect 121637 291211 121703 291214
rect 191649 291274 191715 291277
rect 191649 291272 193660 291274
rect 191649 291216 191654 291272
rect 191710 291216 193660 291272
rect 191649 291214 193660 291216
rect 191649 291211 191715 291214
rect 252878 291108 252938 291348
rect 255405 290730 255471 290733
rect 253460 290728 255471 290730
rect 253460 290672 255410 290728
rect 255466 290672 255471 290728
rect 253460 290670 255471 290672
rect 255405 290667 255471 290670
rect 191741 290322 191807 290325
rect 191741 290320 193660 290322
rect 191741 290264 191746 290320
rect 191802 290264 193660 290320
rect 191741 290262 193660 290264
rect 191741 290259 191807 290262
rect 255681 290186 255747 290189
rect 253460 290184 255747 290186
rect 253460 290128 255686 290184
rect 255742 290128 255747 290184
rect 253460 290126 255747 290128
rect 255681 290123 255747 290126
rect 90817 289914 90883 289917
rect 103830 289914 103836 289916
rect 90817 289912 103836 289914
rect 90817 289856 90822 289912
rect 90878 289856 103836 289912
rect 90817 289854 103836 289856
rect 90817 289851 90883 289854
rect 103830 289852 103836 289854
rect 103900 289852 103906 289916
rect 255405 289778 255471 289781
rect 253460 289776 255471 289778
rect 253460 289720 255410 289776
rect 255466 289720 255471 289776
rect 253460 289718 255471 289720
rect 255405 289715 255471 289718
rect 191741 289370 191807 289373
rect 254209 289370 254275 289373
rect 191741 289368 193660 289370
rect 191741 289312 191746 289368
rect 191802 289312 193660 289368
rect 191741 289310 193660 289312
rect 253460 289368 254275 289370
rect 253460 289312 254214 289368
rect 254270 289312 254275 289368
rect 253460 289310 254275 289312
rect 191741 289307 191807 289310
rect 254209 289307 254275 289310
rect 84101 289098 84167 289101
rect 103513 289098 103579 289101
rect 191649 289098 191715 289101
rect 84101 289096 191715 289098
rect 84101 289040 84106 289096
rect 84162 289040 103518 289096
rect 103574 289040 191654 289096
rect 191710 289040 191715 289096
rect 84101 289038 191715 289040
rect 84101 289035 84167 289038
rect 103513 289035 103579 289038
rect 191649 289035 191715 289038
rect 258574 289036 258580 289100
rect 258644 289098 258650 289100
rect 333973 289098 334039 289101
rect 258644 289096 334039 289098
rect 258644 289040 333978 289096
rect 334034 289040 334039 289096
rect 258644 289038 334039 289040
rect 258644 289036 258650 289038
rect 333973 289035 334039 289038
rect 255681 288826 255747 288829
rect 253460 288824 255747 288826
rect 253460 288768 255686 288824
rect 255742 288768 255747 288824
rect 253460 288766 255747 288768
rect 255681 288763 255747 288766
rect 89621 288554 89687 288557
rect 116577 288554 116643 288557
rect 89621 288552 116643 288554
rect 89621 288496 89626 288552
rect 89682 288496 116582 288552
rect 116638 288496 116643 288552
rect 89621 288494 116643 288496
rect 89621 288491 89687 288494
rect 116577 288491 116643 288494
rect 70158 288356 70164 288420
rect 70228 288418 70234 288420
rect 70393 288418 70459 288421
rect 255405 288418 255471 288421
rect 70228 288416 70459 288418
rect 70228 288360 70398 288416
rect 70454 288360 70459 288416
rect 253460 288416 255471 288418
rect 70228 288358 70459 288360
rect 70228 288356 70234 288358
rect 70393 288355 70459 288358
rect 72918 287676 72924 287740
rect 72988 287738 72994 287740
rect 73797 287738 73863 287741
rect 193630 287738 193690 288388
rect 253460 288360 255410 288416
rect 255466 288360 255471 288416
rect 253460 288358 255471 288360
rect 255405 288355 255471 288358
rect 259545 288010 259611 288013
rect 253460 288008 259611 288010
rect 253460 287952 259550 288008
rect 259606 287952 259611 288008
rect 253460 287950 259611 287952
rect 259545 287947 259611 287950
rect 72988 287736 73863 287738
rect 72988 287680 73802 287736
rect 73858 287680 73863 287736
rect 72988 287678 73863 287680
rect 72988 287676 72994 287678
rect 73797 287675 73863 287678
rect 180750 287678 193690 287738
rect 89161 287466 89227 287469
rect 89437 287466 89503 287469
rect 100569 287466 100635 287469
rect 89161 287464 100635 287466
rect 89161 287408 89166 287464
rect 89222 287408 89442 287464
rect 89498 287408 100574 287464
rect 100630 287408 100635 287464
rect 89161 287406 100635 287408
rect 89161 287403 89227 287406
rect 89437 287403 89503 287406
rect 100569 287403 100635 287406
rect 63125 287330 63191 287333
rect 80789 287330 80855 287333
rect 63125 287328 80855 287330
rect 63125 287272 63130 287328
rect 63186 287272 80794 287328
rect 80850 287272 80855 287328
rect 63125 287270 80855 287272
rect 63125 287267 63191 287270
rect 80789 287267 80855 287270
rect 85297 287330 85363 287333
rect 116025 287330 116091 287333
rect 85297 287328 116091 287330
rect 85297 287272 85302 287328
rect 85358 287272 116030 287328
rect 116086 287272 116091 287328
rect 85297 287270 116091 287272
rect 85297 287267 85363 287270
rect 116025 287267 116091 287270
rect 70158 287132 70164 287196
rect 70228 287194 70234 287196
rect 180750 287194 180810 287678
rect 190821 287466 190887 287469
rect 255681 287466 255747 287469
rect 190821 287464 193660 287466
rect 190821 287408 190826 287464
rect 190882 287408 193660 287464
rect 190821 287406 193660 287408
rect 253460 287464 255747 287466
rect 253460 287408 255686 287464
rect 255742 287408 255747 287464
rect 253460 287406 255747 287408
rect 190821 287403 190887 287406
rect 255681 287403 255747 287406
rect 70228 287134 180810 287194
rect 70228 287132 70234 287134
rect 71630 286996 71636 287060
rect 71700 287058 71706 287060
rect 192569 287058 192635 287061
rect 255589 287058 255655 287061
rect 71700 287056 192635 287058
rect 71700 287000 192574 287056
rect 192630 287000 192635 287056
rect 71700 286998 192635 287000
rect 253460 287056 255655 287058
rect 253460 287000 255594 287056
rect 255650 287000 255655 287056
rect 253460 286998 255655 287000
rect 71700 286996 71706 286998
rect 192569 286995 192635 286998
rect 255589 286995 255655 286998
rect 191741 286514 191807 286517
rect 255497 286514 255563 286517
rect 191741 286512 193660 286514
rect 191741 286456 191746 286512
rect 191802 286456 193660 286512
rect 191741 286454 193660 286456
rect 253460 286512 255563 286514
rect 253460 286456 255502 286512
rect 255558 286456 255563 286512
rect 253460 286454 255563 286456
rect 191741 286451 191807 286454
rect 255497 286451 255563 286454
rect 252829 286378 252895 286381
rect 252829 286376 252938 286378
rect 252829 286320 252834 286376
rect 252890 286320 252938 286376
rect 252829 286315 252938 286320
rect 252878 286076 252938 286315
rect 82629 285970 82695 285973
rect 114645 285970 114711 285973
rect 115841 285970 115907 285973
rect 82629 285968 115907 285970
rect 82629 285912 82634 285968
rect 82690 285912 114650 285968
rect 114706 285912 115846 285968
rect 115902 285912 115907 285968
rect 82629 285910 115907 285912
rect 82629 285907 82695 285910
rect 114645 285907 114711 285910
rect 115841 285907 115907 285910
rect 50705 285834 50771 285837
rect 74073 285834 74139 285837
rect 50705 285832 74139 285834
rect 50705 285776 50710 285832
rect 50766 285776 74078 285832
rect 74134 285776 74139 285832
rect 50705 285774 74139 285776
rect 50705 285771 50771 285774
rect 74073 285771 74139 285774
rect 95049 285698 95115 285701
rect 100017 285698 100083 285701
rect 256877 285698 256943 285701
rect 95049 285696 100083 285698
rect 95049 285640 95054 285696
rect 95110 285640 100022 285696
rect 100078 285640 100083 285696
rect 95049 285638 100083 285640
rect 253460 285696 256943 285698
rect 253460 285640 256882 285696
rect 256938 285640 256943 285696
rect 253460 285638 256943 285640
rect 95049 285635 95115 285638
rect 100017 285635 100083 285638
rect 256877 285635 256943 285638
rect 94129 285562 94195 285565
rect 94957 285562 95023 285565
rect 94129 285560 95023 285562
rect 94129 285504 94134 285560
rect 94190 285504 94962 285560
rect 95018 285504 95023 285560
rect 94129 285502 95023 285504
rect 94129 285499 94195 285502
rect 94957 285499 95023 285502
rect 96705 285562 96771 285565
rect 97717 285562 97783 285565
rect 96705 285560 97783 285562
rect 96705 285504 96710 285560
rect 96766 285504 97722 285560
rect 97778 285504 97783 285560
rect 96705 285502 97783 285504
rect 96705 285499 96771 285502
rect 97717 285499 97783 285502
rect 191649 285562 191715 285565
rect 191649 285560 193660 285562
rect 191649 285504 191654 285560
rect 191710 285504 193660 285560
rect 191649 285502 193660 285504
rect 191649 285499 191715 285502
rect 87505 285426 87571 285429
rect 97942 285426 97948 285428
rect 87505 285424 97948 285426
rect 87505 285368 87510 285424
rect 87566 285368 97948 285424
rect 87505 285366 97948 285368
rect 87505 285363 87571 285366
rect 97942 285364 97948 285366
rect 98012 285364 98018 285428
rect 583520 285276 584960 285516
rect 255405 285154 255471 285157
rect 253460 285152 255471 285154
rect 253460 285096 255410 285152
rect 255466 285096 255471 285152
rect 253460 285094 255471 285096
rect 255405 285091 255471 285094
rect 44081 284882 44147 284885
rect 61837 284882 61903 284885
rect 69013 284882 69079 284885
rect 185669 284882 185735 284885
rect 44081 284880 69079 284882
rect 44081 284824 44086 284880
rect 44142 284824 61842 284880
rect 61898 284824 69018 284880
rect 69074 284824 69079 284880
rect 44081 284822 69079 284824
rect 44081 284819 44147 284822
rect 61837 284819 61903 284822
rect 69013 284819 69079 284822
rect 122790 284880 185735 284882
rect 122790 284824 185674 284880
rect 185730 284824 185735 284880
rect 122790 284822 185735 284824
rect 94129 284474 94195 284477
rect 104934 284474 104940 284476
rect 94129 284472 104940 284474
rect 94129 284416 94134 284472
rect 94190 284416 104940 284472
rect 94129 284414 104940 284416
rect 94129 284411 94195 284414
rect 104934 284412 104940 284414
rect 105004 284412 105010 284476
rect 96705 284338 96771 284341
rect 122598 284338 122604 284340
rect 96705 284336 122604 284338
rect 96705 284280 96710 284336
rect 96766 284280 122604 284336
rect 96705 284278 122604 284280
rect 96705 284275 96771 284278
rect 122598 284276 122604 284278
rect 122668 284338 122674 284340
rect 122790 284338 122850 284822
rect 185669 284819 185735 284822
rect 260230 284820 260236 284884
rect 260300 284882 260306 284884
rect 342253 284882 342319 284885
rect 260300 284880 342319 284882
rect 260300 284824 342258 284880
rect 342314 284824 342319 284880
rect 260300 284822 342319 284824
rect 260300 284820 260306 284822
rect 342253 284819 342319 284822
rect 255405 284746 255471 284749
rect 253460 284744 255471 284746
rect 253460 284688 255410 284744
rect 255466 284688 255471 284744
rect 253460 284686 255471 284688
rect 255405 284683 255471 284686
rect 191741 284474 191807 284477
rect 191741 284472 193660 284474
rect 191741 284416 191746 284472
rect 191802 284416 193660 284472
rect 191741 284414 193660 284416
rect 191741 284411 191807 284414
rect 122668 284278 122850 284338
rect 190361 284338 190427 284341
rect 191649 284338 191715 284341
rect 254117 284338 254183 284341
rect 190361 284336 191715 284338
rect 190361 284280 190366 284336
rect 190422 284280 191654 284336
rect 191710 284280 191715 284336
rect 190361 284278 191715 284280
rect 253460 284336 254183 284338
rect 253460 284280 254122 284336
rect 254178 284280 254183 284336
rect 253460 284278 254183 284280
rect 122668 284276 122674 284278
rect 190361 284275 190427 284278
rect 191649 284275 191715 284278
rect 254117 284275 254183 284278
rect 74257 284204 74323 284205
rect 74206 284202 74212 284204
rect 74166 284142 74212 284202
rect 74276 284200 74323 284204
rect 74318 284144 74323 284200
rect 74206 284140 74212 284142
rect 74276 284140 74323 284144
rect 74257 284139 74323 284140
rect 107009 284202 107075 284205
rect 107561 284202 107627 284205
rect 116117 284202 116183 284205
rect 252921 284202 252987 284205
rect 107009 284200 116183 284202
rect 107009 284144 107014 284200
rect 107070 284144 107566 284200
rect 107622 284144 116122 284200
rect 116178 284144 116183 284200
rect 107009 284142 116183 284144
rect 107009 284139 107075 284142
rect 107561 284139 107627 284142
rect 116117 284139 116183 284142
rect 252878 284200 252987 284202
rect 252878 284144 252926 284200
rect 252982 284144 252987 284200
rect 252878 284139 252987 284144
rect 71175 283794 71241 283797
rect 71630 283794 71636 283796
rect 71175 283792 71636 283794
rect 71175 283736 71180 283792
rect 71236 283736 71636 283792
rect 71175 283734 71636 283736
rect 71175 283731 71241 283734
rect 71630 283732 71636 283734
rect 71700 283732 71706 283796
rect 252878 283764 252938 284139
rect 77385 283658 77451 283661
rect 60690 283656 77451 283658
rect 60690 283600 77390 283656
rect 77446 283600 77451 283656
rect 60690 283598 77451 283600
rect 60457 283522 60523 283525
rect 60690 283522 60750 283598
rect 77385 283595 77451 283598
rect 60457 283520 60750 283522
rect 60457 283464 60462 283520
rect 60518 283464 60750 283520
rect 60457 283462 60750 283464
rect 60457 283459 60523 283462
rect 71078 283460 71084 283524
rect 71148 283522 71154 283524
rect 71865 283522 71931 283525
rect 73521 283524 73587 283525
rect 71148 283520 71931 283522
rect 71148 283464 71870 283520
rect 71926 283464 71931 283520
rect 71148 283462 71931 283464
rect 71148 283460 71154 283462
rect 71865 283459 71931 283462
rect 73470 283460 73476 283524
rect 73540 283522 73587 283524
rect 73540 283520 73632 283522
rect 73582 283464 73632 283520
rect 73540 283462 73632 283464
rect 73540 283460 73587 283462
rect 95182 283460 95188 283524
rect 95252 283522 95258 283524
rect 95693 283522 95759 283525
rect 95252 283520 95759 283522
rect 95252 283464 95698 283520
rect 95754 283464 95759 283520
rect 95252 283462 95759 283464
rect 95252 283460 95258 283462
rect 73521 283459 73587 283460
rect 95693 283459 95759 283462
rect 96654 283460 96660 283524
rect 96724 283522 96730 283524
rect 96797 283522 96863 283525
rect 96724 283520 96863 283522
rect 96724 283464 96802 283520
rect 96858 283464 96863 283520
rect 96724 283462 96863 283464
rect 96724 283460 96730 283462
rect 96797 283459 96863 283462
rect 100569 283522 100635 283525
rect 114553 283522 114619 283525
rect 100569 283520 114619 283522
rect 100569 283464 100574 283520
rect 100630 283464 114558 283520
rect 114614 283464 114619 283520
rect 100569 283462 114619 283464
rect 100569 283459 100635 283462
rect 114553 283459 114619 283462
rect 191741 283522 191807 283525
rect 191741 283520 193660 283522
rect 191741 283464 191746 283520
rect 191802 283464 193660 283520
rect 191741 283462 193660 283464
rect 191741 283459 191807 283462
rect 260046 283460 260052 283524
rect 260116 283522 260122 283524
rect 339493 283522 339559 283525
rect 260116 283520 339559 283522
rect 260116 283464 339498 283520
rect 339554 283464 339559 283520
rect 260116 283462 339559 283464
rect 260116 283460 260122 283462
rect 339493 283459 339559 283462
rect 255405 283386 255471 283389
rect 253460 283384 255471 283386
rect 253460 283328 255410 283384
rect 255466 283328 255471 283384
rect 253460 283326 255471 283328
rect 255405 283323 255471 283326
rect 65926 283188 65932 283252
rect 65996 283250 66002 283252
rect 71037 283250 71103 283253
rect 65996 283248 71103 283250
rect 65996 283192 71042 283248
rect 71098 283192 71103 283248
rect 65996 283190 71103 283192
rect 65996 283188 66002 283190
rect 71037 283187 71103 283190
rect 69062 282437 69122 282948
rect 117998 282916 118004 282980
rect 118068 282978 118074 282980
rect 120165 282978 120231 282981
rect 118068 282976 120231 282978
rect 118068 282920 120170 282976
rect 120226 282920 120231 282976
rect 118068 282918 120231 282920
rect 118068 282916 118074 282918
rect 120165 282915 120231 282918
rect 191281 282842 191347 282845
rect 255405 282842 255471 282845
rect 103470 282840 191347 282842
rect 103470 282784 191286 282840
rect 191342 282784 191347 282840
rect 103470 282782 191347 282784
rect 253460 282840 255471 282842
rect 253460 282784 255410 282840
rect 255466 282784 255471 282840
rect 253460 282782 255471 282784
rect 99966 282706 99972 282708
rect 98716 282646 99972 282706
rect 99966 282644 99972 282646
rect 100036 282706 100042 282708
rect 101990 282706 101996 282708
rect 100036 282646 101996 282706
rect 100036 282644 100042 282646
rect 101990 282644 101996 282646
rect 102060 282706 102066 282708
rect 103470 282706 103530 282782
rect 191281 282779 191347 282782
rect 255405 282779 255471 282782
rect 102060 282646 103530 282706
rect 102060 282644 102066 282646
rect 192477 282570 192543 282573
rect 192477 282568 193660 282570
rect 192477 282512 192482 282568
rect 192538 282512 193660 282568
rect 192477 282510 193660 282512
rect 192477 282507 192543 282510
rect 69013 282432 69122 282437
rect 100661 282434 100727 282437
rect 69013 282376 69018 282432
rect 69074 282376 69122 282432
rect 69013 282374 69122 282376
rect 98686 282432 100727 282434
rect 98686 282376 100666 282432
rect 100722 282376 100727 282432
rect 98686 282374 100727 282376
rect 69013 282371 69079 282374
rect 53557 282162 53623 282165
rect 62982 282162 62988 282164
rect 53557 282160 62988 282162
rect 53557 282104 53562 282160
rect 53618 282104 62988 282160
rect 53557 282102 62988 282104
rect 53557 282099 53623 282102
rect 62982 282100 62988 282102
rect 63052 282162 63058 282164
rect 63052 282102 68908 282162
rect 63052 282100 63058 282102
rect 98686 281860 98746 282374
rect 100661 282371 100727 282374
rect 253430 282298 253490 282404
rect 263593 282298 263659 282301
rect 253430 282296 263659 282298
rect 253430 282240 263598 282296
rect 263654 282240 263659 282296
rect 253430 282238 263659 282240
rect 263593 282235 263659 282238
rect 255497 282026 255563 282029
rect 253460 282024 255563 282026
rect 253460 281968 255502 282024
rect 255558 281968 255563 282024
rect 253460 281966 255563 281968
rect 255497 281963 255563 281966
rect 191465 281618 191531 281621
rect 191465 281616 193660 281618
rect 191465 281560 191470 281616
rect 191526 281560 193660 281616
rect 191465 281558 193660 281560
rect 191465 281555 191531 281558
rect 252878 281349 252938 281452
rect 67541 281346 67607 281349
rect 67541 281344 68908 281346
rect 67541 281288 67546 281344
rect 67602 281288 68908 281344
rect 67541 281286 68908 281288
rect 252829 281344 252938 281349
rect 252829 281288 252834 281344
rect 252890 281288 252938 281344
rect 252829 281286 252938 281288
rect 67541 281283 67607 281286
rect 252829 281283 252895 281286
rect 100753 281074 100819 281077
rect 255497 281074 255563 281077
rect 98716 281072 100819 281074
rect 98716 281016 100758 281072
rect 100814 281016 100819 281072
rect 98716 281014 100819 281016
rect 253460 281072 255563 281074
rect 253460 281016 255502 281072
rect 255558 281016 255563 281072
rect 253460 281014 255563 281016
rect 100753 281011 100819 281014
rect 255497 281011 255563 281014
rect 191557 280666 191623 280669
rect 255405 280666 255471 280669
rect 191557 280664 193660 280666
rect 191557 280608 191562 280664
rect 191618 280608 193660 280664
rect 191557 280606 193660 280608
rect 253460 280664 255471 280666
rect 253460 280608 255410 280664
rect 255466 280608 255471 280664
rect 253460 280606 255471 280608
rect 191557 280603 191623 280606
rect 255405 280603 255471 280606
rect 67950 280468 67956 280532
rect 68020 280530 68026 280532
rect 68020 280470 68908 280530
rect 68020 280468 68026 280470
rect 99373 280258 99439 280261
rect 101489 280258 101555 280261
rect 98716 280256 101555 280258
rect -960 279972 480 280212
rect 98716 280200 99378 280256
rect 99434 280200 101494 280256
rect 101550 280200 101555 280256
rect 98716 280198 101555 280200
rect 99373 280195 99439 280198
rect 101489 280195 101555 280198
rect 255405 280122 255471 280125
rect 253460 280120 255471 280122
rect 253460 280064 255410 280120
rect 255466 280064 255471 280120
rect 253460 280062 255471 280064
rect 255405 280059 255471 280062
rect 66621 279714 66687 279717
rect 191741 279714 191807 279717
rect 255589 279714 255655 279717
rect 66621 279712 68908 279714
rect 66621 279656 66626 279712
rect 66682 279656 68908 279712
rect 66621 279654 68908 279656
rect 191741 279712 193660 279714
rect 191741 279656 191746 279712
rect 191802 279656 193660 279712
rect 191741 279654 193660 279656
rect 253460 279712 255655 279714
rect 253460 279656 255594 279712
rect 255650 279656 255655 279712
rect 253460 279654 255655 279656
rect 66621 279651 66687 279654
rect 191741 279651 191807 279654
rect 255589 279651 255655 279654
rect 101581 279442 101647 279445
rect 98716 279440 101647 279442
rect 98716 279384 101586 279440
rect 101642 279384 101647 279440
rect 98716 279382 101647 279384
rect 101581 279379 101647 279382
rect 255814 279380 255820 279444
rect 255884 279442 255890 279444
rect 583017 279442 583083 279445
rect 255884 279440 583083 279442
rect 255884 279384 583022 279440
rect 583078 279384 583083 279440
rect 255884 279382 583083 279384
rect 255884 279380 255890 279382
rect 583017 279379 583083 279382
rect 255313 279306 255379 279309
rect 253460 279304 255379 279306
rect 253460 279248 255318 279304
rect 255374 279248 255379 279304
rect 253460 279246 255379 279248
rect 255313 279243 255379 279246
rect 66805 278898 66871 278901
rect 66805 278896 68908 278898
rect 66805 278840 66810 278896
rect 66866 278840 68908 278896
rect 66805 278838 68908 278840
rect 66805 278835 66871 278838
rect 100753 278762 100819 278765
rect 135253 278762 135319 278765
rect 100753 278760 135319 278762
rect 100753 278704 100758 278760
rect 100814 278704 135258 278760
rect 135314 278704 135319 278760
rect 100753 278702 135319 278704
rect 100753 278699 100819 278702
rect 135253 278699 135319 278702
rect 191649 278762 191715 278765
rect 255313 278762 255379 278765
rect 191649 278760 193660 278762
rect 191649 278704 191654 278760
rect 191710 278704 193660 278760
rect 191649 278702 193660 278704
rect 253460 278760 255379 278762
rect 253460 278704 255318 278760
rect 255374 278704 255379 278760
rect 253460 278702 255379 278704
rect 191649 278699 191715 278702
rect 255313 278699 255379 278702
rect 101949 278626 102015 278629
rect 98716 278624 102015 278626
rect 98716 278568 101954 278624
rect 102010 278568 102015 278624
rect 98716 278566 102015 278568
rect 101949 278563 102015 278566
rect 255405 278354 255471 278357
rect 253460 278352 255471 278354
rect 253460 278296 255410 278352
rect 255466 278296 255471 278352
rect 253460 278294 255471 278296
rect 255405 278291 255471 278294
rect 66805 278082 66871 278085
rect 256601 278082 256667 278085
rect 272057 278082 272123 278085
rect 66805 278080 68908 278082
rect 66805 278024 66810 278080
rect 66866 278024 68908 278080
rect 66805 278022 68908 278024
rect 256601 278080 272123 278082
rect 256601 278024 256606 278080
rect 256662 278024 272062 278080
rect 272118 278024 272123 278080
rect 256601 278022 272123 278024
rect 66805 278019 66871 278022
rect 256601 278019 256667 278022
rect 272057 278019 272123 278022
rect 102041 277810 102107 277813
rect 98716 277808 102107 277810
rect 98716 277752 102046 277808
rect 102102 277752 102107 277808
rect 98716 277750 102107 277752
rect 102041 277747 102107 277750
rect 191741 277810 191807 277813
rect 255405 277810 255471 277813
rect 191741 277808 193660 277810
rect 191741 277752 191746 277808
rect 191802 277752 193660 277808
rect 191741 277750 193660 277752
rect 253460 277808 255471 277810
rect 253460 277752 255410 277808
rect 255466 277752 255471 277808
rect 253460 277750 255471 277752
rect 191741 277747 191807 277750
rect 255405 277747 255471 277750
rect 68277 277402 68343 277405
rect 255497 277402 255563 277405
rect 68277 277400 68938 277402
rect 68277 277344 68282 277400
rect 68338 277344 68938 277400
rect 68277 277342 68938 277344
rect 253460 277400 255563 277402
rect 253460 277344 255502 277400
rect 255558 277344 255563 277400
rect 253460 277342 255563 277344
rect 68277 277339 68343 277342
rect 68878 277236 68938 277342
rect 255497 277339 255563 277342
rect 255313 276994 255379 276997
rect 253460 276992 255379 276994
rect 66805 276450 66871 276453
rect 98686 276450 98746 276964
rect 253460 276936 255318 276992
rect 255374 276936 255379 276992
rect 253460 276934 255379 276936
rect 255313 276931 255379 276934
rect 191097 276858 191163 276861
rect 193213 276858 193279 276861
rect 191097 276856 193660 276858
rect 191097 276800 191102 276856
rect 191158 276800 193218 276856
rect 193274 276800 193660 276856
rect 191097 276798 193660 276800
rect 191097 276795 191163 276798
rect 193213 276795 193279 276798
rect 156597 276722 156663 276725
rect 193254 276722 193260 276724
rect 156597 276720 193260 276722
rect 156597 276664 156602 276720
rect 156658 276664 193260 276720
rect 156597 276662 193260 276664
rect 156597 276659 156663 276662
rect 193254 276660 193260 276662
rect 193324 276660 193330 276724
rect 256601 276450 256667 276453
rect 66805 276448 68908 276450
rect 66805 276392 66810 276448
rect 66866 276392 68908 276448
rect 66805 276390 68908 276392
rect 98686 276390 103530 276450
rect 253460 276448 256667 276450
rect 253460 276392 256606 276448
rect 256662 276392 256667 276448
rect 253460 276390 256667 276392
rect 66805 276387 66871 276390
rect 52310 276116 52316 276180
rect 52380 276178 52386 276180
rect 52453 276178 52519 276181
rect 102041 276178 102107 276181
rect 52380 276176 52519 276178
rect 52380 276120 52458 276176
rect 52514 276120 52519 276176
rect 52380 276118 52519 276120
rect 98716 276176 102107 276178
rect 98716 276120 102046 276176
rect 102102 276120 102107 276176
rect 98716 276118 102107 276120
rect 52380 276116 52386 276118
rect 52453 276115 52519 276118
rect 102041 276115 102107 276118
rect 103470 276042 103530 276390
rect 256601 276387 256667 276390
rect 118785 276042 118851 276045
rect 257061 276042 257127 276045
rect 103470 276040 118851 276042
rect 103470 275984 118790 276040
rect 118846 275984 118851 276040
rect 103470 275982 118851 275984
rect 253460 276040 257127 276042
rect 253460 275984 257066 276040
rect 257122 275984 257127 276040
rect 253460 275982 257127 275984
rect 118785 275979 118851 275982
rect 257061 275979 257127 275982
rect 257337 276042 257403 276045
rect 258073 276042 258139 276045
rect 257337 276040 258139 276042
rect 257337 275984 257342 276040
rect 257398 275984 258078 276040
rect 258134 275984 258139 276040
rect 257337 275982 258139 275984
rect 257337 275979 257403 275982
rect 258073 275979 258139 275982
rect 57513 275906 57579 275909
rect 67766 275906 67772 275908
rect 57513 275904 67772 275906
rect 57513 275848 57518 275904
rect 57574 275848 67772 275904
rect 57513 275846 67772 275848
rect 57513 275843 57579 275846
rect 67766 275844 67772 275846
rect 67836 275844 67842 275908
rect 101949 275906 102015 275909
rect 121545 275906 121611 275909
rect 101949 275904 121611 275906
rect 101949 275848 101954 275904
rect 102010 275848 121550 275904
rect 121606 275848 121611 275904
rect 101949 275846 121611 275848
rect 101949 275843 102015 275846
rect 121545 275843 121611 275846
rect 191649 275770 191715 275773
rect 191649 275768 193660 275770
rect 191649 275712 191654 275768
rect 191710 275712 193660 275768
rect 191649 275710 193660 275712
rect 191649 275707 191715 275710
rect 66897 275634 66963 275637
rect 255405 275634 255471 275637
rect 66897 275632 68908 275634
rect 66897 275576 66902 275632
rect 66958 275576 68908 275632
rect 66897 275574 68908 275576
rect 253460 275632 255471 275634
rect 253460 275576 255410 275632
rect 255466 275576 255471 275632
rect 253460 275574 255471 275576
rect 66897 275571 66963 275574
rect 255405 275571 255471 275574
rect 100753 275362 100819 275365
rect 98716 275360 100819 275362
rect 98716 275304 100758 275360
rect 100814 275304 100819 275360
rect 98716 275302 100819 275304
rect 100753 275299 100819 275302
rect 32949 275226 33015 275229
rect 57513 275226 57579 275229
rect 32949 275224 57579 275226
rect 32949 275168 32954 275224
rect 33010 275168 57518 275224
rect 57574 275168 57579 275224
rect 32949 275166 57579 275168
rect 32949 275163 33015 275166
rect 57513 275163 57579 275166
rect 255589 275090 255655 275093
rect 253460 275088 255655 275090
rect 253460 275032 255594 275088
rect 255650 275032 255655 275088
rect 253460 275030 255655 275032
rect 255589 275027 255655 275030
rect 67766 274756 67772 274820
rect 67836 274818 67842 274820
rect 191741 274818 191807 274821
rect 67836 274758 68908 274818
rect 191741 274816 193660 274818
rect 191741 274760 191746 274816
rect 191802 274760 193660 274816
rect 191741 274758 193660 274760
rect 67836 274756 67842 274758
rect 191741 274755 191807 274758
rect 118785 274684 118851 274685
rect 118734 274620 118740 274684
rect 118804 274682 118851 274684
rect 121545 274682 121611 274685
rect 121678 274682 121684 274684
rect 118804 274680 118896 274682
rect 118846 274624 118896 274680
rect 118804 274622 118896 274624
rect 121545 274680 121684 274682
rect 121545 274624 121550 274680
rect 121606 274624 121684 274680
rect 121545 274622 121684 274624
rect 118804 274620 118851 274622
rect 118785 274619 118851 274620
rect 121545 274619 121611 274622
rect 121678 274620 121684 274622
rect 121748 274620 121754 274684
rect 256601 274682 256667 274685
rect 253460 274680 256667 274682
rect 253460 274624 256606 274680
rect 256662 274624 256667 274680
rect 253460 274622 256667 274624
rect 256601 274619 256667 274622
rect 100845 274546 100911 274549
rect 98716 274544 100911 274546
rect 98716 274488 100850 274544
rect 100906 274488 100911 274544
rect 98716 274486 100911 274488
rect 100845 274483 100911 274486
rect 255405 274274 255471 274277
rect 253460 274272 255471 274274
rect 253460 274216 255410 274272
rect 255466 274216 255471 274272
rect 253460 274214 255471 274216
rect 255405 274211 255471 274214
rect 66529 274002 66595 274005
rect 66529 274000 68908 274002
rect 66529 273944 66534 274000
rect 66590 273944 68908 274000
rect 66529 273942 68908 273944
rect 66529 273939 66595 273942
rect 193121 273866 193187 273869
rect 193121 273864 193660 273866
rect 193121 273808 193126 273864
rect 193182 273808 193660 273864
rect 193121 273806 193660 273808
rect 193121 273803 193187 273806
rect 100753 273730 100819 273733
rect 254025 273730 254091 273733
rect 98716 273728 100819 273730
rect 98716 273672 100758 273728
rect 100814 273672 100819 273728
rect 98716 273670 100819 273672
rect 253460 273728 254091 273730
rect 253460 273672 254030 273728
rect 254086 273672 254091 273728
rect 253460 273670 254091 273672
rect 100753 273667 100819 273670
rect 254025 273667 254091 273670
rect 60549 273322 60615 273325
rect 99189 273322 99255 273325
rect 102317 273322 102383 273325
rect 253933 273322 253999 273325
rect 60549 273320 62866 273322
rect 60549 273264 60554 273320
rect 60610 273264 62866 273320
rect 60549 273262 62866 273264
rect 60549 273259 60615 273262
rect 62806 273189 62866 273262
rect 99189 273320 102383 273322
rect 99189 273264 99194 273320
rect 99250 273264 102322 273320
rect 102378 273264 102383 273320
rect 99189 273262 102383 273264
rect 253460 273320 253999 273322
rect 253460 273264 253938 273320
rect 253994 273264 253999 273320
rect 253460 273262 253999 273264
rect 99189 273259 99255 273262
rect 102317 273259 102383 273262
rect 253933 273259 253999 273262
rect 62806 273184 62915 273189
rect 62806 273128 62854 273184
rect 62910 273128 62915 273184
rect 62806 273126 62915 273128
rect 62849 273123 62915 273126
rect 66253 273186 66319 273189
rect 109677 273186 109743 273189
rect 66253 273184 68908 273186
rect 66253 273128 66258 273184
rect 66314 273128 68908 273184
rect 66253 273126 68908 273128
rect 98686 273184 109743 273186
rect 98686 273128 109682 273184
rect 109738 273128 109743 273184
rect 98686 273126 109743 273128
rect 66253 273123 66319 273126
rect 98686 272884 98746 273126
rect 109677 273123 109743 273126
rect 191741 272914 191807 272917
rect 191741 272912 193660 272914
rect 191741 272856 191746 272912
rect 191802 272856 193660 272912
rect 191741 272854 193660 272856
rect 191741 272851 191807 272854
rect 253933 272778 253999 272781
rect 253460 272776 253999 272778
rect 253460 272720 253938 272776
rect 253994 272720 253999 272776
rect 253460 272718 253999 272720
rect 253933 272715 253999 272718
rect 256693 272506 256759 272509
rect 266353 272506 266419 272509
rect 256693 272504 266419 272506
rect 256693 272448 256698 272504
rect 256754 272448 266358 272504
rect 266414 272448 266419 272504
rect 256693 272446 266419 272448
rect 256693 272443 256759 272446
rect 266353 272443 266419 272446
rect 66805 272370 66871 272373
rect 255497 272370 255563 272373
rect 66805 272368 68908 272370
rect 66805 272312 66810 272368
rect 66866 272312 68908 272368
rect 66805 272310 68908 272312
rect 253460 272368 255563 272370
rect 253460 272312 255502 272368
rect 255558 272312 255563 272368
rect 253460 272310 255563 272312
rect 66805 272307 66871 272310
rect 255497 272307 255563 272310
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 99189 272098 99255 272101
rect 101397 272098 101463 272101
rect 98716 272096 101463 272098
rect 98716 272040 99194 272096
rect 99250 272040 101402 272096
rect 101458 272040 101463 272096
rect 583520 272084 584960 272174
rect 98716 272038 101463 272040
rect 99189 272035 99255 272038
rect 101397 272035 101463 272038
rect 53465 271962 53531 271965
rect 66253 271962 66319 271965
rect 53465 271960 66319 271962
rect 53465 271904 53470 271960
rect 53526 271904 66258 271960
rect 66314 271904 66319 271960
rect 53465 271902 66319 271904
rect 53465 271899 53531 271902
rect 66253 271899 66319 271902
rect 112253 271964 112319 271965
rect 112253 271960 112300 271964
rect 112364 271962 112370 271964
rect 112253 271904 112258 271960
rect 112253 271900 112300 271904
rect 112364 271902 112410 271962
rect 112364 271900 112370 271902
rect 115974 271900 115980 271964
rect 116044 271962 116050 271964
rect 116853 271962 116919 271965
rect 116044 271960 116919 271962
rect 116044 271904 116858 271960
rect 116914 271904 116919 271960
rect 116044 271902 116919 271904
rect 116044 271900 116050 271902
rect 112253 271899 112319 271900
rect 116853 271899 116919 271902
rect 191189 271962 191255 271965
rect 255405 271962 255471 271965
rect 191189 271960 193660 271962
rect 191189 271904 191194 271960
rect 191250 271904 193660 271960
rect 191189 271902 193660 271904
rect 253460 271960 255471 271962
rect 253460 271904 255410 271960
rect 255466 271904 255471 271960
rect 253460 271902 255471 271904
rect 191189 271899 191255 271902
rect 255405 271899 255471 271902
rect 66161 271554 66227 271557
rect 66161 271552 68908 271554
rect 66161 271496 66166 271552
rect 66222 271496 68908 271552
rect 66161 271494 68908 271496
rect 66161 271491 66227 271494
rect 255497 271418 255563 271421
rect 253460 271416 255563 271418
rect 253460 271360 255502 271416
rect 255558 271360 255563 271416
rect 253460 271358 255563 271360
rect 255497 271355 255563 271358
rect 101673 271282 101739 271285
rect 98716 271280 101739 271282
rect 98716 271224 101678 271280
rect 101734 271224 101739 271280
rect 98716 271222 101739 271224
rect 101673 271219 101739 271222
rect 98494 271084 98500 271148
rect 98564 271146 98570 271148
rect 104341 271146 104407 271149
rect 98564 271144 104407 271146
rect 98564 271088 104346 271144
rect 104402 271088 104407 271144
rect 98564 271086 104407 271088
rect 98564 271084 98570 271086
rect 104341 271083 104407 271086
rect 255814 271084 255820 271148
rect 255884 271146 255890 271148
rect 583569 271146 583635 271149
rect 255884 271144 583635 271146
rect 255884 271088 583574 271144
rect 583630 271088 583635 271144
rect 255884 271086 583635 271088
rect 255884 271084 255890 271086
rect 583569 271083 583635 271086
rect 191097 271010 191163 271013
rect 255313 271010 255379 271013
rect 191097 271008 193660 271010
rect 191097 270952 191102 271008
rect 191158 270952 193660 271008
rect 191097 270950 193660 270952
rect 253460 271008 255379 271010
rect 253460 270952 255318 271008
rect 255374 270952 255379 271008
rect 253460 270950 255379 270952
rect 191097 270947 191163 270950
rect 255313 270947 255379 270950
rect 61745 270738 61811 270741
rect 66161 270738 66227 270741
rect 61745 270736 66227 270738
rect 61745 270680 61750 270736
rect 61806 270680 66166 270736
rect 66222 270680 66227 270736
rect 61745 270678 66227 270680
rect 61745 270675 61811 270678
rect 66161 270675 66227 270678
rect 66805 270738 66871 270741
rect 66805 270736 68908 270738
rect 66805 270680 66810 270736
rect 66866 270680 68908 270736
rect 66805 270678 68908 270680
rect 66805 270675 66871 270678
rect 259637 270602 259703 270605
rect 253460 270600 259703 270602
rect 253460 270544 259642 270600
rect 259698 270544 259703 270600
rect 253460 270542 259703 270544
rect 259637 270539 259703 270542
rect 103973 270466 104039 270469
rect 98716 270464 104039 270466
rect 98716 270408 103978 270464
rect 104034 270408 104039 270464
rect 98716 270406 104039 270408
rect 103973 270403 104039 270406
rect 105629 270466 105695 270469
rect 111742 270466 111748 270468
rect 105629 270464 111748 270466
rect 105629 270408 105634 270464
rect 105690 270408 111748 270464
rect 105629 270406 111748 270408
rect 105629 270403 105695 270406
rect 111742 270404 111748 270406
rect 111812 270404 111818 270468
rect 191741 270058 191807 270061
rect 255405 270058 255471 270061
rect 191741 270056 193660 270058
rect 191741 270000 191746 270056
rect 191802 270000 193660 270056
rect 191741 269998 193660 270000
rect 253460 270056 255471 270058
rect 253460 270000 255410 270056
rect 255466 270000 255471 270056
rect 253460 269998 255471 270000
rect 191741 269995 191807 269998
rect 255405 269995 255471 269998
rect 68878 269378 68938 269892
rect 256509 269786 256575 269789
rect 266445 269786 266511 269789
rect 256509 269784 266511 269786
rect 256509 269728 256514 269784
rect 256570 269728 266450 269784
rect 266506 269728 266511 269784
rect 256509 269726 266511 269728
rect 256509 269723 256575 269726
rect 266445 269723 266511 269726
rect 100753 269650 100819 269653
rect 98716 269648 100819 269650
rect 98716 269592 100758 269648
rect 100814 269592 100819 269648
rect 98716 269590 100819 269592
rect 100753 269587 100819 269590
rect 64830 269318 68938 269378
rect 252878 269381 252938 269620
rect 252878 269376 252987 269381
rect 252878 269320 252926 269376
rect 252982 269320 252987 269376
rect 252878 269318 252987 269320
rect 60549 269242 60615 269245
rect 61878 269242 61884 269244
rect 60549 269240 61884 269242
rect 60549 269184 60554 269240
rect 60610 269184 61884 269240
rect 60549 269182 61884 269184
rect 60549 269179 60615 269182
rect 61878 269180 61884 269182
rect 61948 269242 61954 269244
rect 64830 269242 64890 269318
rect 252921 269315 252987 269318
rect 106825 269244 106891 269245
rect 106774 269242 106780 269244
rect 61948 269182 64890 269242
rect 106734 269182 106780 269242
rect 106844 269240 106891 269244
rect 106886 269184 106891 269240
rect 61948 269180 61954 269182
rect 106774 269180 106780 269182
rect 106844 269180 106891 269184
rect 106825 269179 106891 269180
rect 191649 269106 191715 269109
rect 255497 269106 255563 269109
rect 191649 269104 193660 269106
rect 68878 268562 68938 269076
rect 191649 269048 191654 269104
rect 191710 269048 193660 269104
rect 191649 269046 193660 269048
rect 253460 269104 255563 269106
rect 253460 269048 255502 269104
rect 255558 269048 255563 269104
rect 253460 269046 255563 269048
rect 191649 269043 191715 269046
rect 255497 269043 255563 269046
rect 100845 268834 100911 268837
rect 98716 268832 100911 268834
rect 98716 268776 100850 268832
rect 100906 268776 100911 268832
rect 98716 268774 100911 268776
rect 100845 268771 100911 268774
rect 256601 268698 256667 268701
rect 253460 268696 256667 268698
rect 253460 268640 256606 268696
rect 256662 268640 256667 268696
rect 253460 268638 256667 268640
rect 256601 268635 256667 268638
rect 64830 268502 68938 268562
rect 64830 268018 64890 268502
rect 269757 268426 269823 268429
rect 253430 268424 269823 268426
rect 253430 268368 269762 268424
rect 269818 268368 269823 268424
rect 253430 268366 269823 268368
rect 66161 268290 66227 268293
rect 66161 268288 68908 268290
rect 66161 268232 66166 268288
rect 66222 268232 68908 268288
rect 253430 268260 253490 268366
rect 269757 268363 269823 268366
rect 66161 268230 68908 268232
rect 66161 268227 66227 268230
rect 100753 268018 100819 268021
rect 45510 267958 64890 268018
rect 98716 268016 100819 268018
rect 98716 267960 100758 268016
rect 100814 267960 100819 268016
rect 98716 267958 100819 267960
rect 45510 267885 45570 267958
rect 100753 267955 100819 267958
rect 41045 267882 41111 267885
rect 45461 267882 45570 267885
rect 41045 267880 45570 267882
rect 41045 267824 41050 267880
rect 41106 267824 45466 267880
rect 45522 267824 45570 267880
rect 41045 267822 45570 267824
rect 188521 267882 188587 267885
rect 193630 267882 193690 268124
rect 188521 267880 193690 267882
rect 188521 267824 188526 267880
rect 188582 267824 193690 267880
rect 188521 267822 193690 267824
rect 41045 267819 41111 267822
rect 45461 267819 45527 267822
rect 188521 267819 188587 267822
rect 252878 267613 252938 267716
rect 252829 267608 252938 267613
rect 252829 267552 252834 267608
rect 252890 267552 252938 267608
rect 252829 267550 252938 267552
rect 252829 267547 252895 267550
rect 66805 267474 66871 267477
rect 66805 267472 68908 267474
rect 66805 267416 66810 267472
rect 66866 267416 68908 267472
rect 66805 267414 68908 267416
rect 66805 267411 66871 267414
rect -960 267202 480 267292
rect 100150 267276 100156 267340
rect 100220 267338 100226 267340
rect 110638 267338 110644 267340
rect 100220 267278 110644 267338
rect 100220 267276 100226 267278
rect 110638 267276 110644 267278
rect 110708 267276 110714 267340
rect 255405 267338 255471 267341
rect 253460 267336 255471 267338
rect 253460 267280 255410 267336
rect 255466 267280 255471 267336
rect 253460 267278 255471 267280
rect 255405 267275 255471 267278
rect 3049 267202 3115 267205
rect 101397 267202 101463 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect 98716 267200 101463 267202
rect 98716 267144 101402 267200
rect 101458 267144 101463 267200
rect 98716 267142 101463 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 101397 267139 101463 267142
rect 98729 267066 98795 267069
rect 109534 267066 109540 267068
rect 98729 267064 109540 267066
rect 98729 267008 98734 267064
rect 98790 267008 109540 267064
rect 98729 267006 109540 267008
rect 98729 267003 98795 267006
rect 109534 267004 109540 267006
rect 109604 267004 109610 267068
rect 191465 267066 191531 267069
rect 273437 267066 273503 267069
rect 582557 267066 582623 267069
rect 191465 267064 193660 267066
rect 191465 267008 191470 267064
rect 191526 267008 193660 267064
rect 191465 267006 193660 267008
rect 273437 267064 582623 267066
rect 273437 267008 273442 267064
rect 273498 267008 582562 267064
rect 582618 267008 582623 267064
rect 273437 267006 582623 267008
rect 191465 267003 191531 267006
rect 273437 267003 273503 267006
rect 582557 267003 582623 267006
rect 255405 266930 255471 266933
rect 253460 266928 255471 266930
rect 253460 266872 255410 266928
rect 255466 266872 255471 266928
rect 253460 266870 255471 266872
rect 255405 266867 255471 266870
rect 64638 266460 64644 266524
rect 64708 266522 64714 266524
rect 66253 266522 66319 266525
rect 68878 266522 68938 266628
rect 64708 266520 68938 266522
rect 64708 266464 66258 266520
rect 66314 266464 68938 266520
rect 64708 266462 68938 266464
rect 255497 266522 255563 266525
rect 262213 266522 262279 266525
rect 263358 266522 263364 266524
rect 255497 266520 258090 266522
rect 255497 266464 255502 266520
rect 255558 266464 258090 266520
rect 255497 266462 258090 266464
rect 64708 266460 64714 266462
rect 66253 266459 66319 266462
rect 255497 266459 255563 266462
rect 99230 266386 99236 266388
rect 98716 266326 99236 266386
rect 99230 266324 99236 266326
rect 99300 266324 99306 266388
rect 256509 266386 256575 266389
rect 253460 266384 256575 266386
rect 253460 266328 256514 266384
rect 256570 266328 256575 266384
rect 253460 266326 256575 266328
rect 258030 266386 258090 266462
rect 262213 266520 263364 266522
rect 262213 266464 262218 266520
rect 262274 266464 263364 266520
rect 262213 266462 263364 266464
rect 262213 266459 262279 266462
rect 263358 266460 263364 266462
rect 263428 266522 263434 266524
rect 263726 266522 263732 266524
rect 263428 266462 263732 266522
rect 263428 266460 263434 266462
rect 263726 266460 263732 266462
rect 263796 266460 263802 266524
rect 273437 266386 273503 266389
rect 258030 266384 273503 266386
rect 258030 266328 273442 266384
rect 273498 266328 273503 266384
rect 258030 266326 273503 266328
rect 256509 266323 256575 266326
rect 273437 266323 273503 266326
rect 191741 266114 191807 266117
rect 191741 266112 193660 266114
rect 191741 266056 191746 266112
rect 191802 266056 193660 266112
rect 191741 266054 193660 266056
rect 191741 266051 191807 266054
rect 253974 265978 253980 265980
rect 253460 265918 253980 265978
rect 253974 265916 253980 265918
rect 254044 265978 254050 265980
rect 254044 265918 258090 265978
rect 254044 265916 254050 265918
rect 68878 265298 68938 265812
rect 100017 265570 100083 265573
rect 255313 265570 255379 265573
rect 98716 265568 100083 265570
rect 98716 265512 100022 265568
rect 100078 265512 100083 265568
rect 98716 265510 100083 265512
rect 253460 265568 255379 265570
rect 253460 265512 255318 265568
rect 255374 265512 255379 265568
rect 253460 265510 255379 265512
rect 258030 265570 258090 265918
rect 271137 265570 271203 265573
rect 258030 265568 271203 265570
rect 258030 265512 271142 265568
rect 271198 265512 271203 265568
rect 258030 265510 271203 265512
rect 100017 265507 100083 265510
rect 255313 265507 255379 265510
rect 271137 265507 271203 265510
rect 64830 265238 68938 265298
rect 48221 265026 48287 265029
rect 64830 265026 64890 265238
rect 191281 265162 191347 265165
rect 191281 265160 193660 265162
rect 191281 265104 191286 265160
rect 191342 265104 193660 265160
rect 191281 265102 193660 265104
rect 191281 265099 191347 265102
rect 48221 265024 64890 265026
rect 48221 264968 48226 265024
rect 48282 264968 64890 265024
rect 48221 264966 64890 264968
rect 66805 265026 66871 265029
rect 254158 265026 254164 265028
rect 66805 265024 68908 265026
rect 66805 264968 66810 265024
rect 66866 264968 68908 265024
rect 66805 264966 68908 264968
rect 253460 264966 254164 265026
rect 48221 264963 48287 264966
rect 66805 264963 66871 264966
rect 254158 264964 254164 264966
rect 254228 264964 254234 265028
rect 268377 264890 268443 264893
rect 267690 264888 268443 264890
rect 267690 264832 268382 264888
rect 268438 264832 268443 264888
rect 267690 264830 268443 264832
rect 100753 264754 100819 264757
rect 98716 264752 100819 264754
rect 98716 264696 100758 264752
rect 100814 264696 100819 264752
rect 98716 264694 100819 264696
rect 100753 264691 100819 264694
rect 253430 264346 253490 264588
rect 266353 264346 266419 264349
rect 267690 264346 267750 264830
rect 268377 264827 268443 264830
rect 253430 264344 267750 264346
rect 253430 264288 266358 264344
rect 266414 264288 267750 264344
rect 253430 264286 267750 264288
rect 266353 264283 266419 264286
rect 54845 264210 54911 264213
rect 56409 264210 56475 264213
rect 54845 264208 56475 264210
rect 54845 264152 54850 264208
rect 54906 264152 56414 264208
rect 56470 264152 56475 264208
rect 191005 264210 191071 264213
rect 268561 264210 268627 264213
rect 582649 264210 582715 264213
rect 191005 264208 193660 264210
rect 54845 264150 56475 264152
rect 54845 264147 54911 264150
rect 56409 264147 56475 264150
rect 61929 263666 61995 263669
rect 68878 263666 68938 264180
rect 191005 264152 191010 264208
rect 191066 264152 193660 264208
rect 191005 264150 193660 264152
rect 268561 264208 582715 264210
rect 268561 264152 268566 264208
rect 268622 264152 582654 264208
rect 582710 264152 582715 264208
rect 268561 264150 582715 264152
rect 191005 264147 191071 264150
rect 268561 264147 268627 264150
rect 582649 264147 582715 264150
rect 256601 264074 256667 264077
rect 253460 264072 256667 264074
rect 253460 264016 256606 264072
rect 256662 264016 256667 264072
rect 253460 264014 256667 264016
rect 256601 264011 256667 264014
rect 100753 263938 100819 263941
rect 98716 263936 100819 263938
rect 98716 263880 100758 263936
rect 100814 263880 100819 263936
rect 98716 263878 100819 263880
rect 100753 263875 100819 263878
rect 115013 263668 115079 263669
rect 115013 263666 115060 263668
rect 61929 263664 68938 263666
rect 61929 263608 61934 263664
rect 61990 263608 68938 263664
rect 61929 263606 68938 263608
rect 114968 263664 115060 263666
rect 114968 263608 115018 263664
rect 114968 263606 115060 263608
rect 61929 263603 61995 263606
rect 63358 263533 63418 263606
rect 115013 263604 115060 263606
rect 115124 263604 115130 263668
rect 126830 263604 126836 263668
rect 126900 263666 126906 263668
rect 127065 263666 127131 263669
rect 255405 263666 255471 263669
rect 126900 263664 127131 263666
rect 126900 263608 127070 263664
rect 127126 263608 127131 263664
rect 126900 263606 127131 263608
rect 253460 263664 255471 263666
rect 253460 263608 255410 263664
rect 255466 263608 255471 263664
rect 253460 263606 255471 263608
rect 126900 263604 126906 263606
rect 115013 263603 115079 263604
rect 127065 263603 127131 263606
rect 255405 263603 255471 263606
rect 63358 263528 63467 263533
rect 63358 263472 63406 263528
rect 63462 263472 63467 263528
rect 63358 263470 63467 263472
rect 63401 263467 63467 263470
rect 66621 263394 66687 263397
rect 66621 263392 68908 263394
rect 66621 263336 66626 263392
rect 66682 263336 68908 263392
rect 66621 263334 68908 263336
rect 66621 263331 66687 263334
rect 191189 263258 191255 263261
rect 255405 263258 255471 263261
rect 191189 263256 193660 263258
rect 191189 263200 191194 263256
rect 191250 263200 193660 263256
rect 191189 263198 193660 263200
rect 253460 263256 255471 263258
rect 253460 263200 255410 263256
rect 255466 263200 255471 263256
rect 253460 263198 255471 263200
rect 191189 263195 191255 263198
rect 255405 263195 255471 263198
rect 100753 263122 100819 263125
rect 263542 263122 263548 263124
rect 98716 263120 100819 263122
rect 98716 263064 100758 263120
rect 100814 263064 100819 263120
rect 98716 263062 100819 263064
rect 100753 263059 100819 263062
rect 253430 263062 263548 263122
rect 253430 262684 253490 263062
rect 263542 263060 263548 263062
rect 263612 263060 263618 263124
rect 66897 262578 66963 262581
rect 66897 262576 68908 262578
rect 66897 262520 66902 262576
rect 66958 262520 68908 262576
rect 66897 262518 68908 262520
rect 66897 262515 66963 262518
rect 100845 262306 100911 262309
rect 98716 262304 100911 262306
rect 98716 262248 100850 262304
rect 100906 262248 100911 262304
rect 98716 262246 100911 262248
rect 100845 262243 100911 262246
rect 191005 262306 191071 262309
rect 256734 262306 256740 262308
rect 191005 262304 193660 262306
rect 191005 262248 191010 262304
rect 191066 262248 193660 262304
rect 191005 262246 193660 262248
rect 253460 262246 256740 262306
rect 191005 262243 191071 262246
rect 256734 262244 256740 262246
rect 256804 262244 256810 262308
rect 98085 262170 98151 262173
rect 98637 262170 98703 262173
rect 98085 262168 98703 262170
rect 98085 262112 98090 262168
rect 98146 262112 98642 262168
rect 98698 262112 98703 262168
rect 98085 262110 98703 262112
rect 98085 262107 98151 262110
rect 98637 262107 98703 262110
rect 104341 262170 104407 262173
rect 105077 262170 105143 262173
rect 104341 262168 105143 262170
rect 104341 262112 104346 262168
rect 104402 262112 105082 262168
rect 105138 262112 105143 262168
rect 104341 262110 105143 262112
rect 104341 262107 104407 262110
rect 105077 262107 105143 262110
rect 255814 261898 255820 261900
rect 252908 261868 255820 261898
rect 252878 261838 255820 261868
rect 252878 261764 252938 261838
rect 255814 261836 255820 261838
rect 255884 261836 255890 261900
rect 34237 261490 34303 261493
rect 61878 261490 61884 261492
rect 34237 261488 61884 261490
rect 34237 261432 34242 261488
rect 34298 261432 61884 261488
rect 34237 261430 61884 261432
rect 34237 261427 34303 261430
rect 61878 261428 61884 261430
rect 61948 261490 61954 261492
rect 68878 261490 68938 261732
rect 252870 261700 252876 261764
rect 252940 261700 252946 261764
rect 100753 261490 100819 261493
rect 61948 261430 68938 261490
rect 98716 261488 100819 261490
rect 98716 261432 100758 261488
rect 100814 261432 100819 261488
rect 98716 261430 100819 261432
rect 61948 261428 61954 261430
rect 100753 261427 100819 261430
rect 191373 261354 191439 261357
rect 256877 261354 256943 261357
rect 191373 261352 193660 261354
rect 191373 261296 191378 261352
rect 191434 261296 193660 261352
rect 191373 261294 193660 261296
rect 253460 261352 256943 261354
rect 253460 261296 256882 261352
rect 256938 261296 256943 261352
rect 253460 261294 256943 261296
rect 191373 261291 191439 261294
rect 256877 261291 256943 261294
rect 98637 261082 98703 261085
rect 181529 261082 181595 261085
rect 98637 261080 181595 261082
rect 98637 261024 98642 261080
rect 98698 261024 181534 261080
rect 181590 261024 181595 261080
rect 98637 261022 181595 261024
rect 98637 261019 98703 261022
rect 181529 261019 181595 261022
rect 66713 260946 66779 260949
rect 259678 260946 259684 260948
rect 66713 260944 68908 260946
rect 66713 260888 66718 260944
rect 66774 260888 68908 260944
rect 66713 260886 68908 260888
rect 253460 260886 259684 260946
rect 66713 260883 66779 260886
rect 259678 260884 259684 260886
rect 259748 260884 259754 260948
rect 100845 260674 100911 260677
rect 98716 260672 100911 260674
rect 98716 260616 100850 260672
rect 100906 260616 100911 260672
rect 98716 260614 100911 260616
rect 100845 260611 100911 260614
rect 191741 260402 191807 260405
rect 191741 260400 193660 260402
rect 191741 260344 191746 260400
rect 191802 260344 193660 260400
rect 191741 260342 193660 260344
rect 191741 260339 191807 260342
rect 253430 260266 253490 260508
rect 253430 260206 258090 260266
rect 66437 260130 66503 260133
rect 258030 260130 258090 260206
rect 269297 260130 269363 260133
rect 309777 260130 309843 260133
rect 66437 260128 68908 260130
rect 66437 260072 66442 260128
rect 66498 260072 68908 260128
rect 66437 260070 68908 260072
rect 258030 260128 309843 260130
rect 258030 260072 269302 260128
rect 269358 260072 309782 260128
rect 309838 260072 309843 260128
rect 258030 260070 309843 260072
rect 66437 260067 66503 260070
rect 269297 260067 269363 260070
rect 309777 260067 309843 260070
rect 255262 259994 255268 259996
rect 253460 259934 255268 259994
rect 255262 259932 255268 259934
rect 255332 259994 255338 259996
rect 255865 259994 255931 259997
rect 255332 259992 255931 259994
rect 255332 259936 255870 259992
rect 255926 259936 255931 259992
rect 255332 259934 255931 259936
rect 255332 259932 255338 259934
rect 255865 259931 255931 259934
rect 98134 259589 98194 259828
rect 98085 259584 98194 259589
rect 255405 259586 255471 259589
rect 98085 259528 98090 259584
rect 98146 259528 98194 259584
rect 98085 259526 98194 259528
rect 253460 259584 255471 259586
rect 253460 259528 255410 259584
rect 255466 259528 255471 259584
rect 253460 259526 255471 259528
rect 98085 259523 98151 259526
rect 255405 259523 255471 259526
rect 57646 259388 57652 259452
rect 57716 259450 57722 259452
rect 59118 259450 59124 259452
rect 57716 259390 59124 259450
rect 57716 259388 57722 259390
rect 59118 259388 59124 259390
rect 59188 259388 59194 259452
rect 68185 258770 68251 258773
rect 68878 258770 68938 259284
rect 100845 259042 100911 259045
rect 98716 259040 100911 259042
rect 98716 258984 100850 259040
rect 100906 258984 100911 259040
rect 98716 258982 100911 258984
rect 100845 258979 100911 258982
rect 193397 258906 193463 258909
rect 193630 258906 193690 259420
rect 255405 259042 255471 259045
rect 253460 259040 255471 259042
rect 253460 258984 255410 259040
rect 255466 258984 255471 259040
rect 253460 258982 255471 258984
rect 255405 258979 255471 258982
rect 193397 258904 193690 258906
rect 193397 258848 193402 258904
rect 193458 258848 193690 258904
rect 193397 258846 193690 258848
rect 582465 258906 582531 258909
rect 583520 258906 584960 258996
rect 582465 258904 584960 258906
rect 582465 258848 582470 258904
rect 582526 258848 584960 258904
rect 582465 258846 584960 258848
rect 193397 258843 193463 258846
rect 582465 258843 582531 258846
rect 132585 258770 132651 258773
rect 133781 258770 133847 258773
rect 68185 258768 68938 258770
rect 68185 258712 68190 258768
rect 68246 258712 68938 258768
rect 68185 258710 68938 258712
rect 125550 258768 133847 258770
rect 125550 258712 132590 258768
rect 132646 258712 133786 258768
rect 133842 258712 133847 258768
rect 583520 258756 584960 258846
rect 125550 258710 133847 258712
rect 68185 258707 68251 258710
rect 57646 258164 57652 258228
rect 57716 258226 57722 258228
rect 68878 258226 68938 258468
rect 100753 258226 100819 258229
rect 57716 258166 68938 258226
rect 98716 258224 100819 258226
rect 98716 258168 100758 258224
rect 100814 258168 100819 258224
rect 98716 258166 100819 258168
rect 57716 258164 57722 258166
rect 100753 258163 100819 258166
rect 124438 258028 124444 258092
rect 124508 258028 124514 258092
rect 124446 257954 124506 258028
rect 125550 257954 125610 258710
rect 132585 258707 132651 258710
rect 133781 258707 133847 258710
rect 255497 258634 255563 258637
rect 253460 258632 255563 258634
rect 253460 258576 255502 258632
rect 255558 258576 255563 258632
rect 253460 258574 255563 258576
rect 255497 258571 255563 258574
rect 190637 258362 190703 258365
rect 190637 258360 193660 258362
rect 190637 258304 190642 258360
rect 190698 258304 193660 258360
rect 190637 258302 193660 258304
rect 190637 258299 190703 258302
rect 254526 258226 254532 258228
rect 253460 258166 254532 258226
rect 254526 258164 254532 258166
rect 254596 258164 254602 258228
rect 103470 257894 125610 257954
rect 66621 257682 66687 257685
rect 66621 257680 68908 257682
rect 66621 257624 66626 257680
rect 66682 257624 68908 257680
rect 66621 257622 68908 257624
rect 66621 257619 66687 257622
rect 100845 257410 100911 257413
rect 98716 257408 100911 257410
rect 98716 257352 100850 257408
rect 100906 257352 100911 257408
rect 98716 257350 100911 257352
rect 100845 257347 100911 257350
rect 101029 257274 101095 257277
rect 103470 257274 103530 257894
rect 255405 257682 255471 257685
rect 253460 257680 255471 257682
rect 253460 257624 255410 257680
rect 255466 257624 255471 257680
rect 253460 257622 255471 257624
rect 255405 257619 255471 257622
rect 191741 257410 191807 257413
rect 191741 257408 193660 257410
rect 191741 257352 191746 257408
rect 191802 257352 193660 257408
rect 191741 257350 193660 257352
rect 191741 257347 191807 257350
rect 101029 257272 103530 257274
rect 101029 257216 101034 257272
rect 101090 257216 103530 257272
rect 101029 257214 103530 257216
rect 157977 257274 158043 257277
rect 184289 257274 184355 257277
rect 267825 257274 267891 257277
rect 268561 257274 268627 257277
rect 157977 257272 184355 257274
rect 157977 257216 157982 257272
rect 158038 257216 184294 257272
rect 184350 257216 184355 257272
rect 157977 257214 184355 257216
rect 253460 257272 268627 257274
rect 253460 257216 267830 257272
rect 267886 257216 268566 257272
rect 268622 257216 268627 257272
rect 253460 257214 268627 257216
rect 101029 257211 101095 257214
rect 157977 257211 158043 257214
rect 184289 257211 184355 257214
rect 267825 257211 267891 257214
rect 268561 257211 268627 257214
rect 66345 256866 66411 256869
rect 258390 256866 258396 256868
rect 66345 256864 68908 256866
rect 66345 256808 66350 256864
rect 66406 256808 68908 256864
rect 66345 256806 68908 256808
rect 253460 256806 258396 256866
rect 66345 256803 66411 256806
rect 258390 256804 258396 256806
rect 258460 256804 258466 256868
rect 262254 256668 262260 256732
rect 262324 256730 262330 256732
rect 262673 256730 262739 256733
rect 262324 256728 262739 256730
rect 262324 256672 262678 256728
rect 262734 256672 262739 256728
rect 262324 256670 262739 256672
rect 262324 256668 262330 256670
rect 262673 256667 262739 256670
rect 100937 256594 101003 256597
rect 98716 256592 101003 256594
rect 98716 256536 100942 256592
rect 100998 256536 101003 256592
rect 98716 256534 101003 256536
rect 100937 256531 101003 256534
rect 106089 256324 106155 256325
rect 106038 256322 106044 256324
rect 105998 256262 106044 256322
rect 106108 256320 106155 256324
rect 106150 256264 106155 256320
rect 106038 256260 106044 256262
rect 106108 256260 106155 256264
rect 106089 256259 106155 256260
rect 66805 256050 66871 256053
rect 66805 256048 68908 256050
rect 66805 255992 66810 256048
rect 66866 255992 68908 256048
rect 66805 255990 68908 255992
rect 66805 255987 66871 255990
rect 100845 255778 100911 255781
rect 98716 255776 100911 255778
rect 98716 255720 100850 255776
rect 100906 255720 100911 255776
rect 98716 255718 100911 255720
rect 100845 255715 100911 255718
rect 189717 255778 189783 255781
rect 193630 255778 193690 256428
rect 255405 256322 255471 256325
rect 253460 256320 255471 256322
rect 253460 256264 255410 256320
rect 255466 256264 255471 256320
rect 253460 256262 255471 256264
rect 255405 256259 255471 256262
rect 258349 256052 258415 256053
rect 258349 256050 258396 256052
rect 258304 256048 258396 256050
rect 258304 255992 258354 256048
rect 258304 255990 258396 255992
rect 258349 255988 258396 255990
rect 258460 255988 258466 256052
rect 258349 255987 258415 255988
rect 255497 255914 255563 255917
rect 253460 255912 255563 255914
rect 253460 255856 255502 255912
rect 255558 255856 255563 255912
rect 253460 255854 255563 255856
rect 255497 255851 255563 255854
rect 189717 255776 193690 255778
rect 189717 255720 189722 255776
rect 189778 255720 193690 255776
rect 189717 255718 193690 255720
rect 189717 255715 189783 255718
rect 191741 255506 191807 255509
rect 191741 255504 193660 255506
rect 191741 255448 191746 255504
rect 191802 255448 193660 255504
rect 191741 255446 193660 255448
rect 191741 255443 191807 255446
rect 258390 255370 258396 255372
rect 253460 255310 258396 255370
rect 258390 255308 258396 255310
rect 258460 255308 258466 255372
rect 66805 255234 66871 255237
rect 66805 255232 68908 255234
rect 66805 255176 66810 255232
rect 66866 255176 68908 255232
rect 66805 255174 68908 255176
rect 66805 255171 66871 255174
rect 101489 254962 101555 254965
rect 255405 254962 255471 254965
rect 98716 254960 101555 254962
rect 98716 254904 101494 254960
rect 101550 254904 101555 254960
rect 98716 254902 101555 254904
rect 253460 254960 255471 254962
rect 253460 254904 255410 254960
rect 255466 254904 255471 254960
rect 253460 254902 255471 254904
rect 101489 254899 101555 254902
rect 255405 254899 255471 254902
rect 41270 254492 41276 254556
rect 41340 254554 41346 254556
rect 49509 254554 49575 254557
rect 41340 254552 49575 254554
rect 41340 254496 49514 254552
rect 49570 254496 49575 254552
rect 41340 254494 49575 254496
rect 41340 254492 41346 254494
rect 49509 254491 49575 254494
rect 191557 254554 191623 254557
rect 255589 254554 255655 254557
rect 255957 254554 256023 254557
rect 267917 254554 267983 254557
rect 191557 254552 193660 254554
rect 191557 254496 191562 254552
rect 191618 254496 193660 254552
rect 191557 254494 193660 254496
rect 253460 254552 256023 254554
rect 253460 254496 255594 254552
rect 255650 254496 255962 254552
rect 256018 254496 256023 254552
rect 253460 254494 256023 254496
rect 191557 254491 191623 254494
rect 255589 254491 255655 254494
rect 255957 254491 256023 254494
rect 258030 254552 267983 254554
rect 258030 254496 267922 254552
rect 267978 254496 267983 254552
rect 258030 254494 267983 254496
rect 258030 254418 258090 254494
rect 267917 254491 267983 254494
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 57830 253948 57836 254012
rect 57900 254010 57906 254012
rect 60365 254010 60431 254013
rect 68878 254010 68938 254388
rect 253430 254358 258090 254418
rect 101029 254146 101095 254149
rect 98716 254144 101095 254146
rect 98716 254088 101034 254144
rect 101090 254088 101095 254144
rect 98716 254086 101095 254088
rect 101029 254083 101095 254086
rect 57900 254008 68938 254010
rect 57900 253952 60370 254008
rect 60426 253952 68938 254008
rect 253430 253980 253490 254358
rect 57900 253950 68938 253952
rect 57900 253948 57906 253950
rect 60365 253947 60431 253950
rect 66989 253602 67055 253605
rect 191005 253602 191071 253605
rect 255497 253602 255563 253605
rect 66989 253600 68908 253602
rect 66989 253544 66994 253600
rect 67050 253544 68908 253600
rect 66989 253542 68908 253544
rect 191005 253600 193660 253602
rect 191005 253544 191010 253600
rect 191066 253544 193660 253600
rect 191005 253542 193660 253544
rect 253460 253600 255563 253602
rect 253460 253544 255502 253600
rect 255558 253544 255563 253600
rect 253460 253542 255563 253544
rect 66989 253539 67055 253542
rect 191005 253539 191071 253542
rect 255497 253539 255563 253542
rect 100702 253330 100708 253332
rect 98716 253270 100708 253330
rect 100702 253268 100708 253270
rect 100772 253268 100778 253332
rect 255405 253194 255471 253197
rect 253460 253192 255471 253194
rect 253460 253136 255410 253192
rect 255466 253136 255471 253192
rect 253460 253134 255471 253136
rect 255405 253131 255471 253134
rect 61837 252786 61903 252789
rect 64781 252786 64847 252789
rect 61837 252784 68908 252786
rect 61837 252728 61842 252784
rect 61898 252728 64786 252784
rect 64842 252728 68908 252784
rect 61837 252726 68908 252728
rect 61837 252723 61903 252726
rect 64781 252723 64847 252726
rect 191741 252650 191807 252653
rect 255681 252650 255747 252653
rect 191741 252648 193660 252650
rect 191741 252592 191746 252648
rect 191802 252592 193660 252648
rect 253092 252648 255747 252650
rect 253092 252620 255686 252648
rect 191741 252590 193660 252592
rect 253062 252592 255686 252620
rect 255742 252592 255747 252648
rect 253062 252590 255747 252592
rect 191741 252587 191807 252590
rect 99465 252514 99531 252517
rect 100385 252514 100451 252517
rect 98716 252512 100451 252514
rect 98716 252456 99470 252512
rect 99526 252456 100390 252512
rect 100446 252456 100451 252512
rect 98716 252454 100451 252456
rect 99465 252451 99531 252454
rect 100385 252451 100451 252454
rect 252921 252514 252987 252517
rect 253062 252514 253122 252590
rect 255681 252587 255747 252590
rect 252921 252512 253122 252514
rect 252921 252456 252926 252512
rect 252982 252456 253122 252512
rect 252921 252454 253122 252456
rect 252921 252451 252987 252454
rect 255497 252242 255563 252245
rect 253460 252240 255563 252242
rect 253460 252184 255502 252240
rect 255558 252184 255563 252240
rect 253460 252182 255563 252184
rect 255497 252179 255563 252182
rect 68878 251426 68938 251940
rect 125777 251834 125843 251837
rect 142981 251834 143047 251837
rect 255405 251834 255471 251837
rect 122790 251832 143047 251834
rect 122790 251776 125782 251832
rect 125838 251776 142986 251832
rect 143042 251776 143047 251832
rect 122790 251774 143047 251776
rect 253460 251832 255471 251834
rect 253460 251776 255410 251832
rect 255466 251776 255471 251832
rect 253460 251774 255471 251776
rect 64830 251366 68938 251426
rect 98686 251426 98746 251668
rect 122790 251426 122850 251774
rect 125777 251771 125843 251774
rect 142981 251771 143047 251774
rect 255405 251771 255471 251774
rect 262489 251834 262555 251837
rect 291837 251834 291903 251837
rect 262489 251832 291903 251834
rect 262489 251776 262494 251832
rect 262550 251776 291842 251832
rect 291898 251776 291903 251832
rect 262489 251774 291903 251776
rect 262489 251771 262555 251774
rect 291837 251771 291903 251774
rect 191557 251698 191623 251701
rect 191557 251696 193660 251698
rect 191557 251640 191562 251696
rect 191618 251640 193660 251696
rect 191557 251638 193660 251640
rect 191557 251635 191623 251638
rect 98686 251366 122850 251426
rect 59118 251228 59124 251292
rect 59188 251290 59194 251292
rect 63309 251290 63375 251293
rect 64830 251290 64890 251366
rect 255313 251290 255379 251293
rect 59188 251288 64890 251290
rect 59188 251232 63314 251288
rect 63370 251232 64890 251288
rect 59188 251230 64890 251232
rect 253460 251288 255379 251290
rect 253460 251232 255318 251288
rect 255374 251232 255379 251288
rect 253460 251230 255379 251232
rect 59188 251228 59194 251230
rect 63309 251227 63375 251230
rect 255313 251227 255379 251230
rect 66805 251154 66871 251157
rect 66805 251152 68908 251154
rect 66805 251096 66810 251152
rect 66866 251096 68908 251152
rect 66805 251094 68908 251096
rect 66805 251091 66871 251094
rect 100845 250882 100911 250885
rect 98716 250880 100911 250882
rect 98716 250824 100850 250880
rect 100906 250824 100911 250880
rect 98716 250822 100911 250824
rect 100845 250819 100911 250822
rect 191741 250746 191807 250749
rect 191741 250744 193660 250746
rect 191741 250688 191746 250744
rect 191802 250688 193660 250744
rect 191741 250686 193660 250688
rect 191741 250683 191807 250686
rect 253430 250610 253490 250852
rect 263869 250610 263935 250613
rect 253430 250608 263935 250610
rect 253430 250552 263874 250608
rect 263930 250552 263935 250608
rect 253430 250550 263935 250552
rect 263869 250547 263935 250550
rect 255313 250338 255379 250341
rect 253460 250336 255379 250338
rect 64873 249930 64939 249933
rect 66110 249930 66116 249932
rect 64873 249928 66116 249930
rect 64873 249872 64878 249928
rect 64934 249872 66116 249928
rect 64873 249870 66116 249872
rect 64873 249867 64939 249870
rect 66110 249868 66116 249870
rect 66180 249930 66186 249932
rect 68878 249930 68938 250308
rect 253460 250280 255318 250336
rect 255374 250280 255379 250336
rect 253460 250278 255379 250280
rect 255313 250275 255379 250278
rect 100845 250066 100911 250069
rect 98716 250064 100911 250066
rect 98716 250008 100850 250064
rect 100906 250008 100911 250064
rect 98716 250006 100911 250008
rect 100845 250003 100911 250006
rect 255405 249930 255471 249933
rect 66180 249870 68938 249930
rect 253460 249928 255471 249930
rect 253460 249872 255410 249928
rect 255466 249872 255471 249928
rect 253460 249870 255471 249872
rect 66180 249868 66186 249870
rect 255405 249867 255471 249870
rect 190637 249658 190703 249661
rect 190637 249656 193660 249658
rect 190637 249600 190642 249656
rect 190698 249600 193660 249656
rect 190637 249598 193660 249600
rect 190637 249595 190703 249598
rect 66713 249522 66779 249525
rect 66713 249520 68908 249522
rect 66713 249464 66718 249520
rect 66774 249464 68908 249520
rect 66713 249462 68908 249464
rect 66713 249459 66779 249462
rect 100845 249250 100911 249253
rect 98716 249248 100911 249250
rect 98716 249192 100850 249248
rect 100906 249192 100911 249248
rect 98716 249190 100911 249192
rect 253430 249250 253490 249492
rect 254577 249250 254643 249253
rect 253430 249248 254643 249250
rect 253430 249192 254582 249248
rect 254638 249192 254643 249248
rect 253430 249190 254643 249192
rect 100845 249187 100911 249190
rect 254577 249187 254643 249190
rect 106641 249114 106707 249117
rect 108246 249114 108252 249116
rect 106641 249112 108252 249114
rect 106641 249056 106646 249112
rect 106702 249056 108252 249112
rect 106641 249054 108252 249056
rect 106641 249051 106707 249054
rect 108246 249052 108252 249054
rect 108316 249052 108322 249116
rect 255313 248978 255379 248981
rect 253460 248976 255379 248978
rect 253460 248920 255318 248976
rect 255374 248920 255379 248976
rect 253460 248918 255379 248920
rect 255313 248915 255379 248918
rect 55213 248434 55279 248437
rect 56501 248434 56567 248437
rect 68878 248434 68938 248676
rect 189809 248570 189875 248573
rect 193630 248570 193690 248676
rect 255681 248570 255747 248573
rect 189809 248568 193690 248570
rect 189809 248512 189814 248568
rect 189870 248512 193690 248568
rect 189809 248510 193690 248512
rect 253460 248568 255747 248570
rect 253460 248512 255686 248568
rect 255742 248512 255747 248568
rect 253460 248510 255747 248512
rect 189809 248507 189875 248510
rect 255681 248507 255747 248510
rect 100937 248434 101003 248437
rect 55213 248432 68938 248434
rect 55213 248376 55218 248432
rect 55274 248376 56506 248432
rect 56562 248376 68938 248432
rect 55213 248374 68938 248376
rect 98716 248432 101003 248434
rect 98716 248376 100942 248432
rect 100998 248376 101003 248432
rect 98716 248374 101003 248376
rect 55213 248371 55279 248374
rect 56501 248371 56567 248374
rect 100937 248371 101003 248374
rect 99230 248236 99236 248300
rect 99300 248298 99306 248300
rect 143533 248298 143599 248301
rect 99300 248296 143599 248298
rect 99300 248240 143538 248296
rect 143594 248240 143599 248296
rect 99300 248238 143599 248240
rect 99300 248236 99306 248238
rect 143533 248235 143599 248238
rect 253246 247893 253306 248132
rect 253197 247888 253306 247893
rect 68878 247346 68938 247860
rect 253197 247832 253202 247888
rect 253258 247832 253306 247888
rect 253197 247830 253306 247832
rect 253197 247827 253263 247830
rect 191741 247754 191807 247757
rect 191741 247752 193660 247754
rect 191741 247696 191746 247752
rect 191802 247696 193660 247752
rect 191741 247694 193660 247696
rect 191741 247691 191807 247694
rect 100845 247618 100911 247621
rect 98716 247616 100911 247618
rect 98716 247560 100850 247616
rect 100906 247560 100911 247616
rect 98716 247558 100911 247560
rect 100845 247555 100911 247558
rect 143533 247618 143599 247621
rect 192334 247618 192340 247620
rect 143533 247616 192340 247618
rect 143533 247560 143538 247616
rect 143594 247560 192340 247616
rect 143533 247558 192340 247560
rect 143533 247555 143599 247558
rect 192334 247556 192340 247558
rect 192404 247556 192410 247620
rect 255405 247618 255471 247621
rect 253460 247616 255471 247618
rect 253460 247560 255410 247616
rect 255466 247560 255471 247616
rect 253460 247558 255471 247560
rect 255405 247555 255471 247558
rect 64830 247286 68938 247346
rect 52453 247210 52519 247213
rect 53557 247210 53623 247213
rect 64830 247210 64890 247286
rect 258349 247210 258415 247213
rect 52453 247208 64890 247210
rect 52453 247152 52458 247208
rect 52514 247152 53562 247208
rect 53618 247152 64890 247208
rect 52453 247150 64890 247152
rect 253460 247208 258415 247210
rect 253460 247152 258354 247208
rect 258410 247152 258415 247208
rect 253460 247150 258415 247152
rect 52453 247147 52519 247150
rect 53557 247147 53623 247150
rect 258349 247147 258415 247150
rect 67449 247074 67515 247077
rect 67449 247072 68908 247074
rect 67449 247016 67454 247072
rect 67510 247016 68908 247072
rect 67449 247014 68908 247016
rect 67449 247011 67515 247014
rect 109534 247012 109540 247076
rect 109604 247074 109610 247076
rect 184381 247074 184447 247077
rect 109604 247072 184447 247074
rect 109604 247016 184386 247072
rect 184442 247016 184447 247072
rect 109604 247014 184447 247016
rect 109604 247012 109610 247014
rect 184381 247011 184447 247014
rect 100845 246802 100911 246805
rect 255313 246802 255379 246805
rect 98716 246800 100911 246802
rect 98716 246744 100850 246800
rect 100906 246744 100911 246800
rect 253460 246800 255379 246802
rect 98716 246742 100911 246744
rect 100845 246739 100911 246742
rect 57697 246258 57763 246261
rect 66662 246258 66668 246260
rect 57697 246256 66668 246258
rect 57697 246200 57702 246256
rect 57758 246200 66668 246256
rect 57697 246198 66668 246200
rect 57697 246195 57763 246198
rect 66662 246196 66668 246198
rect 66732 246196 66738 246260
rect 66989 246258 67055 246261
rect 109033 246258 109099 246261
rect 111006 246258 111012 246260
rect 66989 246256 68908 246258
rect 66989 246200 66994 246256
rect 67050 246200 68908 246256
rect 66989 246198 68908 246200
rect 109033 246256 111012 246258
rect 109033 246200 109038 246256
rect 109094 246200 111012 246256
rect 109033 246198 111012 246200
rect 66989 246195 67055 246198
rect 109033 246195 109099 246198
rect 111006 246196 111012 246198
rect 111076 246258 111082 246260
rect 120165 246258 120231 246261
rect 193438 246258 193444 246260
rect 111076 246256 120231 246258
rect 111076 246200 120170 246256
rect 120226 246200 120231 246256
rect 111076 246198 120231 246200
rect 111076 246196 111082 246198
rect 120165 246195 120231 246198
rect 180750 246198 193444 246258
rect 111190 246060 111196 246124
rect 111260 246122 111266 246124
rect 180750 246122 180810 246198
rect 193438 246196 193444 246198
rect 193508 246196 193514 246260
rect 193630 246122 193690 246772
rect 253460 246744 255318 246800
rect 255374 246744 255379 246800
rect 253460 246742 255379 246744
rect 255313 246739 255379 246742
rect 111260 246062 180810 246122
rect 191422 246062 193690 246122
rect 253062 246125 253122 246228
rect 253062 246120 253171 246125
rect 253062 246064 253110 246120
rect 253166 246064 253171 246120
rect 253062 246062 253171 246064
rect 111260 246060 111266 246062
rect 100845 245986 100911 245989
rect 98716 245984 100911 245986
rect 98716 245928 100850 245984
rect 100906 245928 100911 245984
rect 98716 245926 100911 245928
rect 100845 245923 100911 245926
rect 189901 245714 189967 245717
rect 191422 245714 191482 246062
rect 253105 246059 253171 246062
rect 191557 245850 191623 245853
rect 255405 245850 255471 245853
rect 191557 245848 193660 245850
rect 191557 245792 191562 245848
rect 191618 245792 193660 245848
rect 191557 245790 193660 245792
rect 253460 245848 255471 245850
rect 253460 245792 255410 245848
rect 255466 245792 255471 245848
rect 253460 245790 255471 245792
rect 191557 245787 191623 245790
rect 255405 245787 255471 245790
rect 189901 245712 191482 245714
rect 189901 245656 189906 245712
rect 189962 245656 191482 245712
rect 189901 245654 191482 245656
rect 189901 245651 189967 245654
rect 582373 245578 582439 245581
rect 583520 245578 584960 245668
rect 582373 245576 584960 245578
rect 582373 245520 582378 245576
rect 582434 245520 584960 245576
rect 582373 245518 584960 245520
rect 582373 245515 582439 245518
rect 583520 245428 584960 245518
rect 68878 244898 68938 245412
rect 255497 245306 255563 245309
rect 253460 245304 255563 245306
rect 253460 245248 255502 245304
rect 255558 245248 255563 245304
rect 253460 245246 255563 245248
rect 255497 245243 255563 245246
rect 100845 245170 100911 245173
rect 98716 245168 100911 245170
rect 98716 245112 100850 245168
rect 100906 245112 100911 245168
rect 98716 245110 100911 245112
rect 100845 245107 100911 245110
rect 64830 244838 68938 244898
rect 48037 244490 48103 244493
rect 64830 244490 64890 244838
rect 108246 244836 108252 244900
rect 108316 244898 108322 244900
rect 135345 244898 135411 244901
rect 108316 244896 135411 244898
rect 108316 244840 135350 244896
rect 135406 244840 135411 244896
rect 108316 244838 135411 244840
rect 108316 244836 108322 244838
rect 135345 244835 135411 244838
rect 191046 244836 191052 244900
rect 191116 244898 191122 244900
rect 255589 244898 255655 244901
rect 191116 244838 193660 244898
rect 253460 244896 255655 244898
rect 253460 244840 255594 244896
rect 255650 244840 255655 244896
rect 253460 244838 255655 244840
rect 191116 244836 191122 244838
rect 255589 244835 255655 244838
rect 253606 244700 253612 244764
rect 253676 244762 253682 244764
rect 255262 244762 255268 244764
rect 253676 244702 255268 244762
rect 253676 244700 253682 244702
rect 255262 244700 255268 244702
rect 255332 244700 255338 244764
rect 66897 244626 66963 244629
rect 66897 244624 68908 244626
rect 66897 244568 66902 244624
rect 66958 244568 68908 244624
rect 66897 244566 68908 244568
rect 66897 244563 66963 244566
rect 255262 244490 255268 244492
rect 48037 244488 64890 244490
rect 48037 244432 48042 244488
rect 48098 244432 64890 244488
rect 48037 244430 64890 244432
rect 253460 244430 255268 244490
rect 48037 244427 48103 244430
rect 255262 244428 255268 244430
rect 255332 244428 255338 244492
rect 100937 244354 101003 244357
rect 124305 244356 124371 244357
rect 98716 244352 101003 244354
rect 98716 244296 100942 244352
rect 100998 244296 101003 244352
rect 98716 244294 101003 244296
rect 100937 244291 101003 244294
rect 124254 244292 124260 244356
rect 124324 244354 124371 244356
rect 255313 244354 255379 244357
rect 259494 244354 259500 244356
rect 124324 244352 124416 244354
rect 124366 244296 124416 244352
rect 124324 244294 124416 244296
rect 255313 244352 259500 244354
rect 255313 244296 255318 244352
rect 255374 244296 259500 244352
rect 255313 244294 259500 244296
rect 124324 244292 124371 244294
rect 124305 244291 124371 244292
rect 255313 244291 255379 244294
rect 259494 244292 259500 244294
rect 259564 244354 259570 244356
rect 260741 244354 260807 244357
rect 259564 244352 260807 244354
rect 259564 244296 260746 244352
rect 260802 244296 260807 244352
rect 259564 244294 260807 244296
rect 259564 244292 259570 244294
rect 260741 244291 260807 244294
rect 191741 243946 191807 243949
rect 191741 243944 193660 243946
rect 191741 243888 191746 243944
rect 191802 243888 193660 243944
rect 191741 243886 193660 243888
rect 191741 243883 191807 243886
rect 253062 243813 253122 243916
rect 66805 243810 66871 243813
rect 66805 243808 68908 243810
rect 66805 243752 66810 243808
rect 66866 243752 68908 243808
rect 66805 243750 68908 243752
rect 253013 243808 253122 243813
rect 253013 243752 253018 243808
rect 253074 243752 253122 243808
rect 253013 243750 253122 243752
rect 66805 243747 66871 243750
rect 253013 243747 253079 243750
rect 100886 243538 100892 243540
rect 98716 243478 100892 243538
rect 100886 243476 100892 243478
rect 100956 243476 100962 243540
rect 255405 243538 255471 243541
rect 253460 243536 255471 243538
rect 253460 243480 255410 243536
rect 255466 243480 255471 243536
rect 253460 243478 255471 243480
rect 255405 243475 255471 243478
rect 255814 243130 255820 243132
rect 253460 243070 255820 243130
rect 255814 243068 255820 243070
rect 255884 243068 255890 243132
rect 66110 242932 66116 242996
rect 66180 242994 66186 242996
rect 66662 242994 66668 242996
rect 66180 242934 66668 242994
rect 66180 242932 66186 242934
rect 66662 242932 66668 242934
rect 66732 242994 66738 242996
rect 66732 242934 68908 242994
rect 66732 242932 66738 242934
rect 191230 242932 191236 242996
rect 191300 242994 191306 242996
rect 191300 242934 193660 242994
rect 191300 242932 191306 242934
rect 160921 242858 160987 242861
rect 193673 242858 193739 242861
rect 160921 242856 193739 242858
rect 160921 242800 160926 242856
rect 160982 242800 193678 242856
rect 193734 242800 193739 242856
rect 160921 242798 193739 242800
rect 160921 242795 160987 242798
rect 193673 242795 193739 242798
rect 100845 242722 100911 242725
rect 98716 242720 100911 242722
rect 98716 242664 100850 242720
rect 100906 242664 100911 242720
rect 98716 242662 100911 242664
rect 100845 242659 100911 242662
rect 255313 242586 255379 242589
rect 253460 242584 255379 242586
rect 253460 242528 255318 242584
rect 255374 242528 255379 242584
rect 253460 242526 255379 242528
rect 255313 242523 255379 242526
rect 255957 242178 256023 242181
rect 253460 242176 256023 242178
rect 65926 241708 65932 241772
rect 65996 241770 66002 241772
rect 68553 241770 68619 241773
rect 65996 241768 68619 241770
rect 65996 241712 68558 241768
rect 68614 241712 68619 241768
rect 65996 241710 68619 241712
rect 65996 241708 66002 241710
rect 68553 241707 68619 241710
rect 61694 241572 61700 241636
rect 61764 241634 61770 241636
rect 64781 241634 64847 241637
rect 68878 241634 68938 242148
rect 253460 242120 255962 242176
rect 256018 242120 256023 242176
rect 253460 242118 256023 242120
rect 255957 242115 256023 242118
rect 253013 242042 253079 242045
rect 255405 242042 255471 242045
rect 253013 242040 255471 242042
rect 100845 241906 100911 241909
rect 98716 241904 100911 241906
rect 98716 241848 100850 241904
rect 100906 241848 100911 241904
rect 98716 241846 100911 241848
rect 100845 241843 100911 241846
rect 70117 241772 70183 241773
rect 70117 241770 70164 241772
rect 70072 241768 70164 241770
rect 70072 241712 70122 241768
rect 70072 241710 70164 241712
rect 70117 241708 70164 241710
rect 70228 241708 70234 241772
rect 70894 241708 70900 241772
rect 70964 241770 70970 241772
rect 71129 241770 71195 241773
rect 71446 241770 71452 241772
rect 70964 241768 71452 241770
rect 70964 241712 71134 241768
rect 71190 241712 71452 241768
rect 70964 241710 71452 241712
rect 70964 241708 70970 241710
rect 70117 241707 70183 241708
rect 71129 241707 71195 241710
rect 71446 241708 71452 241710
rect 71516 241708 71522 241772
rect 72785 241770 72851 241773
rect 74257 241772 74323 241773
rect 91553 241772 91619 241773
rect 72918 241770 72924 241772
rect 72785 241768 72924 241770
rect 72785 241712 72790 241768
rect 72846 241712 72924 241768
rect 72785 241710 72924 241712
rect 72785 241707 72851 241710
rect 72918 241708 72924 241710
rect 72988 241708 72994 241772
rect 74206 241708 74212 241772
rect 74276 241770 74323 241772
rect 74276 241768 74368 241770
rect 74318 241712 74368 241768
rect 74276 241710 74368 241712
rect 74276 241708 74323 241710
rect 91502 241708 91508 241772
rect 91572 241770 91619 241772
rect 95877 241770 95943 241773
rect 102726 241770 102732 241772
rect 91572 241768 91664 241770
rect 91614 241712 91664 241768
rect 91572 241710 91664 241712
rect 95877 241768 102732 241770
rect 95877 241712 95882 241768
rect 95938 241712 102732 241768
rect 95877 241710 102732 241712
rect 91572 241708 91619 241710
rect 74257 241707 74323 241708
rect 91553 241707 91619 241708
rect 95877 241707 95943 241710
rect 102726 241708 102732 241710
rect 102796 241708 102802 241772
rect 94957 241636 95023 241637
rect 94957 241634 95004 241636
rect 61764 241632 68938 241634
rect 61764 241576 64786 241632
rect 64842 241576 68938 241632
rect 61764 241574 68938 241576
rect 94912 241632 95004 241634
rect 94912 241576 94962 241632
rect 94912 241574 95004 241576
rect 61764 241572 61770 241574
rect 64781 241571 64847 241574
rect 94957 241572 95004 241574
rect 95068 241572 95074 241636
rect 178677 241634 178743 241637
rect 193630 241634 193690 242012
rect 253013 241984 253018 242040
rect 253074 241984 255410 242040
rect 255466 241984 255471 242040
rect 253013 241982 255471 241984
rect 253013 241979 253079 241982
rect 255405 241979 255471 241982
rect 255405 241770 255471 241773
rect 253460 241768 255471 241770
rect 253460 241712 255410 241768
rect 255466 241712 255471 241768
rect 253460 241710 255471 241712
rect 255405 241707 255471 241710
rect 178677 241632 193690 241634
rect 178677 241576 178682 241632
rect 178738 241576 193690 241632
rect 178677 241574 193690 241576
rect 94957 241571 95023 241572
rect 178677 241571 178743 241574
rect 67766 241436 67772 241500
rect 67836 241498 67842 241500
rect 68369 241498 68435 241501
rect 67836 241496 68435 241498
rect 67836 241440 68374 241496
rect 68430 241440 68435 241496
rect 67836 241438 68435 241440
rect 67836 241436 67842 241438
rect 68369 241435 68435 241438
rect 76879 241498 76945 241501
rect 107694 241498 107700 241500
rect 76879 241496 107700 241498
rect 76879 241440 76884 241496
rect 76940 241440 107700 241496
rect 76879 241438 107700 241440
rect 76879 241435 76945 241438
rect 107694 241436 107700 241438
rect 107764 241498 107770 241500
rect 253974 241498 253980 241500
rect 107764 241438 253980 241498
rect 107764 241436 107770 241438
rect 253974 241436 253980 241438
rect 254044 241436 254050 241500
rect 67633 241362 67699 241365
rect 68783 241362 68849 241365
rect 126237 241362 126303 241365
rect 67633 241360 126303 241362
rect 67633 241304 67638 241360
rect 67694 241304 68788 241360
rect 68844 241304 126242 241360
rect 126298 241304 126303 241360
rect 67633 241302 126303 241304
rect 67633 241299 67699 241302
rect 68783 241299 68849 241302
rect 126237 241299 126303 241302
rect 142889 241362 142955 241365
rect 256877 241362 256943 241365
rect 142889 241360 256943 241362
rect 142889 241304 142894 241360
rect 142950 241304 256882 241360
rect 256938 241304 256943 241360
rect 142889 241302 256943 241304
rect 142889 241299 142955 241302
rect 256877 241299 256943 241302
rect 250529 241226 250595 241229
rect 253606 241226 253612 241228
rect 250529 241224 253612 241226
rect -960 241090 480 241180
rect 250529 241168 250534 241224
rect 250590 241168 253612 241224
rect 250529 241166 253612 241168
rect 250529 241163 250595 241166
rect 253606 241164 253612 241166
rect 253676 241164 253682 241228
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 64137 240818 64203 240821
rect 70577 240818 70643 240821
rect 64137 240816 70643 240818
rect 64137 240760 64142 240816
rect 64198 240760 70582 240816
rect 70638 240760 70643 240816
rect 64137 240758 70643 240760
rect 64137 240755 64203 240758
rect 70577 240755 70643 240758
rect 253606 240756 253612 240820
rect 253676 240818 253682 240820
rect 266629 240818 266695 240821
rect 253676 240816 266695 240818
rect 253676 240760 266634 240816
rect 266690 240760 266695 240816
rect 253676 240758 266695 240760
rect 253676 240756 253682 240758
rect 266629 240755 266695 240758
rect 78029 240274 78095 240277
rect 78029 240272 78138 240274
rect 78029 240216 78034 240272
rect 78090 240216 78138 240272
rect 78029 240211 78138 240216
rect 65977 240138 66043 240141
rect 69381 240138 69447 240141
rect 69790 240138 69796 240140
rect 65977 240136 69796 240138
rect 65977 240080 65982 240136
rect 66038 240080 69386 240136
rect 69442 240080 69796 240136
rect 65977 240078 69796 240080
rect 65977 240075 66043 240078
rect 69381 240075 69447 240078
rect 69790 240076 69796 240078
rect 69860 240076 69866 240140
rect 70393 240138 70459 240141
rect 71037 240138 71103 240141
rect 70393 240136 71103 240138
rect 70393 240080 70398 240136
rect 70454 240080 71042 240136
rect 71098 240080 71103 240136
rect 70393 240078 71103 240080
rect 78078 240138 78138 240211
rect 82077 240138 82143 240141
rect 78078 240136 82143 240138
rect 78078 240080 82082 240136
rect 82138 240080 82143 240136
rect 78078 240078 82143 240080
rect 70393 240075 70459 240078
rect 71037 240075 71103 240078
rect 82077 240075 82143 240078
rect 97809 240138 97875 240141
rect 104157 240138 104223 240141
rect 220813 240140 220879 240141
rect 234705 240140 234771 240141
rect 220813 240138 220860 240140
rect 97809 240136 104223 240138
rect 97809 240080 97814 240136
rect 97870 240080 104162 240136
rect 104218 240080 104223 240136
rect 97809 240078 104223 240080
rect 97809 240075 97875 240078
rect 104157 240075 104223 240078
rect 113130 240078 219450 240138
rect 220768 240136 220860 240138
rect 220768 240080 220818 240136
rect 220768 240078 220860 240080
rect 55070 239940 55076 240004
rect 55140 240002 55146 240004
rect 72417 240002 72483 240005
rect 72693 240002 72759 240005
rect 55140 240000 72759 240002
rect 55140 239944 72422 240000
rect 72478 239944 72698 240000
rect 72754 239944 72759 240000
rect 55140 239942 72759 239944
rect 55140 239940 55146 239942
rect 72417 239939 72483 239942
rect 72693 239939 72759 239942
rect 85481 240002 85547 240005
rect 86861 240002 86927 240005
rect 107653 240002 107719 240005
rect 113130 240002 113190 240078
rect 85481 240000 113190 240002
rect 85481 239944 85486 240000
rect 85542 239944 86866 240000
rect 86922 239944 107658 240000
rect 107714 239944 113190 240000
rect 85481 239942 113190 239944
rect 187141 240002 187207 240005
rect 204897 240002 204963 240005
rect 187141 240000 204963 240002
rect 187141 239944 187146 240000
rect 187202 239944 204902 240000
rect 204958 239944 204963 240000
rect 187141 239942 204963 239944
rect 85481 239939 85547 239942
rect 86861 239939 86927 239942
rect 107653 239939 107719 239942
rect 187141 239939 187207 239942
rect 204897 239939 204963 239942
rect 206369 240002 206435 240005
rect 207054 240002 207060 240004
rect 206369 240000 207060 240002
rect 206369 239944 206374 240000
rect 206430 239944 207060 240000
rect 206369 239942 207060 239944
rect 206369 239939 206435 239942
rect 207054 239940 207060 239942
rect 207124 239940 207130 240004
rect 219390 240002 219450 240078
rect 220813 240076 220860 240078
rect 220924 240076 220930 240140
rect 234654 240138 234660 240140
rect 234614 240078 234660 240138
rect 234724 240136 234771 240140
rect 234766 240080 234771 240136
rect 234654 240076 234660 240078
rect 234724 240076 234771 240080
rect 220813 240075 220879 240076
rect 234705 240075 234771 240076
rect 227253 240002 227319 240005
rect 219390 240000 227319 240002
rect 219390 239944 227258 240000
rect 227314 239944 227319 240000
rect 219390 239942 227319 239944
rect 227253 239939 227319 239942
rect 43989 239866 44055 239869
rect 70393 239866 70459 239869
rect 43989 239864 70459 239866
rect 43989 239808 43994 239864
rect 44050 239808 70398 239864
rect 70454 239808 70459 239864
rect 43989 239806 70459 239808
rect 43989 239803 44055 239806
rect 70393 239803 70459 239806
rect 191833 239866 191899 239869
rect 192702 239866 192708 239868
rect 191833 239864 192708 239866
rect 191833 239808 191838 239864
rect 191894 239808 192708 239864
rect 191833 239806 192708 239808
rect 191833 239803 191899 239806
rect 192702 239804 192708 239806
rect 192772 239804 192778 239868
rect 246389 239594 246455 239597
rect 252502 239594 252508 239596
rect 246389 239592 252508 239594
rect 246389 239536 246394 239592
rect 246450 239536 252508 239592
rect 246389 239534 252508 239536
rect 246389 239531 246455 239534
rect 252502 239532 252508 239534
rect 252572 239532 252578 239596
rect 240777 239458 240843 239461
rect 259729 239458 259795 239461
rect 240777 239456 259795 239458
rect 240777 239400 240782 239456
rect 240838 239400 259734 239456
rect 259790 239400 259795 239456
rect 240777 239398 259795 239400
rect 240777 239395 240843 239398
rect 259729 239395 259795 239398
rect 74257 238778 74323 238781
rect 74625 238778 74691 238781
rect 74257 238776 74691 238778
rect 74257 238720 74262 238776
rect 74318 238720 74630 238776
rect 74686 238720 74691 238776
rect 74257 238718 74691 238720
rect 74257 238715 74323 238718
rect 74625 238715 74691 238718
rect 48221 238642 48287 238645
rect 252645 238642 252711 238645
rect 48221 238640 252711 238642
rect 48221 238584 48226 238640
rect 48282 238584 252650 238640
rect 252706 238584 252711 238640
rect 48221 238582 252711 238584
rect 48221 238579 48287 238582
rect 252645 238579 252711 238582
rect 193806 238444 193812 238508
rect 193876 238506 193882 238508
rect 250437 238506 250503 238509
rect 193876 238504 250503 238506
rect 193876 238448 250442 238504
rect 250498 238448 250503 238504
rect 193876 238446 250503 238448
rect 193876 238444 193882 238446
rect 250437 238443 250503 238446
rect 238661 238370 238727 238373
rect 238886 238370 238892 238372
rect 238616 238368 238892 238370
rect 238616 238312 238666 238368
rect 238722 238312 238892 238368
rect 238616 238310 238892 238312
rect 238661 238307 238727 238310
rect 238886 238308 238892 238310
rect 238956 238308 238962 238372
rect 102726 238036 102732 238100
rect 102796 238098 102802 238100
rect 118734 238098 118740 238100
rect 102796 238038 118740 238098
rect 102796 238036 102802 238038
rect 118734 238036 118740 238038
rect 118804 238036 118810 238100
rect 81433 237962 81499 237965
rect 107653 237962 107719 237965
rect 117957 237962 118023 237965
rect 81433 237960 118023 237962
rect 81433 237904 81438 237960
rect 81494 237904 107658 237960
rect 107714 237904 117962 237960
rect 118018 237904 118023 237960
rect 81433 237902 118023 237904
rect 81433 237899 81499 237902
rect 107653 237899 107719 237902
rect 117957 237899 118023 237902
rect 255262 237900 255268 237964
rect 255332 237962 255338 237964
rect 582833 237962 582899 237965
rect 255332 237960 582899 237962
rect 255332 237904 582838 237960
rect 582894 237904 582899 237960
rect 255332 237902 582899 237904
rect 255332 237900 255338 237902
rect 582833 237899 582899 237902
rect 47945 237418 48011 237421
rect 48221 237418 48287 237421
rect 47945 237416 48287 237418
rect 47945 237360 47950 237416
rect 48006 237360 48226 237416
rect 48282 237360 48287 237416
rect 47945 237358 48287 237360
rect 47945 237355 48011 237358
rect 48221 237355 48287 237358
rect 90909 237418 90975 237421
rect 91185 237418 91251 237421
rect 90909 237416 91251 237418
rect 90909 237360 90914 237416
rect 90970 237360 91190 237416
rect 91246 237360 91251 237416
rect 90909 237358 91251 237360
rect 90909 237355 90975 237358
rect 91185 237355 91251 237358
rect 242014 237356 242020 237420
rect 242084 237418 242090 237420
rect 244273 237418 244339 237421
rect 242084 237416 244339 237418
rect 242084 237360 244278 237416
rect 244334 237360 244339 237416
rect 242084 237358 244339 237360
rect 242084 237356 242090 237358
rect 244273 237355 244339 237358
rect 249057 237418 249123 237421
rect 255262 237418 255268 237420
rect 249057 237416 255268 237418
rect 249057 237360 249062 237416
rect 249118 237360 255268 237416
rect 249057 237358 255268 237360
rect 249057 237355 249123 237358
rect 255262 237356 255268 237358
rect 255332 237356 255338 237420
rect 59077 237282 59143 237285
rect 111190 237282 111196 237284
rect 59077 237280 111196 237282
rect 59077 237224 59082 237280
rect 59138 237224 111196 237280
rect 59077 237222 111196 237224
rect 59077 237219 59143 237222
rect 111190 237220 111196 237222
rect 111260 237220 111266 237284
rect 173341 237282 173407 237285
rect 253606 237282 253612 237284
rect 173341 237280 253612 237282
rect 173341 237224 173346 237280
rect 173402 237224 253612 237280
rect 173341 237222 253612 237224
rect 173341 237219 173407 237222
rect 253606 237220 253612 237222
rect 253676 237220 253682 237284
rect 89713 237146 89779 237149
rect 102777 237146 102843 237149
rect 89713 237144 102843 237146
rect 89713 237088 89718 237144
rect 89774 237088 102782 237144
rect 102838 237088 102843 237144
rect 89713 237086 102843 237088
rect 89713 237083 89779 237086
rect 102777 237083 102843 237086
rect 111558 236676 111564 236740
rect 111628 236738 111634 236740
rect 188521 236738 188587 236741
rect 111628 236736 188587 236738
rect 111628 236680 188526 236736
rect 188582 236680 188587 236736
rect 111628 236678 188587 236680
rect 111628 236676 111634 236678
rect 188521 236675 188587 236678
rect 105537 236602 105603 236605
rect 191373 236602 191439 236605
rect 105537 236600 191439 236602
rect 105537 236544 105542 236600
rect 105598 236544 191378 236600
rect 191434 236544 191439 236600
rect 105537 236542 191439 236544
rect 105537 236539 105603 236542
rect 191373 236539 191439 236542
rect 192477 236602 192543 236605
rect 285673 236602 285739 236605
rect 192477 236600 285739 236602
rect 192477 236544 192482 236600
rect 192538 236544 285678 236600
rect 285734 236544 285739 236600
rect 192477 236542 285739 236544
rect 192477 236539 192543 236542
rect 285673 236539 285739 236542
rect 258349 235922 258415 235925
rect 142110 235920 258415 235922
rect 142110 235864 258354 235920
rect 258410 235864 258415 235920
rect 142110 235862 258415 235864
rect 92657 235514 92723 235517
rect 96654 235514 96660 235516
rect 92657 235512 96660 235514
rect 92657 235456 92662 235512
rect 92718 235456 96660 235512
rect 92657 235454 96660 235456
rect 92657 235451 92723 235454
rect 96654 235452 96660 235454
rect 96724 235452 96730 235516
rect 101397 235514 101463 235517
rect 118734 235514 118740 235516
rect 101397 235512 118740 235514
rect 101397 235456 101402 235512
rect 101458 235456 118740 235512
rect 101397 235454 118740 235456
rect 101397 235451 101463 235454
rect 118734 235452 118740 235454
rect 118804 235514 118810 235516
rect 118804 235454 122850 235514
rect 118804 235452 118810 235454
rect 88333 235378 88399 235381
rect 117681 235378 117747 235381
rect 88333 235376 117747 235378
rect 88333 235320 88338 235376
rect 88394 235320 117686 235376
rect 117742 235320 117747 235376
rect 88333 235318 117747 235320
rect 122790 235378 122850 235454
rect 140773 235378 140839 235381
rect 142110 235378 142170 235862
rect 258349 235859 258415 235862
rect 192334 235724 192340 235788
rect 192404 235786 192410 235788
rect 255405 235786 255471 235789
rect 192404 235784 255471 235786
rect 192404 235728 255410 235784
rect 255466 235728 255471 235784
rect 192404 235726 255471 235728
rect 192404 235724 192410 235726
rect 255405 235723 255471 235726
rect 122790 235376 142170 235378
rect 122790 235320 140778 235376
rect 140834 235320 142170 235376
rect 122790 235318 142170 235320
rect 88333 235315 88399 235318
rect 117681 235315 117747 235318
rect 140773 235315 140839 235318
rect 15101 235242 15167 235245
rect 191230 235242 191236 235244
rect 15101 235240 191236 235242
rect 15101 235184 15106 235240
rect 15162 235184 191236 235240
rect 15101 235182 191236 235184
rect 15101 235179 15167 235182
rect 191230 235180 191236 235182
rect 191300 235180 191306 235244
rect 97901 234698 97967 234701
rect 99465 234698 99531 234701
rect 97901 234696 99531 234698
rect 97901 234640 97906 234696
rect 97962 234640 99470 234696
rect 99526 234640 99531 234696
rect 97901 234638 99531 234640
rect 97901 234635 97967 234638
rect 99465 234635 99531 234638
rect 255814 234636 255820 234700
rect 255884 234698 255890 234700
rect 582649 234698 582715 234701
rect 255884 234696 582715 234698
rect 255884 234640 582654 234696
rect 582710 234640 582715 234696
rect 255884 234638 582715 234640
rect 255884 234636 255890 234638
rect 582649 234635 582715 234638
rect 45277 234562 45343 234565
rect 78765 234562 78831 234565
rect 45277 234560 78831 234562
rect 45277 234504 45282 234560
rect 45338 234504 78770 234560
rect 78826 234504 78831 234560
rect 45277 234502 78831 234504
rect 45277 234499 45343 234502
rect 78765 234499 78831 234502
rect 114502 234500 114508 234564
rect 114572 234562 114578 234564
rect 114645 234562 114711 234565
rect 114572 234560 114711 234562
rect 114572 234504 114650 234560
rect 114706 234504 114711 234560
rect 114572 234502 114711 234504
rect 114572 234500 114578 234502
rect 114645 234499 114711 234502
rect 122925 234562 122991 234565
rect 129733 234562 129799 234565
rect 262254 234562 262260 234564
rect 122925 234560 262260 234562
rect 122925 234504 122930 234560
rect 122986 234504 129738 234560
rect 129794 234504 262260 234560
rect 122925 234502 262260 234504
rect 122925 234499 122991 234502
rect 129733 234499 129799 234502
rect 262254 234500 262260 234502
rect 262324 234500 262330 234564
rect 117998 234426 118004 234428
rect 93810 234366 118004 234426
rect 86769 234154 86835 234157
rect 93810 234154 93870 234366
rect 117998 234364 118004 234366
rect 118068 234364 118074 234428
rect 86769 234152 93870 234154
rect 86769 234096 86774 234152
rect 86830 234096 93870 234152
rect 86769 234094 93870 234096
rect 86769 234091 86835 234094
rect 100017 234018 100083 234021
rect 100017 234016 109050 234018
rect 100017 233960 100022 234016
rect 100078 233960 109050 234016
rect 100017 233958 109050 233960
rect 100017 233955 100083 233958
rect 71681 233882 71747 233885
rect 73102 233882 73108 233884
rect 71681 233880 73108 233882
rect 71681 233824 71686 233880
rect 71742 233824 73108 233880
rect 71681 233822 73108 233824
rect 71681 233819 71747 233822
rect 73102 233820 73108 233822
rect 73172 233820 73178 233884
rect 93853 233882 93919 233885
rect 98637 233882 98703 233885
rect 93853 233880 98703 233882
rect 93853 233824 93858 233880
rect 93914 233824 98642 233880
rect 98698 233824 98703 233880
rect 93853 233822 98703 233824
rect 93853 233819 93919 233822
rect 98637 233819 98703 233822
rect 99097 233882 99163 233885
rect 100886 233882 100892 233884
rect 99097 233880 100892 233882
rect 99097 233824 99102 233880
rect 99158 233824 100892 233880
rect 99097 233822 100892 233824
rect 99097 233819 99163 233822
rect 100886 233820 100892 233822
rect 100956 233820 100962 233884
rect 108990 233882 109050 233958
rect 122925 233882 122991 233885
rect 108990 233880 122991 233882
rect 108990 233824 122930 233880
rect 122986 233824 122991 233880
rect 108990 233822 122991 233824
rect 122925 233819 122991 233822
rect 85665 233338 85731 233341
rect 86769 233338 86835 233341
rect 85665 233336 86835 233338
rect 85665 233280 85670 233336
rect 85726 233280 86774 233336
rect 86830 233280 86835 233336
rect 85665 233278 86835 233280
rect 85665 233275 85731 233278
rect 86769 233275 86835 233278
rect 256734 233202 256740 233204
rect 122790 233142 256740 233202
rect 106774 232732 106780 232796
rect 106844 232794 106850 232796
rect 121678 232794 121684 232796
rect 106844 232734 121684 232794
rect 106844 232732 106850 232734
rect 121678 232732 121684 232734
rect 121748 232794 121754 232796
rect 122790 232794 122850 233142
rect 256734 233140 256740 233142
rect 256804 233140 256810 233204
rect 146293 233066 146359 233069
rect 260925 233066 260991 233069
rect 121748 232734 122850 232794
rect 142110 233064 260991 233066
rect 142110 233008 146298 233064
rect 146354 233008 260930 233064
rect 260986 233008 260991 233064
rect 142110 233006 260991 233008
rect 121748 232732 121754 232734
rect 68645 232658 68711 232661
rect 77569 232658 77635 232661
rect 68645 232656 77635 232658
rect 68645 232600 68650 232656
rect 68706 232600 77574 232656
rect 77630 232600 77635 232656
rect 68645 232598 77635 232600
rect 68645 232595 68711 232598
rect 77569 232595 77635 232598
rect 97993 232658 98059 232661
rect 129733 232658 129799 232661
rect 142110 232658 142170 233006
rect 146293 233003 146359 233006
rect 260925 233003 260991 233006
rect 97993 232656 142170 232658
rect 97993 232600 97998 232656
rect 98054 232600 129738 232656
rect 129794 232600 142170 232656
rect 97993 232598 142170 232600
rect 97993 232595 98059 232598
rect 129733 232595 129799 232598
rect 33041 232522 33107 232525
rect 189901 232522 189967 232525
rect 33041 232520 189967 232522
rect 33041 232464 33046 232520
rect 33102 232464 189906 232520
rect 189962 232464 189967 232520
rect 33041 232462 189967 232464
rect 33041 232459 33107 232462
rect 189901 232459 189967 232462
rect 582373 232386 582439 232389
rect 583520 232386 584960 232476
rect 582373 232384 584960 232386
rect 582373 232328 582378 232384
rect 582434 232328 584960 232384
rect 582373 232326 584960 232328
rect 582373 232323 582439 232326
rect 583520 232236 584960 232326
rect 116526 231842 116532 231844
rect 113130 231782 116532 231842
rect 85573 231298 85639 231301
rect 93894 231298 93900 231300
rect 85573 231296 93900 231298
rect 85573 231240 85578 231296
rect 85634 231240 93900 231296
rect 85573 231238 93900 231240
rect 85573 231235 85639 231238
rect 93894 231236 93900 231238
rect 93964 231298 93970 231300
rect 111742 231298 111748 231300
rect 93964 231238 111748 231298
rect 93964 231236 93970 231238
rect 111742 231236 111748 231238
rect 111812 231236 111818 231300
rect 85573 231162 85639 231165
rect 113130 231162 113190 231782
rect 116526 231780 116532 231782
rect 116596 231842 116602 231844
rect 258390 231842 258396 231844
rect 116596 231782 258396 231842
rect 116596 231780 116602 231782
rect 258390 231780 258396 231782
rect 258460 231780 258466 231844
rect 85573 231160 113190 231162
rect 85573 231104 85578 231160
rect 85634 231104 113190 231160
rect 85573 231102 113190 231104
rect 85573 231099 85639 231102
rect 72417 230618 72483 230621
rect 74533 230618 74599 230621
rect 255497 230618 255563 230621
rect 72417 230616 255563 230618
rect 72417 230560 72422 230616
rect 72478 230560 74538 230616
rect 74594 230560 255502 230616
rect 255558 230560 255563 230616
rect 72417 230558 255563 230560
rect 72417 230555 72483 230558
rect 74533 230555 74599 230558
rect 255497 230555 255563 230558
rect 61878 230420 61884 230484
rect 61948 230482 61954 230484
rect 269389 230482 269455 230485
rect 61948 230480 269455 230482
rect 61948 230424 269394 230480
rect 269450 230424 269455 230480
rect 61948 230422 269455 230424
rect 61948 230420 61954 230422
rect 269389 230419 269455 230422
rect 97441 230346 97507 230349
rect 99966 230346 99972 230348
rect 97441 230344 99972 230346
rect 97441 230288 97446 230344
rect 97502 230288 99972 230344
rect 97441 230286 99972 230288
rect 97441 230283 97507 230286
rect 99966 230284 99972 230286
rect 100036 230284 100042 230348
rect 100569 229802 100635 229805
rect 100702 229802 100708 229804
rect 100569 229800 100708 229802
rect 100569 229744 100574 229800
rect 100630 229744 100708 229800
rect 100569 229742 100708 229744
rect 100569 229739 100635 229742
rect 100702 229740 100708 229742
rect 100772 229740 100778 229804
rect 238661 229124 238727 229125
rect 238661 229122 238708 229124
rect 238616 229120 238708 229122
rect 238772 229122 238778 229124
rect 238616 229064 238666 229120
rect 238616 229062 238708 229064
rect 238661 229060 238708 229062
rect 238772 229062 238854 229122
rect 238772 229060 238778 229062
rect 238661 229059 238727 229060
rect 52085 228986 52151 228989
rect 262489 228986 262555 228989
rect 52085 228984 262555 228986
rect 52085 228928 52090 228984
rect 52146 228928 262494 228984
rect 262550 228928 262555 228984
rect 52085 228926 262555 228928
rect 52085 228923 52151 228926
rect 262489 228923 262555 228926
rect 103830 228850 103836 228852
rect 80010 228790 103836 228850
rect 79317 228306 79383 228309
rect 80010 228306 80070 228790
rect 103830 228788 103836 228790
rect 103900 228850 103906 228852
rect 234613 228850 234679 228853
rect 238661 228852 238727 228853
rect 238661 228850 238708 228852
rect 103900 228848 234679 228850
rect 103900 228792 234618 228848
rect 234674 228792 234679 228848
rect 103900 228790 234679 228792
rect 238616 228848 238708 228850
rect 238772 228850 238778 228852
rect 238616 228792 238666 228848
rect 238616 228790 238708 228792
rect 103900 228788 103906 228790
rect 234613 228787 234679 228790
rect 238661 228788 238708 228790
rect 238772 228790 238854 228850
rect 238772 228788 238778 228790
rect 238661 228787 238727 228788
rect 79317 228304 80070 228306
rect 79317 228248 79322 228304
rect 79378 228248 80070 228304
rect 79317 228246 80070 228248
rect 104801 228306 104867 228309
rect 214414 228306 214420 228308
rect 104801 228304 214420 228306
rect 104801 228248 104806 228304
rect 104862 228248 214420 228304
rect 104801 228246 214420 228248
rect 79317 228243 79383 228246
rect 104801 228243 104867 228246
rect 214414 228244 214420 228246
rect 214484 228244 214490 228308
rect -960 227884 480 228124
rect 92289 227762 92355 227765
rect 94681 227762 94747 227765
rect 92289 227760 94747 227762
rect 92289 227704 92294 227760
rect 92350 227704 94686 227760
rect 94742 227704 94747 227760
rect 92289 227702 94747 227704
rect 92289 227699 92355 227702
rect 94681 227699 94747 227702
rect 92289 227082 92355 227085
rect 95182 227082 95188 227084
rect 92289 227080 95188 227082
rect 92289 227024 92294 227080
rect 92350 227024 95188 227080
rect 92289 227022 95188 227024
rect 92289 227019 92355 227022
rect 95182 227020 95188 227022
rect 95252 227020 95258 227084
rect 200757 227082 200823 227085
rect 249241 227082 249307 227085
rect 200757 227080 249307 227082
rect 200757 227024 200762 227080
rect 200818 227024 249246 227080
rect 249302 227024 249307 227080
rect 200757 227022 249307 227024
rect 200757 227019 200823 227022
rect 249241 227019 249307 227022
rect 78581 226946 78647 226949
rect 259678 226946 259684 226948
rect 78581 226944 259684 226946
rect 78581 226888 78586 226944
rect 78642 226888 259684 226944
rect 78581 226886 259684 226888
rect 78581 226883 78647 226886
rect 259678 226884 259684 226886
rect 259748 226884 259754 226948
rect 60457 226266 60523 226269
rect 251817 226266 251883 226269
rect 60457 226264 251883 226266
rect 60457 226208 60462 226264
rect 60518 226208 251822 226264
rect 251878 226208 251883 226264
rect 60457 226206 251883 226208
rect 60457 226203 60523 226206
rect 251817 226203 251883 226206
rect 81525 226130 81591 226133
rect 115974 226130 115980 226132
rect 80010 226128 115980 226130
rect 80010 226072 81530 226128
rect 81586 226072 115980 226128
rect 80010 226070 115980 226072
rect 76557 225586 76623 225589
rect 80010 225586 80070 226070
rect 81525 226067 81591 226070
rect 115974 226068 115980 226070
rect 116044 226068 116050 226132
rect 103421 225994 103487 225997
rect 104934 225994 104940 225996
rect 103421 225992 104940 225994
rect 103421 225936 103426 225992
rect 103482 225936 104940 225992
rect 103421 225934 104940 225936
rect 103421 225931 103487 225934
rect 104934 225932 104940 225934
rect 105004 225932 105010 225996
rect 76557 225584 80070 225586
rect 76557 225528 76562 225584
rect 76618 225528 80070 225584
rect 76557 225526 80070 225528
rect 141417 225586 141483 225589
rect 216806 225586 216812 225588
rect 141417 225584 216812 225586
rect 141417 225528 141422 225584
rect 141478 225528 216812 225584
rect 141417 225526 216812 225528
rect 76557 225523 76623 225526
rect 141417 225523 141483 225526
rect 216806 225524 216812 225526
rect 216876 225524 216882 225588
rect 52177 224906 52243 224909
rect 259637 224906 259703 224909
rect 52177 224904 259703 224906
rect 52177 224848 52182 224904
rect 52238 224848 259642 224904
rect 259698 224848 259703 224904
rect 52177 224846 259703 224848
rect 52177 224843 52243 224846
rect 259637 224843 259703 224846
rect 268009 224770 268075 224773
rect 268377 224770 268443 224773
rect 113130 224768 268443 224770
rect 113130 224712 268014 224768
rect 268070 224712 268382 224768
rect 268438 224712 268443 224768
rect 113130 224710 268443 224712
rect 78857 224226 78923 224229
rect 110638 224226 110644 224228
rect 78857 224224 110644 224226
rect 78857 224168 78862 224224
rect 78918 224168 110644 224224
rect 78857 224166 110644 224168
rect 78857 224163 78923 224166
rect 110638 224164 110644 224166
rect 110708 224226 110714 224228
rect 113130 224226 113190 224710
rect 268009 224707 268075 224710
rect 268377 224707 268443 224710
rect 110708 224166 113190 224226
rect 115841 224226 115907 224229
rect 216070 224226 216076 224228
rect 115841 224224 216076 224226
rect 115841 224168 115846 224224
rect 115902 224168 216076 224224
rect 115841 224166 216076 224168
rect 110708 224164 110714 224166
rect 115841 224163 115907 224166
rect 216070 224164 216076 224166
rect 216140 224164 216146 224228
rect 49417 223546 49483 223549
rect 49601 223546 49667 223549
rect 270769 223546 270835 223549
rect 49417 223544 270835 223546
rect 49417 223488 49422 223544
rect 49478 223488 49606 223544
rect 49662 223488 270774 223544
rect 270830 223488 270835 223544
rect 49417 223486 270835 223488
rect 49417 223483 49483 223486
rect 49601 223483 49667 223486
rect 270769 223483 270835 223486
rect 4061 222866 4127 222869
rect 186814 222866 186820 222868
rect 4061 222864 186820 222866
rect 4061 222808 4066 222864
rect 4122 222808 186820 222864
rect 4061 222806 186820 222808
rect 4061 222803 4127 222806
rect 186814 222804 186820 222806
rect 186884 222804 186890 222868
rect 57605 222188 57671 222189
rect 57605 222186 57652 222188
rect 57560 222184 57652 222186
rect 57716 222186 57722 222188
rect 240777 222186 240843 222189
rect 57716 222184 240843 222186
rect 57560 222128 57610 222184
rect 57716 222128 240782 222184
rect 240838 222128 240843 222184
rect 57560 222126 57652 222128
rect 57605 222124 57652 222126
rect 57716 222126 240843 222128
rect 57716 222124 57722 222126
rect 57605 222123 57671 222124
rect 240777 222123 240843 222126
rect 126881 222052 126947 222053
rect 126830 222050 126836 222052
rect 126754 221990 126836 222050
rect 126900 222050 126947 222052
rect 258390 222050 258396 222052
rect 126900 222048 258396 222050
rect 126942 221992 258396 222048
rect 126830 221988 126836 221990
rect 126900 221990 258396 221992
rect 126900 221988 126947 221990
rect 258390 221988 258396 221990
rect 258460 221988 258466 222052
rect 126881 221987 126947 221988
rect 50705 220826 50771 220829
rect 267917 220826 267983 220829
rect 50705 220824 267983 220826
rect 50705 220768 50710 220824
rect 50766 220768 267922 220824
rect 267978 220768 267983 220824
rect 50705 220766 267983 220768
rect 50705 220763 50771 220766
rect 267917 220763 267983 220766
rect 92473 220690 92539 220693
rect 93710 220690 93716 220692
rect 92473 220688 93716 220690
rect 92473 220632 92478 220688
rect 92534 220632 93716 220688
rect 92473 220630 93716 220632
rect 92473 220627 92539 220630
rect 93710 220628 93716 220630
rect 93780 220690 93786 220692
rect 106406 220690 106412 220692
rect 93780 220630 106412 220690
rect 93780 220628 93786 220630
rect 106406 220628 106412 220630
rect 106476 220628 106482 220692
rect 263726 220690 263732 220692
rect 142110 220630 263732 220690
rect 96705 220282 96771 220285
rect 121678 220282 121684 220284
rect 96705 220280 121684 220282
rect 96705 220224 96710 220280
rect 96766 220224 121684 220280
rect 96705 220222 121684 220224
rect 96705 220219 96771 220222
rect 121678 220220 121684 220222
rect 121748 220282 121754 220284
rect 138013 220282 138079 220285
rect 142110 220282 142170 220630
rect 263726 220628 263732 220630
rect 263796 220628 263802 220692
rect 121748 220280 142170 220282
rect 121748 220224 138018 220280
rect 138074 220224 142170 220280
rect 121748 220222 142170 220224
rect 121748 220220 121754 220222
rect 138013 220219 138079 220222
rect 117078 220084 117084 220148
rect 117148 220146 117154 220148
rect 234838 220146 234844 220148
rect 117148 220086 234844 220146
rect 117148 220084 117154 220086
rect 234838 220084 234844 220086
rect 234908 220084 234914 220148
rect 238661 219466 238727 219469
rect 238886 219466 238892 219468
rect 238616 219464 238892 219466
rect 238616 219408 238666 219464
rect 238722 219408 238892 219464
rect 238616 219406 238892 219408
rect 238661 219403 238727 219406
rect 238886 219404 238892 219406
rect 238956 219404 238962 219468
rect 69974 219268 69980 219332
rect 70044 219330 70050 219332
rect 251909 219330 251975 219333
rect 70044 219328 251975 219330
rect 70044 219272 251914 219328
rect 251970 219272 251975 219328
rect 70044 219270 251975 219272
rect 70044 219268 70050 219270
rect 251909 219267 251975 219270
rect 131113 219194 131179 219197
rect 269297 219194 269363 219197
rect 131113 219192 269363 219194
rect 131113 219136 131118 219192
rect 131174 219136 269302 219192
rect 269358 219136 269363 219192
rect 131113 219134 269363 219136
rect 131113 219131 131179 219134
rect 269297 219131 269363 219134
rect 238661 219058 238727 219061
rect 238886 219058 238892 219060
rect 238616 219056 238892 219058
rect 238616 219000 238666 219056
rect 238722 219000 238892 219056
rect 238616 218998 238892 219000
rect 238661 218995 238727 218998
rect 238886 218996 238892 218998
rect 238956 218996 238962 219060
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 100569 218650 100635 218653
rect 125685 218650 125751 218653
rect 131113 218650 131179 218653
rect 100569 218648 131179 218650
rect 100569 218592 100574 218648
rect 100630 218592 125690 218648
rect 125746 218592 131118 218648
rect 131174 218592 131179 218648
rect 100569 218590 131179 218592
rect 100569 218587 100635 218590
rect 125685 218587 125751 218590
rect 131113 218587 131179 218590
rect 95877 217290 95943 217293
rect 244406 217290 244412 217292
rect 95877 217288 244412 217290
rect 95877 217232 95882 217288
rect 95938 217232 244412 217288
rect 95877 217230 244412 217232
rect 95877 217227 95943 217230
rect 244406 217228 244412 217230
rect 244476 217228 244482 217292
rect 95325 216746 95391 216749
rect 95877 216746 95943 216749
rect 95325 216744 95943 216746
rect 95325 216688 95330 216744
rect 95386 216688 95882 216744
rect 95938 216688 95943 216744
rect 95325 216686 95943 216688
rect 95325 216683 95391 216686
rect 95877 216683 95943 216686
rect 244406 216684 244412 216748
rect 244476 216746 244482 216748
rect 244917 216746 244983 216749
rect 244476 216744 244983 216746
rect 244476 216688 244922 216744
rect 244978 216688 244983 216744
rect 244476 216686 244983 216688
rect 244476 216684 244482 216686
rect 244917 216683 244983 216686
rect 42609 216610 42675 216613
rect 48037 216610 48103 216613
rect 246389 216610 246455 216613
rect 42609 216608 246455 216610
rect 42609 216552 42614 216608
rect 42670 216552 48042 216608
rect 48098 216552 246394 216608
rect 246450 216552 246455 216608
rect 42609 216550 246455 216552
rect 42609 216547 42675 216550
rect 48037 216547 48103 216550
rect 246389 216547 246455 216550
rect 134517 215930 134583 215933
rect 236494 215930 236500 215932
rect 134517 215928 236500 215930
rect 134517 215872 134522 215928
rect 134578 215872 236500 215928
rect 134517 215870 236500 215872
rect 134517 215867 134583 215870
rect 236494 215868 236500 215870
rect 236564 215868 236570 215932
rect 133822 215250 133828 215252
rect 122790 215190 133828 215250
rect -960 214978 480 215068
rect 3141 214978 3207 214981
rect -960 214976 3207 214978
rect -960 214920 3146 214976
rect 3202 214920 3207 214976
rect -960 214918 3207 214920
rect -960 214828 480 214918
rect 3141 214915 3207 214918
rect 99097 214706 99163 214709
rect 111885 214706 111951 214709
rect 122790 214706 122850 215190
rect 133822 215188 133828 215190
rect 133892 215250 133898 215252
rect 266353 215250 266419 215253
rect 133892 215248 266419 215250
rect 133892 215192 266358 215248
rect 266414 215192 266419 215248
rect 133892 215190 266419 215192
rect 133892 215188 133898 215190
rect 266353 215187 266419 215190
rect 99097 214704 122850 214706
rect 99097 214648 99102 214704
rect 99158 214648 111890 214704
rect 111946 214648 122850 214704
rect 99097 214646 122850 214648
rect 99097 214643 99163 214646
rect 111885 214643 111951 214646
rect 38561 214570 38627 214573
rect 221222 214570 221228 214572
rect 38561 214568 221228 214570
rect 38561 214512 38566 214568
rect 38622 214512 221228 214568
rect 38561 214510 221228 214512
rect 38561 214507 38627 214510
rect 221222 214508 221228 214510
rect 221292 214508 221298 214572
rect 139485 213890 139551 213893
rect 258257 213890 258323 213893
rect 139485 213888 258323 213890
rect 139485 213832 139490 213888
rect 139546 213832 258262 213888
rect 258318 213832 258323 213888
rect 139485 213830 258323 213832
rect 139485 213827 139551 213830
rect 258257 213827 258323 213830
rect 86217 213210 86283 213213
rect 139485 213210 139551 213213
rect 86217 213208 139551 213210
rect 86217 213152 86222 213208
rect 86278 213152 139490 213208
rect 139546 213152 139551 213208
rect 86217 213150 139551 213152
rect 86217 213147 86283 213150
rect 139485 213147 139551 213150
rect 188981 213210 189047 213213
rect 583477 213210 583543 213213
rect 188981 213208 583543 213210
rect 188981 213152 188986 213208
rect 189042 213152 583482 213208
rect 583538 213152 583543 213208
rect 188981 213150 583543 213152
rect 188981 213147 189047 213150
rect 583477 213147 583543 213150
rect 124305 212530 124371 212533
rect 262213 212530 262279 212533
rect 122790 212528 262279 212530
rect 122790 212472 124310 212528
rect 124366 212472 262218 212528
rect 262274 212472 262279 212528
rect 122790 212470 262279 212472
rect 108246 211924 108252 211988
rect 108316 211986 108322 211988
rect 122790 211986 122850 212470
rect 124305 212467 124371 212470
rect 262213 212467 262279 212470
rect 108316 211926 122850 211986
rect 108316 211924 108322 211926
rect 90817 211850 90883 211853
rect 128629 211852 128695 211853
rect 114502 211850 114508 211852
rect 90817 211848 114508 211850
rect 90817 211792 90822 211848
rect 90878 211792 114508 211848
rect 90817 211790 114508 211792
rect 90817 211787 90883 211790
rect 114502 211788 114508 211790
rect 114572 211850 114578 211852
rect 128629 211850 128676 211852
rect 114572 211848 128676 211850
rect 128740 211850 128746 211852
rect 114572 211792 128634 211848
rect 114572 211790 128676 211792
rect 114572 211788 114578 211790
rect 128629 211788 128676 211790
rect 128740 211790 128822 211850
rect 128740 211788 128746 211790
rect 128629 211787 128695 211788
rect 120349 211034 120415 211037
rect 120717 211034 120783 211037
rect 260833 211034 260899 211037
rect 120349 211032 260899 211034
rect 120349 210976 120354 211032
rect 120410 210976 120722 211032
rect 120778 210976 260838 211032
rect 260894 210976 260899 211032
rect 120349 210974 260899 210976
rect 120349 210971 120415 210974
rect 120717 210971 120783 210974
rect 260833 210971 260899 210974
rect 84009 210354 84075 210357
rect 104014 210354 104020 210356
rect 84009 210352 104020 210354
rect 84009 210296 84014 210352
rect 84070 210296 104020 210352
rect 84009 210294 104020 210296
rect 84009 210291 84075 210294
rect 104014 210292 104020 210294
rect 104084 210354 104090 210356
rect 120349 210354 120415 210357
rect 104084 210352 120415 210354
rect 104084 210296 120354 210352
rect 120410 210296 120415 210352
rect 104084 210294 120415 210296
rect 104084 210292 104090 210294
rect 120349 210291 120415 210294
rect 238661 209812 238727 209813
rect 238661 209810 238708 209812
rect 238616 209808 238708 209810
rect 238772 209810 238778 209812
rect 238616 209752 238666 209808
rect 238616 209750 238708 209752
rect 238661 209748 238708 209750
rect 238772 209750 238854 209810
rect 238772 209748 238778 209750
rect 238661 209747 238727 209748
rect 49509 209674 49575 209677
rect 255814 209674 255820 209676
rect 49509 209672 255820 209674
rect 49509 209616 49514 209672
rect 49570 209616 255820 209672
rect 49509 209614 255820 209616
rect 49509 209611 49575 209614
rect 255814 209612 255820 209614
rect 255884 209612 255890 209676
rect 238661 209538 238727 209541
rect 238886 209538 238892 209540
rect 238616 209536 238892 209538
rect 238616 209480 238666 209536
rect 238722 209480 238892 209536
rect 238616 209478 238892 209480
rect 238661 209475 238727 209478
rect 238886 209476 238892 209478
rect 238956 209476 238962 209540
rect 119061 208314 119127 208317
rect 273345 208314 273411 208317
rect 119061 208312 273411 208314
rect 119061 208256 119066 208312
rect 119122 208256 273350 208312
rect 273406 208256 273411 208312
rect 119061 208254 273411 208256
rect 119061 208251 119127 208254
rect 273345 208251 273411 208254
rect 128353 208178 128419 208181
rect 252737 208178 252803 208181
rect 128353 208176 252803 208178
rect 128353 208120 128358 208176
rect 128414 208120 252742 208176
rect 252798 208120 252803 208176
rect 128353 208118 252803 208120
rect 128353 208115 128419 208118
rect 252737 208115 252803 208118
rect 93761 207770 93827 207773
rect 109033 207770 109099 207773
rect 128353 207770 128419 207773
rect 93761 207768 128419 207770
rect 93761 207712 93766 207768
rect 93822 207712 109038 207768
rect 109094 207712 128358 207768
rect 128414 207712 128419 207768
rect 93761 207710 128419 207712
rect 93761 207707 93827 207710
rect 109033 207707 109099 207710
rect 128353 207707 128419 207710
rect 84193 207634 84259 207637
rect 104985 207634 105051 207637
rect 119061 207634 119127 207637
rect 84193 207632 119127 207634
rect 84193 207576 84198 207632
rect 84254 207576 104990 207632
rect 105046 207576 119066 207632
rect 119122 207576 119127 207632
rect 84193 207574 119127 207576
rect 84193 207571 84259 207574
rect 104985 207571 105051 207574
rect 119061 207571 119127 207574
rect 117405 206954 117471 206957
rect 257061 206954 257127 206957
rect 117405 206952 257127 206954
rect 117405 206896 117410 206952
rect 117466 206896 257066 206952
rect 257122 206896 257127 206952
rect 117405 206894 257127 206896
rect 117405 206891 117471 206894
rect 257061 206891 257127 206894
rect 259494 206818 259500 206820
rect 122790 206758 259500 206818
rect 90909 206410 90975 206413
rect 114553 206410 114619 206413
rect 117405 206410 117471 206413
rect 90909 206408 117471 206410
rect 90909 206352 90914 206408
rect 90970 206352 114558 206408
rect 114614 206352 117410 206408
rect 117466 206352 117471 206408
rect 90909 206350 117471 206352
rect 90909 206347 90975 206350
rect 114553 206347 114619 206350
rect 117405 206347 117471 206350
rect 83089 206274 83155 206277
rect 109309 206274 109375 206277
rect 121453 206274 121519 206277
rect 122790 206274 122850 206758
rect 259494 206756 259500 206758
rect 259564 206756 259570 206820
rect 83089 206272 122850 206274
rect 83089 206216 83094 206272
rect 83150 206216 109314 206272
rect 109370 206216 121458 206272
rect 121514 206216 122850 206272
rect 83089 206214 122850 206216
rect 83089 206211 83155 206214
rect 109309 206211 109375 206214
rect 121453 206211 121519 206214
rect 582465 205730 582531 205733
rect 583520 205730 584960 205820
rect 582465 205728 584960 205730
rect 582465 205672 582470 205728
rect 582526 205672 584960 205728
rect 582465 205670 584960 205672
rect 582465 205667 582531 205670
rect 57697 205594 57763 205597
rect 270677 205594 270743 205597
rect 57697 205592 270743 205594
rect 57697 205536 57702 205592
rect 57758 205536 270682 205592
rect 270738 205536 270743 205592
rect 583520 205580 584960 205670
rect 57697 205534 270743 205536
rect 57697 205531 57763 205534
rect 270677 205531 270743 205534
rect 97349 204914 97415 204917
rect 99373 204914 99439 204917
rect 97349 204912 99439 204914
rect 97349 204856 97354 204912
rect 97410 204856 99378 204912
rect 99434 204856 99439 204912
rect 97349 204854 99439 204856
rect 97349 204851 97415 204854
rect 99373 204851 99439 204854
rect 92974 204172 92980 204236
rect 93044 204234 93050 204236
rect 93710 204234 93716 204236
rect 93044 204174 93716 204234
rect 93044 204172 93050 204174
rect 93710 204172 93716 204174
rect 93780 204234 93786 204236
rect 250529 204234 250595 204237
rect 93780 204232 250595 204234
rect 93780 204176 250534 204232
rect 250590 204176 250595 204232
rect 93780 204174 250595 204176
rect 93780 204172 93786 204174
rect 250529 204171 250595 204174
rect 213177 202874 213243 202877
rect 218646 202874 218652 202876
rect 213177 202872 218652 202874
rect 213177 202816 213182 202872
rect 213238 202816 218652 202872
rect 213177 202814 218652 202816
rect 213177 202811 213243 202814
rect 218646 202812 218652 202814
rect 218716 202812 218722 202876
rect 88190 202132 88196 202196
rect 88260 202194 88266 202196
rect 103830 202194 103836 202196
rect 88260 202134 103836 202194
rect 88260 202132 88266 202134
rect 103830 202132 103836 202134
rect 103900 202132 103906 202196
rect -960 201922 480 202012
rect 3233 201922 3299 201925
rect -960 201920 3299 201922
rect -960 201864 3238 201920
rect 3294 201864 3299 201920
rect -960 201862 3299 201864
rect -960 201772 480 201862
rect 3233 201859 3299 201862
rect 92749 200698 92815 200701
rect 109534 200698 109540 200700
rect 92749 200696 109540 200698
rect 92749 200640 92754 200696
rect 92810 200640 109540 200696
rect 92749 200638 109540 200640
rect 92749 200635 92815 200638
rect 109534 200636 109540 200638
rect 109604 200636 109610 200700
rect 195237 200698 195303 200701
rect 205582 200698 205588 200700
rect 195237 200696 205588 200698
rect 195237 200640 195242 200696
rect 195298 200640 205588 200696
rect 195237 200638 205588 200640
rect 195237 200635 195303 200638
rect 205582 200636 205588 200638
rect 205652 200636 205658 200700
rect 206277 200698 206343 200701
rect 230974 200698 230980 200700
rect 206277 200696 230980 200698
rect 206277 200640 206282 200696
rect 206338 200640 230980 200696
rect 206277 200638 230980 200640
rect 206277 200635 206343 200638
rect 230974 200636 230980 200638
rect 231044 200636 231050 200700
rect 238661 200154 238727 200157
rect 238886 200154 238892 200156
rect 238616 200152 238892 200154
rect 238616 200096 238666 200152
rect 238722 200096 238892 200152
rect 238616 200094 238892 200096
rect 238661 200091 238727 200094
rect 238886 200092 238892 200094
rect 238956 200092 238962 200156
rect 102726 199956 102732 200020
rect 102796 200018 102802 200020
rect 102869 200018 102935 200021
rect 254526 200018 254532 200020
rect 102796 200016 254532 200018
rect 102796 199960 102874 200016
rect 102930 199960 254532 200016
rect 102796 199958 254532 199960
rect 102796 199956 102802 199958
rect 102869 199955 102935 199958
rect 254526 199956 254532 199958
rect 254596 199956 254602 200020
rect 238661 199882 238727 199885
rect 238886 199882 238892 199884
rect 238616 199880 238892 199882
rect 238616 199824 238666 199880
rect 238722 199824 238892 199880
rect 238616 199822 238892 199824
rect 238661 199819 238727 199822
rect 238886 199820 238892 199822
rect 238956 199820 238962 199884
rect 67950 192476 67956 192540
rect 68020 192538 68026 192540
rect 136633 192538 136699 192541
rect 68020 192536 136699 192538
rect 68020 192480 136638 192536
rect 136694 192480 136699 192536
rect 68020 192478 136699 192480
rect 68020 192476 68026 192478
rect 136633 192475 136699 192478
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 238661 190500 238727 190501
rect 238661 190498 238708 190500
rect 238616 190496 238708 190498
rect 238772 190498 238778 190500
rect 238616 190440 238666 190496
rect 238616 190438 238708 190440
rect 238661 190436 238708 190438
rect 238772 190438 238854 190498
rect 238772 190436 238778 190438
rect 238661 190435 238727 190436
rect 238661 190362 238727 190365
rect 238616 190360 238770 190362
rect 238616 190304 238666 190360
rect 238722 190304 238770 190360
rect 238616 190302 238770 190304
rect 238661 190299 238770 190302
rect 238710 190228 238770 190299
rect 238702 190164 238708 190228
rect 238772 190164 238778 190228
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 5441 188322 5507 188325
rect 219566 188322 219572 188324
rect 5441 188320 219572 188322
rect 5441 188264 5446 188320
rect 5502 188264 219572 188320
rect 5441 188262 219572 188264
rect 5441 188259 5507 188262
rect 219566 188260 219572 188262
rect 219636 188260 219642 188324
rect 111701 186962 111767 186965
rect 213678 186962 213684 186964
rect 111701 186960 213684 186962
rect 111701 186904 111706 186960
rect 111762 186904 213684 186960
rect 111701 186902 213684 186904
rect 111701 186899 111767 186902
rect 213678 186900 213684 186902
rect 213748 186900 213754 186964
rect 21357 185602 21423 185605
rect 198774 185602 198780 185604
rect 21357 185600 198780 185602
rect 21357 185544 21362 185600
rect 21418 185544 198780 185600
rect 21357 185542 198780 185544
rect 21357 185539 21423 185542
rect 198774 185540 198780 185542
rect 198844 185540 198850 185604
rect 238661 180844 238727 180845
rect 238661 180842 238708 180844
rect 238616 180840 238708 180842
rect 238772 180842 238778 180844
rect 238616 180784 238666 180840
rect 238616 180782 238708 180784
rect 238661 180780 238708 180782
rect 238772 180782 238854 180842
rect 238772 180780 238778 180782
rect 238661 180779 238727 180780
rect 238661 180706 238727 180709
rect 238616 180704 238770 180706
rect 238616 180648 238666 180704
rect 238722 180648 238770 180704
rect 238616 180646 238770 180648
rect 238661 180643 238770 180646
rect 238710 180572 238770 180643
rect 238702 180508 238708 180572
rect 238772 180508 238778 180572
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 238661 171188 238727 171189
rect 238661 171186 238708 171188
rect 238616 171184 238708 171186
rect 238772 171186 238778 171188
rect 238616 171128 238666 171184
rect 238616 171126 238708 171128
rect 238661 171124 238708 171126
rect 238772 171126 238854 171186
rect 238772 171124 238778 171126
rect 238661 171123 238727 171124
rect 238661 171052 238727 171053
rect 238661 171050 238708 171052
rect 238616 171048 238708 171050
rect 238772 171050 238778 171052
rect 238616 170992 238666 171048
rect 238616 170990 238708 170992
rect 238661 170988 238708 170990
rect 238772 170990 238854 171050
rect 238772 170988 238778 170990
rect 238661 170987 238727 170988
rect 580349 165882 580415 165885
rect 583520 165882 584960 165972
rect 580349 165880 584960 165882
rect 580349 165824 580354 165880
rect 580410 165824 584960 165880
rect 580349 165822 584960 165824
rect 580349 165819 580415 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 238661 161530 238727 161533
rect 238886 161530 238892 161532
rect 238616 161528 238892 161530
rect 238616 161472 238666 161528
rect 238722 161472 238892 161528
rect 238616 161470 238892 161472
rect 238661 161467 238727 161470
rect 238886 161468 238892 161470
rect 238956 161468 238962 161532
rect 238661 161394 238727 161397
rect 238616 161392 238770 161394
rect 238616 161336 238666 161392
rect 238722 161336 238770 161392
rect 238616 161334 238770 161336
rect 238661 161331 238770 161334
rect 238710 161260 238770 161331
rect 238702 161196 238708 161260
rect 238772 161196 238778 161260
rect 40677 153778 40743 153781
rect 203006 153778 203012 153780
rect 40677 153776 203012 153778
rect 40677 153720 40682 153776
rect 40738 153720 203012 153776
rect 40677 153718 203012 153720
rect 40677 153715 40743 153718
rect 203006 153716 203012 153718
rect 203076 153716 203082 153780
rect 583385 152690 583451 152693
rect 583520 152690 584960 152780
rect 583385 152688 584960 152690
rect 583385 152632 583390 152688
rect 583446 152632 584960 152688
rect 583385 152630 584960 152632
rect 583385 152627 583451 152630
rect 583520 152540 584960 152630
rect 238661 151876 238727 151877
rect 238661 151874 238708 151876
rect 238616 151872 238708 151874
rect 238772 151874 238778 151876
rect 238616 151816 238666 151872
rect 238616 151814 238708 151816
rect 238661 151812 238708 151814
rect 238772 151814 238854 151874
rect 238772 151812 238778 151814
rect 238661 151811 238727 151812
rect 238661 151738 238727 151741
rect 238616 151736 238770 151738
rect 238616 151680 238666 151736
rect 238722 151680 238770 151736
rect 238616 151678 238770 151680
rect 238661 151675 238770 151678
rect 238710 151604 238770 151675
rect 238702 151540 238708 151604
rect 238772 151540 238778 151604
rect 16389 151058 16455 151061
rect 197486 151058 197492 151060
rect 16389 151056 197492 151058
rect 16389 151000 16394 151056
rect 16450 151000 197492 151056
rect 16389 150998 197492 151000
rect 16389 150995 16455 150998
rect 197486 150996 197492 150998
rect 197556 150996 197562 151060
rect -960 149834 480 149924
rect 2957 149834 3023 149837
rect -960 149832 3023 149834
rect -960 149776 2962 149832
rect 3018 149776 3023 149832
rect -960 149774 3023 149776
rect -960 149684 480 149774
rect 2957 149771 3023 149774
rect 50337 149698 50403 149701
rect 191046 149698 191052 149700
rect 50337 149696 191052 149698
rect 50337 149640 50342 149696
rect 50398 149640 191052 149696
rect 50337 149638 191052 149640
rect 50337 149635 50403 149638
rect 191046 149636 191052 149638
rect 191116 149636 191122 149700
rect 92473 148338 92539 148341
rect 122598 148338 122604 148340
rect 92473 148336 122604 148338
rect 92473 148280 92478 148336
rect 92534 148280 122604 148336
rect 92473 148278 122604 148280
rect 92473 148275 92539 148278
rect 122598 148276 122604 148278
rect 122668 148276 122674 148340
rect 48221 146978 48287 146981
rect 223798 146978 223804 146980
rect 48221 146976 223804 146978
rect 48221 146920 48226 146976
rect 48282 146920 223804 146976
rect 48221 146918 223804 146920
rect 48221 146915 48287 146918
rect 223798 146916 223804 146918
rect 223868 146916 223874 146980
rect 66161 145618 66227 145621
rect 238661 145618 238727 145621
rect 239254 145618 239260 145620
rect 66161 145616 239260 145618
rect 66161 145560 66166 145616
rect 66222 145560 238666 145616
rect 238722 145560 239260 145616
rect 66161 145558 239260 145560
rect 66161 145555 66227 145558
rect 238661 145555 238727 145558
rect 239254 145556 239260 145558
rect 239324 145556 239330 145620
rect 84469 141402 84535 141405
rect 121637 141402 121703 141405
rect 295333 141402 295399 141405
rect 84469 141400 295399 141402
rect 84469 141344 84474 141400
rect 84530 141344 121642 141400
rect 121698 141344 295338 141400
rect 295394 141344 295399 141400
rect 84469 141342 295399 141344
rect 84469 141339 84535 141342
rect 121637 141339 121703 141342
rect 295333 141339 295399 141342
rect 68553 140858 68619 140861
rect 71957 140858 72023 140861
rect 68553 140856 72023 140858
rect 68553 140800 68558 140856
rect 68614 140800 71962 140856
rect 72018 140800 72023 140856
rect 68553 140798 72023 140800
rect 68553 140795 68619 140798
rect 71957 140795 72023 140798
rect 88793 140042 88859 140045
rect 125593 140042 125659 140045
rect 88793 140040 125659 140042
rect 88793 139984 88798 140040
rect 88854 139984 125598 140040
rect 125654 139984 125659 140040
rect 88793 139982 125659 139984
rect 88793 139979 88859 139982
rect 125593 139979 125659 139982
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 81065 138682 81131 138685
rect 117313 138682 117379 138685
rect 81065 138680 117379 138682
rect 81065 138624 81070 138680
rect 81126 138624 117318 138680
rect 117374 138624 117379 138680
rect 81065 138622 117379 138624
rect 81065 138619 81131 138622
rect 117313 138619 117379 138622
rect 239254 138620 239260 138684
rect 239324 138682 239330 138684
rect 249057 138682 249123 138685
rect 239324 138680 249123 138682
rect 239324 138624 249062 138680
rect 249118 138624 249123 138680
rect 239324 138622 249123 138624
rect 239324 138620 239330 138622
rect 249057 138619 249123 138622
rect 68870 138076 68876 138140
rect 68940 138138 68946 138140
rect 72141 138138 72207 138141
rect 68940 138136 72207 138138
rect 68940 138080 72146 138136
rect 72202 138080 72207 138136
rect 68940 138078 72207 138080
rect 68940 138076 68946 138078
rect 72141 138075 72207 138078
rect 80421 137458 80487 137461
rect 94957 137458 95023 137461
rect 80421 137456 95023 137458
rect 80421 137400 80426 137456
rect 80482 137400 94962 137456
rect 95018 137400 95023 137456
rect 80421 137398 95023 137400
rect 80421 137395 80487 137398
rect 94957 137395 95023 137398
rect 52085 137322 52151 137325
rect 73797 137322 73863 137325
rect 52085 137320 73863 137322
rect 52085 137264 52090 137320
rect 52146 137264 73802 137320
rect 73858 137264 73863 137320
rect 52085 137262 73863 137264
rect 52085 137259 52151 137262
rect 73797 137259 73863 137262
rect 86861 137322 86927 137325
rect 104157 137322 104223 137325
rect 86861 137320 104223 137322
rect 86861 137264 86866 137320
rect 86922 137264 104162 137320
rect 104218 137264 104223 137320
rect 86861 137262 104223 137264
rect 86861 137259 86927 137262
rect 104157 137259 104223 137262
rect 69841 136914 69907 136917
rect 71078 136914 71084 136916
rect 69841 136912 71084 136914
rect -960 136778 480 136868
rect 69841 136856 69846 136912
rect 69902 136856 71084 136912
rect 69841 136854 71084 136856
rect 69841 136851 69907 136854
rect 71078 136852 71084 136854
rect 71148 136852 71154 136916
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 87321 136778 87387 136781
rect 88190 136778 88196 136780
rect 87321 136776 88196 136778
rect 87321 136720 87326 136776
rect 87382 136720 88196 136776
rect 87321 136718 88196 136720
rect 87321 136715 87387 136718
rect 88190 136716 88196 136718
rect 88260 136716 88266 136780
rect 63309 135962 63375 135965
rect 73245 135962 73311 135965
rect 63309 135960 73311 135962
rect 63309 135904 63314 135960
rect 63370 135904 73250 135960
rect 73306 135904 73311 135960
rect 63309 135902 73311 135904
rect 63309 135899 63375 135902
rect 73245 135899 73311 135902
rect 92381 135282 92447 135285
rect 94078 135282 94084 135284
rect 92381 135280 94084 135282
rect 92381 135224 92386 135280
rect 92442 135224 94084 135280
rect 92381 135222 94084 135224
rect 92381 135219 92447 135222
rect 94078 135220 94084 135222
rect 94148 135220 94154 135284
rect 71681 134740 71747 134741
rect 71630 134738 71636 134740
rect 71590 134678 71636 134738
rect 71700 134736 71747 134740
rect 71742 134680 71747 134736
rect 71630 134676 71636 134678
rect 71700 134676 71747 134680
rect 71681 134675 71747 134676
rect 94865 134602 94931 134605
rect 100753 134602 100819 134605
rect 94865 134600 100819 134602
rect 94865 134544 94870 134600
rect 94926 134544 100758 134600
rect 100814 134544 100819 134600
rect 94865 134542 100819 134544
rect 94865 134539 94931 134542
rect 100753 134539 100819 134542
rect 66253 134466 66319 134469
rect 66253 134464 68908 134466
rect 66253 134408 66258 134464
rect 66314 134408 68908 134464
rect 66253 134406 68908 134408
rect 66253 134403 66319 134406
rect 97441 133922 97507 133925
rect 94668 133920 97507 133922
rect 94668 133864 97446 133920
rect 97502 133864 97507 133920
rect 94668 133862 97507 133864
rect 97441 133859 97507 133862
rect 66253 133650 66319 133653
rect 66253 133648 68908 133650
rect 66253 133592 66258 133648
rect 66314 133592 68908 133648
rect 66253 133590 68908 133592
rect 66253 133587 66319 133590
rect 96705 133106 96771 133109
rect 94668 133104 96771 133106
rect 94668 133048 96710 133104
rect 96766 133048 96771 133104
rect 94668 133046 96771 133048
rect 96705 133043 96771 133046
rect 67766 132772 67772 132836
rect 67836 132834 67842 132836
rect 67836 132774 68908 132834
rect 67836 132772 67842 132774
rect 96613 132290 96679 132293
rect 94668 132288 96679 132290
rect 94668 132232 96618 132288
rect 96674 132232 96679 132288
rect 94668 132230 96679 132232
rect 96613 132227 96679 132230
rect 66253 132018 66319 132021
rect 66253 132016 68908 132018
rect 66253 131960 66258 132016
rect 66314 131960 68908 132016
rect 66253 131958 68908 131960
rect 66253 131955 66319 131958
rect 97349 131474 97415 131477
rect 94668 131472 97415 131474
rect 94668 131416 97354 131472
rect 97410 131416 97415 131472
rect 94668 131414 97415 131416
rect 97349 131411 97415 131414
rect 66345 131202 66411 131205
rect 66345 131200 68908 131202
rect 66345 131144 66350 131200
rect 66406 131144 68908 131200
rect 66345 131142 68908 131144
rect 66345 131139 66411 131142
rect 97257 130930 97323 130933
rect 94668 130928 97323 130930
rect 94668 130872 97262 130928
rect 97318 130872 97323 130928
rect 94668 130870 97323 130872
rect 97257 130867 97323 130870
rect 62982 130596 62988 130660
rect 63052 130658 63058 130660
rect 63052 130598 68908 130658
rect 63052 130596 63058 130598
rect 94638 129978 94698 130084
rect 106774 129978 106780 129980
rect 94638 129918 106780 129978
rect 106774 129916 106780 129918
rect 106844 129916 106850 129980
rect 67541 129842 67607 129845
rect 67541 129840 68908 129842
rect 67541 129784 67546 129840
rect 67602 129784 68908 129840
rect 67541 129782 68908 129784
rect 67541 129779 67607 129782
rect 96705 129298 96771 129301
rect 94668 129296 96771 129298
rect 94668 129240 96710 129296
rect 96766 129240 96771 129296
rect 94668 129238 96771 129240
rect 96705 129235 96771 129238
rect 65977 129026 66043 129029
rect 65977 129024 68908 129026
rect 65977 128968 65982 129024
rect 66038 128968 68908 129024
rect 65977 128966 68908 128968
rect 65977 128963 66043 128966
rect 102869 128482 102935 128485
rect 94668 128480 102935 128482
rect 94668 128424 102874 128480
rect 102930 128424 102935 128480
rect 94668 128422 102935 128424
rect 102869 128419 102935 128422
rect 66437 128210 66503 128213
rect 66437 128208 68908 128210
rect 66437 128152 66442 128208
rect 66498 128152 68908 128208
rect 66437 128150 68908 128152
rect 66437 128147 66503 128150
rect 66897 127666 66963 127669
rect 97165 127666 97231 127669
rect 66897 127664 68908 127666
rect 66897 127608 66902 127664
rect 66958 127608 68908 127664
rect 66897 127606 68908 127608
rect 94668 127664 97231 127666
rect 94668 127608 97170 127664
rect 97226 127608 97231 127664
rect 94668 127606 97231 127608
rect 66897 127603 66963 127606
rect 97165 127603 97231 127606
rect 97533 127122 97599 127125
rect 94668 127120 97599 127122
rect 94668 127064 97538 127120
rect 97594 127064 97599 127120
rect 94668 127062 97599 127064
rect 97533 127059 97599 127062
rect 66713 126850 66779 126853
rect 66713 126848 68908 126850
rect 66713 126792 66718 126848
rect 66774 126792 68908 126848
rect 66713 126790 68908 126792
rect 66713 126787 66779 126790
rect 97809 126306 97875 126309
rect 94668 126304 97875 126306
rect 94668 126248 97814 126304
rect 97870 126248 97875 126304
rect 94668 126246 97875 126248
rect 97809 126243 97875 126246
rect 66069 126034 66135 126037
rect 583293 126034 583359 126037
rect 583520 126034 584960 126124
rect 66069 126032 68908 126034
rect 66069 125976 66074 126032
rect 66130 125976 68908 126032
rect 66069 125974 68908 125976
rect 583293 126032 584960 126034
rect 583293 125976 583298 126032
rect 583354 125976 584960 126032
rect 583293 125974 584960 125976
rect 66069 125971 66135 125974
rect 583293 125971 583359 125974
rect 583520 125884 584960 125974
rect 96797 125490 96863 125493
rect 94668 125488 96863 125490
rect 94668 125432 96802 125488
rect 96858 125432 96863 125488
rect 94668 125430 96863 125432
rect 96797 125427 96863 125430
rect 66897 125218 66963 125221
rect 66897 125216 68908 125218
rect 66897 125160 66902 125216
rect 66958 125160 68908 125216
rect 66897 125158 68908 125160
rect 66897 125155 66963 125158
rect 104157 124810 104223 124813
rect 318793 124810 318859 124813
rect 104157 124808 318859 124810
rect 104157 124752 104162 124808
rect 104218 124752 318798 124808
rect 318854 124752 318859 124808
rect 104157 124750 318859 124752
rect 104157 124747 104223 124750
rect 318793 124747 318859 124750
rect 97441 124674 97507 124677
rect 94668 124672 97507 124674
rect 94668 124616 97446 124672
rect 97502 124616 97507 124672
rect 94668 124614 97507 124616
rect 97441 124611 97507 124614
rect 66253 124402 66319 124405
rect 66253 124400 68908 124402
rect 66253 124344 66258 124400
rect 66314 124344 68908 124400
rect 66253 124342 68908 124344
rect 66253 124339 66319 124342
rect 95233 124132 95299 124133
rect 95182 124130 95188 124132
rect 94638 123994 94698 124100
rect 95142 124070 95188 124130
rect 95252 124128 95299 124132
rect 95294 124072 95299 124128
rect 95182 124068 95188 124070
rect 95252 124068 95299 124072
rect 95233 124067 95299 124068
rect 96613 123994 96679 123997
rect 94638 123992 96679 123994
rect 94638 123936 96618 123992
rect 96674 123936 96679 123992
rect 94638 123934 96679 123936
rect 96613 123931 96679 123934
rect 65517 123858 65583 123861
rect 65517 123856 68908 123858
rect -960 123572 480 123812
rect 65517 123800 65522 123856
rect 65578 123800 68908 123856
rect 65517 123798 68908 123800
rect 65517 123795 65583 123798
rect 97809 123314 97875 123317
rect 94668 123312 97875 123314
rect 94668 123256 97814 123312
rect 97870 123256 97875 123312
rect 94668 123254 97875 123256
rect 97809 123251 97875 123254
rect 66897 123042 66963 123045
rect 66897 123040 68908 123042
rect 66897 122984 66902 123040
rect 66958 122984 68908 123040
rect 66897 122982 68908 122984
rect 66897 122979 66963 122982
rect 97809 122498 97875 122501
rect 94668 122496 97875 122498
rect 94668 122440 97814 122496
rect 97870 122440 97875 122496
rect 94668 122438 97875 122440
rect 97809 122435 97875 122438
rect 66897 122226 66963 122229
rect 66897 122224 68908 122226
rect 66897 122168 66902 122224
rect 66958 122168 68908 122224
rect 66897 122166 68908 122168
rect 66897 122163 66963 122166
rect 94638 121546 94698 121652
rect 120257 121546 120323 121549
rect 94638 121544 120323 121546
rect 94638 121488 120262 121544
rect 120318 121488 120323 121544
rect 94638 121486 120323 121488
rect 120257 121483 120323 121486
rect 68878 120866 68938 121380
rect 97809 120866 97875 120869
rect 64830 120806 68938 120866
rect 94668 120864 97875 120866
rect 94668 120808 97814 120864
rect 97870 120808 97875 120864
rect 94668 120806 97875 120808
rect 63125 120186 63191 120189
rect 64830 120186 64890 120806
rect 97809 120803 97875 120806
rect 66713 120594 66779 120597
rect 66713 120592 68908 120594
rect 66713 120536 66718 120592
rect 66774 120536 68908 120592
rect 66713 120534 68908 120536
rect 66713 120531 66779 120534
rect 97809 120322 97875 120325
rect 94668 120320 97875 120322
rect 94668 120264 97814 120320
rect 97870 120264 97875 120320
rect 94668 120262 97875 120264
rect 97809 120259 97875 120262
rect 63125 120184 64890 120186
rect 63125 120128 63130 120184
rect 63186 120128 64890 120184
rect 63125 120126 64890 120128
rect 63125 120123 63191 120126
rect 66897 120050 66963 120053
rect 66897 120048 68908 120050
rect 66897 119992 66902 120048
rect 66958 119992 68908 120048
rect 66897 119990 68908 119992
rect 66897 119987 66963 119990
rect 66069 119234 66135 119237
rect 66253 119234 66319 119237
rect 66069 119232 68908 119234
rect 66069 119176 66074 119232
rect 66130 119176 66258 119232
rect 66314 119176 68908 119232
rect 66069 119174 68908 119176
rect 66069 119171 66135 119174
rect 66253 119171 66319 119174
rect 94638 118962 94698 119476
rect 118734 118962 118740 118964
rect 94638 118902 118740 118962
rect 118734 118900 118740 118902
rect 118804 118900 118810 118964
rect 98494 118690 98500 118692
rect 94668 118630 98500 118690
rect 98494 118628 98500 118630
rect 98564 118628 98570 118692
rect 66897 118418 66963 118421
rect 66897 118416 68908 118418
rect 66897 118360 66902 118416
rect 66958 118360 68908 118416
rect 66897 118358 68908 118360
rect 66897 118355 66963 118358
rect 97809 117874 97875 117877
rect 94668 117872 97875 117874
rect 94668 117816 97814 117872
rect 97870 117816 97875 117872
rect 94668 117814 97875 117816
rect 97809 117811 97875 117814
rect 66161 117602 66227 117605
rect 66161 117600 68908 117602
rect 66161 117544 66166 117600
rect 66222 117544 68908 117600
rect 66161 117542 68908 117544
rect 66161 117539 66227 117542
rect 66897 117058 66963 117061
rect 96613 117058 96679 117061
rect 66897 117056 68908 117058
rect 66897 117000 66902 117056
rect 66958 117000 68908 117056
rect 66897 116998 68908 117000
rect 94668 117056 96679 117058
rect 94668 117000 96618 117056
rect 96674 117000 96679 117056
rect 94668 116998 96679 117000
rect 66897 116995 66963 116998
rect 96613 116995 96679 116998
rect 97809 116514 97875 116517
rect 94668 116512 97875 116514
rect 94668 116456 97814 116512
rect 97870 116456 97875 116512
rect 94668 116454 97875 116456
rect 97809 116451 97875 116454
rect 64638 116044 64644 116108
rect 64708 116106 64714 116108
rect 68878 116106 68938 116212
rect 64708 116046 68938 116106
rect 64708 116044 64714 116046
rect 97809 115698 97875 115701
rect 94668 115696 97875 115698
rect 94668 115640 97814 115696
rect 97870 115640 97875 115696
rect 94668 115638 97875 115640
rect 97809 115635 97875 115638
rect 66897 115426 66963 115429
rect 66897 115424 68908 115426
rect 66897 115368 66902 115424
rect 66958 115368 68908 115424
rect 66897 115366 68908 115368
rect 66897 115363 66963 115366
rect 98637 115154 98703 115157
rect 114502 115154 114508 115156
rect 98637 115152 114508 115154
rect 98637 115096 98642 115152
rect 98698 115096 114508 115152
rect 98637 115094 114508 115096
rect 98637 115091 98703 115094
rect 114502 115092 114508 115094
rect 114572 115092 114578 115156
rect 97717 114882 97783 114885
rect 94668 114880 97783 114882
rect 94668 114824 97722 114880
rect 97778 114824 97783 114880
rect 94668 114822 97783 114824
rect 97717 114819 97783 114822
rect 67173 114610 67239 114613
rect 67173 114608 68908 114610
rect 67173 114552 67178 114608
rect 67234 114552 68908 114608
rect 67173 114550 68908 114552
rect 67173 114547 67239 114550
rect 96613 114066 96679 114069
rect 94668 114064 96679 114066
rect 94668 114008 96618 114064
rect 96674 114008 96679 114064
rect 94668 114006 96679 114008
rect 96613 114003 96679 114006
rect 68878 113522 68938 113764
rect 64830 113462 68938 113522
rect 64597 113250 64663 113253
rect 64830 113250 64890 113462
rect 94638 113386 94698 113492
rect 133873 113386 133939 113389
rect 94638 113384 133939 113386
rect 94638 113328 133878 113384
rect 133934 113328 133939 113384
rect 94638 113326 133939 113328
rect 133873 113323 133939 113326
rect 64597 113248 64890 113250
rect 64597 113192 64602 113248
rect 64658 113192 64890 113248
rect 64597 113190 64890 113192
rect 66621 113250 66687 113253
rect 66621 113248 68908 113250
rect 66621 113192 66626 113248
rect 66682 113192 68908 113248
rect 66621 113190 68908 113192
rect 64597 113187 64663 113190
rect 66621 113187 66687 113190
rect 61878 113052 61884 113116
rect 61948 113114 61954 113116
rect 66846 113114 66852 113116
rect 61948 113054 66852 113114
rect 61948 113052 61954 113054
rect 66846 113052 66852 113054
rect 66916 113052 66922 113116
rect 583109 112842 583175 112845
rect 583520 112842 584960 112932
rect 583109 112840 584960 112842
rect 583109 112784 583114 112840
rect 583170 112784 584960 112840
rect 583109 112782 584960 112784
rect 583109 112779 583175 112782
rect 97809 112706 97875 112709
rect 94668 112704 97875 112706
rect 94668 112648 97814 112704
rect 97870 112648 97875 112704
rect 583520 112692 584960 112782
rect 94668 112646 97875 112648
rect 97809 112643 97875 112646
rect 66897 112434 66963 112437
rect 66897 112432 68908 112434
rect 66897 112376 66902 112432
rect 66958 112376 68908 112432
rect 66897 112374 68908 112376
rect 66897 112371 66963 112374
rect 95969 111890 96035 111893
rect 94668 111888 96035 111890
rect 94668 111832 95974 111888
rect 96030 111832 96035 111888
rect 94668 111830 96035 111832
rect 95969 111827 96035 111830
rect 66846 111556 66852 111620
rect 66916 111618 66922 111620
rect 66916 111558 68908 111618
rect 66916 111556 66922 111558
rect 97901 111074 97967 111077
rect 94668 111072 97967 111074
rect 94668 111016 97906 111072
rect 97962 111016 97967 111072
rect 94668 111014 97967 111016
rect 97901 111011 97967 111014
rect 98729 111074 98795 111077
rect 116761 111074 116827 111077
rect 98729 111072 116827 111074
rect 98729 111016 98734 111072
rect 98790 111016 116766 111072
rect 116822 111016 116827 111072
rect 98729 111014 116827 111016
rect 98729 111011 98795 111014
rect 116761 111011 116827 111014
rect 66897 110802 66963 110805
rect 66897 110800 68908 110802
rect -960 110666 480 110756
rect 66897 110744 66902 110800
rect 66958 110744 68908 110800
rect 66897 110742 68908 110744
rect 66897 110739 66963 110742
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 66253 110258 66319 110261
rect 97901 110258 97967 110261
rect 66253 110256 68908 110258
rect 66253 110200 66258 110256
rect 66314 110200 68908 110256
rect 66253 110198 68908 110200
rect 94668 110256 97967 110258
rect 94668 110200 97906 110256
rect 97962 110200 97967 110256
rect 94668 110198 97967 110200
rect 66253 110195 66319 110198
rect 97901 110195 97967 110198
rect 97809 109714 97875 109717
rect 94668 109712 97875 109714
rect 94668 109656 97814 109712
rect 97870 109656 97875 109712
rect 94668 109654 97875 109656
rect 97809 109651 97875 109654
rect 66897 109442 66963 109445
rect 66897 109440 68908 109442
rect 66897 109384 66902 109440
rect 66958 109384 68908 109440
rect 66897 109382 68908 109384
rect 66897 109379 66963 109382
rect 97901 108898 97967 108901
rect 94668 108896 97967 108898
rect 94668 108840 97906 108896
rect 97962 108840 97967 108896
rect 94668 108838 97967 108840
rect 97901 108835 97967 108838
rect 66897 108626 66963 108629
rect 66897 108624 68908 108626
rect 66897 108568 66902 108624
rect 66958 108568 68908 108624
rect 66897 108566 68908 108568
rect 66897 108563 66963 108566
rect 97206 108292 97212 108356
rect 97276 108354 97282 108356
rect 128997 108354 129063 108357
rect 97276 108352 129063 108354
rect 97276 108296 129002 108352
rect 129058 108296 129063 108352
rect 97276 108294 129063 108296
rect 97276 108292 97282 108294
rect 128997 108291 129063 108294
rect 97717 108082 97783 108085
rect 94668 108080 97783 108082
rect 94668 108024 97722 108080
rect 97778 108024 97783 108080
rect 94668 108022 97783 108024
rect 97717 108019 97783 108022
rect 66989 107810 67055 107813
rect 66989 107808 68908 107810
rect 66989 107752 66994 107808
rect 67050 107752 68908 107808
rect 66989 107750 68908 107752
rect 66989 107747 67055 107750
rect 66897 106994 66963 106997
rect 94638 106994 94698 107236
rect 66897 106992 68908 106994
rect 66897 106936 66902 106992
rect 66958 106936 68908 106992
rect 66897 106934 68908 106936
rect 94638 106934 103530 106994
rect 66897 106931 66963 106934
rect 97533 106722 97599 106725
rect 94668 106720 97599 106722
rect 94668 106664 97538 106720
rect 97594 106664 97599 106720
rect 94668 106662 97599 106664
rect 97533 106659 97599 106662
rect 66713 106450 66779 106453
rect 66713 106448 68908 106450
rect 66713 106392 66718 106448
rect 66774 106392 68908 106448
rect 66713 106390 68908 106392
rect 66713 106387 66779 106390
rect 103470 106314 103530 106934
rect 124438 106314 124444 106316
rect 103470 106254 124444 106314
rect 124438 106252 124444 106254
rect 124508 106252 124514 106316
rect 97901 105906 97967 105909
rect 94668 105904 97967 105906
rect 94668 105848 97906 105904
rect 97962 105848 97967 105904
rect 94668 105846 97967 105848
rect 97901 105843 97967 105846
rect 66897 105634 66963 105637
rect 66897 105632 68908 105634
rect 66897 105576 66902 105632
rect 66958 105576 68908 105632
rect 66897 105574 68908 105576
rect 66897 105571 66963 105574
rect 97625 105090 97691 105093
rect 94668 105088 97691 105090
rect 94668 105032 97630 105088
rect 97686 105032 97691 105088
rect 94668 105030 97691 105032
rect 97625 105027 97691 105030
rect 66253 104818 66319 104821
rect 66253 104816 68908 104818
rect 66253 104760 66258 104816
rect 66314 104760 68908 104816
rect 66253 104758 68908 104760
rect 66253 104755 66319 104758
rect 97165 104274 97231 104277
rect 94668 104272 97231 104274
rect 94668 104216 97170 104272
rect 97226 104216 97231 104272
rect 94668 104214 97231 104216
rect 97165 104211 97231 104214
rect 102041 104138 102107 104141
rect 233366 104138 233372 104140
rect 102041 104136 233372 104138
rect 102041 104080 102046 104136
rect 102102 104080 233372 104136
rect 102041 104078 233372 104080
rect 102041 104075 102107 104078
rect 233366 104076 233372 104078
rect 233436 104076 233442 104140
rect 67357 104002 67423 104005
rect 67357 104000 68908 104002
rect 67357 103944 67362 104000
rect 67418 103944 68908 104000
rect 67357 103942 68908 103944
rect 67357 103939 67423 103942
rect 97206 103458 97212 103460
rect 94668 103398 97212 103458
rect 97206 103396 97212 103398
rect 97276 103396 97282 103460
rect 66897 103186 66963 103189
rect 66897 103184 68908 103186
rect 66897 103128 66902 103184
rect 66958 103128 68908 103184
rect 66897 103126 68908 103128
rect 66897 103123 66963 103126
rect 97165 102914 97231 102917
rect 94668 102912 97231 102914
rect 94668 102856 97170 102912
rect 97226 102856 97231 102912
rect 94668 102854 97231 102856
rect 97165 102851 97231 102854
rect 67541 102642 67607 102645
rect 67541 102640 68908 102642
rect 67541 102584 67546 102640
rect 67602 102584 68908 102640
rect 67541 102582 68908 102584
rect 67541 102579 67607 102582
rect 59118 102172 59124 102236
rect 59188 102234 59194 102236
rect 67541 102234 67607 102237
rect 59188 102232 67607 102234
rect 59188 102176 67546 102232
rect 67602 102176 67607 102232
rect 59188 102174 67607 102176
rect 59188 102172 59194 102174
rect 67541 102171 67607 102174
rect 97901 102098 97967 102101
rect 94668 102096 97967 102098
rect 94668 102040 97906 102096
rect 97962 102040 97967 102096
rect 94668 102038 97967 102040
rect 97901 102035 97967 102038
rect 66805 101826 66871 101829
rect 66805 101824 68908 101826
rect 66805 101768 66810 101824
rect 66866 101768 68908 101824
rect 66805 101766 68908 101768
rect 66805 101763 66871 101766
rect 95969 101418 96035 101421
rect 109309 101418 109375 101421
rect 95969 101416 109375 101418
rect 95969 101360 95974 101416
rect 96030 101360 109314 101416
rect 109370 101360 109375 101416
rect 95969 101358 109375 101360
rect 95969 101355 96035 101358
rect 109309 101355 109375 101358
rect 233141 101418 233207 101421
rect 238518 101418 238524 101420
rect 233141 101416 238524 101418
rect 233141 101360 233146 101416
rect 233202 101360 238524 101416
rect 233141 101358 238524 101360
rect 233141 101355 233207 101358
rect 238518 101356 238524 101358
rect 238588 101356 238594 101420
rect 97809 101282 97875 101285
rect 94668 101280 97875 101282
rect 94668 101224 97814 101280
rect 97870 101224 97875 101280
rect 94668 101222 97875 101224
rect 97809 101219 97875 101222
rect 66437 101010 66503 101013
rect 66437 101008 68908 101010
rect 66437 100952 66442 101008
rect 66498 100952 68908 101008
rect 66437 100950 68908 100952
rect 66437 100947 66503 100950
rect 97901 100466 97967 100469
rect 94668 100464 97967 100466
rect 94668 100408 97906 100464
rect 97962 100408 97967 100464
rect 94668 100406 97967 100408
rect 97901 100403 97967 100406
rect 66805 100194 66871 100197
rect 66805 100192 68908 100194
rect 66805 100136 66810 100192
rect 66866 100136 68908 100192
rect 66805 100134 68908 100136
rect 66805 100131 66871 100134
rect 97349 100058 97415 100061
rect 121678 100058 121684 100060
rect 97349 100056 121684 100058
rect 97349 100000 97354 100056
rect 97410 100000 121684 100056
rect 97349 99998 121684 100000
rect 97349 99995 97415 99998
rect 121678 99996 121684 99998
rect 121748 99996 121754 100060
rect 66805 99650 66871 99653
rect 97717 99650 97783 99653
rect 66805 99648 68908 99650
rect 66805 99592 66810 99648
rect 66866 99592 68908 99648
rect 66805 99590 68908 99592
rect 94668 99648 97783 99650
rect 94668 99592 97722 99648
rect 97778 99592 97783 99648
rect 94668 99590 97783 99592
rect 66805 99587 66871 99590
rect 97717 99587 97783 99590
rect 583201 99514 583267 99517
rect 583520 99514 584960 99604
rect 583201 99512 584960 99514
rect 583201 99456 583206 99512
rect 583262 99456 584960 99512
rect 583201 99454 584960 99456
rect 583201 99451 583267 99454
rect 583520 99364 584960 99454
rect 66805 98834 66871 98837
rect 66805 98832 68908 98834
rect 66805 98776 66810 98832
rect 66866 98776 68908 98832
rect 66805 98774 68908 98776
rect 66805 98771 66871 98774
rect 94638 98562 94698 99076
rect 108246 98562 108252 98564
rect 94638 98502 108252 98562
rect 108246 98500 108252 98502
rect 108316 98500 108322 98564
rect 97533 98290 97599 98293
rect 94668 98288 97599 98290
rect 94668 98232 97538 98288
rect 97594 98232 97599 98288
rect 94668 98230 97599 98232
rect 97533 98227 97599 98230
rect 67449 98018 67515 98021
rect 67449 98016 68908 98018
rect 67449 97960 67454 98016
rect 67510 97960 68908 98016
rect 67449 97958 68908 97960
rect 67449 97955 67515 97958
rect -960 97610 480 97700
rect 3049 97610 3115 97613
rect -960 97608 3115 97610
rect -960 97552 3054 97608
rect 3110 97552 3115 97608
rect -960 97550 3115 97552
rect -960 97460 480 97550
rect 3049 97547 3115 97550
rect 97901 97474 97967 97477
rect 94668 97472 97967 97474
rect 94668 97416 97906 97472
rect 97962 97416 97967 97472
rect 94668 97414 97967 97416
rect 97901 97411 97967 97414
rect 66897 97202 66963 97205
rect 66897 97200 68908 97202
rect 66897 97144 66902 97200
rect 66958 97144 68908 97200
rect 66897 97142 68908 97144
rect 66897 97139 66963 97142
rect 99046 97140 99052 97204
rect 99116 97202 99122 97204
rect 232078 97202 232084 97204
rect 99116 97142 232084 97202
rect 99116 97140 99122 97142
rect 232078 97140 232084 97142
rect 232148 97140 232154 97204
rect 97533 96658 97599 96661
rect 94668 96656 97599 96658
rect 94668 96600 97538 96656
rect 97594 96600 97599 96656
rect 94668 96598 97599 96600
rect 97533 96595 97599 96598
rect 66253 96386 66319 96389
rect 66253 96384 68908 96386
rect 66253 96328 66258 96384
rect 66314 96328 68908 96384
rect 66253 96326 68908 96328
rect 66253 96323 66319 96326
rect 66805 95842 66871 95845
rect 66805 95840 68908 95842
rect 66805 95784 66810 95840
rect 66866 95784 68908 95840
rect 66805 95782 68908 95784
rect 66805 95779 66871 95782
rect 94638 95570 94698 96084
rect 127249 95570 127315 95573
rect 94638 95568 127315 95570
rect 94638 95512 127254 95568
rect 127310 95512 127315 95568
rect 94638 95510 127315 95512
rect 127249 95507 127315 95510
rect 66110 95236 66116 95300
rect 66180 95298 66186 95300
rect 97901 95298 97967 95301
rect 66180 95238 66316 95298
rect 94668 95296 97967 95298
rect 94668 95240 97906 95296
rect 97962 95240 97967 95296
rect 94668 95238 97967 95240
rect 66180 95236 66186 95238
rect 66256 94890 66316 95238
rect 97901 95235 97967 95238
rect 66437 95026 66503 95029
rect 66437 95024 68908 95026
rect 66437 94968 66442 95024
rect 66498 94968 68908 95024
rect 66437 94966 68908 94968
rect 66437 94963 66503 94966
rect 66256 94830 68938 94890
rect 68878 94180 68938 94830
rect 97901 94482 97967 94485
rect 232262 94482 232268 94484
rect 94668 94480 97967 94482
rect 94668 94424 97906 94480
rect 97962 94424 97967 94480
rect 94668 94422 97967 94424
rect 97901 94419 97967 94422
rect 103470 94422 232268 94482
rect 95141 94346 95207 94349
rect 103470 94346 103530 94422
rect 232262 94420 232268 94422
rect 232332 94420 232338 94484
rect 95141 94344 103530 94346
rect 95141 94288 95146 94344
rect 95202 94288 103530 94344
rect 95141 94286 103530 94288
rect 95141 94283 95207 94286
rect 97901 93666 97967 93669
rect 94668 93664 97967 93666
rect 94668 93608 97906 93664
rect 97962 93608 97967 93664
rect 94668 93606 97967 93608
rect 97901 93603 97967 93606
rect 66805 93394 66871 93397
rect 66805 93392 69460 93394
rect 66805 93336 66810 93392
rect 66866 93364 69460 93392
rect 66866 93336 69490 93364
rect 66805 93334 69490 93336
rect 66805 93331 66871 93334
rect 69430 92714 69490 93334
rect 97349 92850 97415 92853
rect 94668 92848 97415 92850
rect 94668 92792 97354 92848
rect 97410 92792 97415 92848
rect 94668 92790 97415 92792
rect 97349 92787 97415 92790
rect 69565 92714 69631 92717
rect 69430 92712 69631 92714
rect 69430 92656 69570 92712
rect 69626 92656 69631 92712
rect 69430 92654 69631 92656
rect 69565 92651 69631 92654
rect 69703 92714 69769 92717
rect 69974 92714 69980 92716
rect 69703 92712 69980 92714
rect 69703 92656 69708 92712
rect 69764 92656 69980 92712
rect 69703 92654 69980 92656
rect 69703 92651 69769 92654
rect 69974 92652 69980 92654
rect 70044 92652 70050 92716
rect 70894 92714 70900 92716
rect 70856 92683 70900 92714
rect 70807 92678 70900 92683
rect 70807 92622 70812 92678
rect 70868 92652 70900 92678
rect 70964 92652 70970 92716
rect 70868 92622 70916 92652
rect 70807 92620 70916 92622
rect 70807 92617 70873 92620
rect 69606 92516 69612 92580
rect 69676 92578 69682 92580
rect 70301 92578 70367 92581
rect 69676 92576 70367 92578
rect 69676 92520 70306 92576
rect 70362 92520 70367 92576
rect 69676 92518 70367 92520
rect 69676 92516 69682 92518
rect 70301 92515 70367 92518
rect 68553 92442 68619 92445
rect 75729 92442 75795 92445
rect 68553 92440 75795 92442
rect 68553 92384 68558 92440
rect 68614 92384 75734 92440
rect 75790 92384 75795 92440
rect 68553 92382 75795 92384
rect 68553 92379 68619 92382
rect 75729 92379 75795 92382
rect 91277 92442 91343 92445
rect 92974 92442 92980 92444
rect 91277 92440 92980 92442
rect 91277 92384 91282 92440
rect 91338 92384 92980 92440
rect 91277 92382 92980 92384
rect 91277 92379 91343 92382
rect 92974 92380 92980 92382
rect 93044 92380 93050 92444
rect 93853 92442 93919 92445
rect 95182 92442 95188 92444
rect 93853 92440 95188 92442
rect 93853 92384 93858 92440
rect 93914 92384 95188 92440
rect 93853 92382 95188 92384
rect 93853 92379 93919 92382
rect 95182 92380 95188 92382
rect 95252 92380 95258 92444
rect 89805 92306 89871 92309
rect 114553 92306 114619 92309
rect 89805 92304 114619 92306
rect 89805 92248 89810 92304
rect 89866 92248 114558 92304
rect 114614 92248 114619 92304
rect 89805 92246 114619 92248
rect 89805 92243 89871 92246
rect 114553 92243 114619 92246
rect 54477 91762 54543 91765
rect 220813 91762 220879 91765
rect 54477 91760 220879 91762
rect 54477 91704 54482 91760
rect 54538 91704 220818 91760
rect 220874 91704 220879 91760
rect 54477 91702 220879 91704
rect 54477 91699 54543 91702
rect 220813 91699 220879 91702
rect 92565 91490 92631 91493
rect 95049 91490 95115 91493
rect 92565 91488 95115 91490
rect 92565 91432 92570 91488
rect 92626 91432 95054 91488
rect 95110 91432 95115 91488
rect 92565 91430 95115 91432
rect 92565 91427 92631 91430
rect 95049 91427 95115 91430
rect 68870 91020 68876 91084
rect 68940 91082 68946 91084
rect 72233 91082 72299 91085
rect 68940 91080 72299 91082
rect 68940 91024 72238 91080
rect 72294 91024 72299 91080
rect 68940 91022 72299 91024
rect 68940 91020 68946 91022
rect 72233 91019 72299 91022
rect 92749 91082 92815 91085
rect 109033 91082 109099 91085
rect 92749 91080 109099 91082
rect 92749 91024 92754 91080
rect 92810 91024 109038 91080
rect 109094 91024 109099 91080
rect 92749 91022 109099 91024
rect 92749 91019 92815 91022
rect 109033 91019 109099 91022
rect 57697 90946 57763 90949
rect 71129 90946 71195 90949
rect 57697 90944 71195 90946
rect 57697 90888 57702 90944
rect 57758 90888 71134 90944
rect 71190 90888 71195 90944
rect 57697 90886 71195 90888
rect 57697 90883 57763 90886
rect 71129 90883 71195 90886
rect 71630 90884 71636 90948
rect 71700 90946 71706 90948
rect 81433 90946 81499 90949
rect 71700 90944 81499 90946
rect 71700 90888 81438 90944
rect 81494 90888 81499 90944
rect 71700 90886 81499 90888
rect 71700 90884 71706 90886
rect 81433 90883 81499 90886
rect 90725 90946 90791 90949
rect 98637 90946 98703 90949
rect 90725 90944 98703 90946
rect 90725 90888 90730 90944
rect 90786 90888 98642 90944
rect 98698 90888 98703 90944
rect 90725 90886 98703 90888
rect 90725 90883 90791 90886
rect 98637 90883 98703 90886
rect 50981 90810 51047 90813
rect 77937 90810 78003 90813
rect 50981 90808 78003 90810
rect 50981 90752 50986 90808
rect 51042 90752 77942 90808
rect 77998 90752 78003 90808
rect 50981 90750 78003 90752
rect 50981 90747 51047 90750
rect 77937 90747 78003 90750
rect 80605 90810 80671 90813
rect 94078 90810 94084 90812
rect 80605 90808 94084 90810
rect 80605 90752 80610 90808
rect 80666 90752 94084 90808
rect 80605 90750 94084 90752
rect 80605 90747 80671 90750
rect 94078 90748 94084 90750
rect 94148 90748 94154 90812
rect 77477 90674 77543 90677
rect 92565 90674 92631 90677
rect 77477 90672 92631 90674
rect 77477 90616 77482 90672
rect 77538 90616 92570 90672
rect 92626 90616 92631 90672
rect 77477 90614 92631 90616
rect 77477 90611 77543 90614
rect 92565 90611 92631 90614
rect 82077 89722 82143 89725
rect 103830 89722 103836 89724
rect 82077 89720 103836 89722
rect 82077 89664 82082 89720
rect 82138 89664 103836 89720
rect 82077 89662 103836 89664
rect 82077 89659 82143 89662
rect 103830 89660 103836 89662
rect 103900 89660 103906 89724
rect 89529 89586 89595 89589
rect 93894 89586 93900 89588
rect 89529 89584 93900 89586
rect 89529 89528 89534 89584
rect 89590 89528 93900 89584
rect 89529 89526 93900 89528
rect 89529 89523 89595 89526
rect 93894 89524 93900 89526
rect 93964 89524 93970 89588
rect 58617 89042 58683 89045
rect 224902 89042 224908 89044
rect 58617 89040 224908 89042
rect 58617 88984 58622 89040
rect 58678 88984 224908 89040
rect 58617 88982 224908 88984
rect 58617 88979 58683 88982
rect 224902 88980 224908 88982
rect 224972 88980 224978 89044
rect 58985 88226 59051 88229
rect 74809 88226 74875 88229
rect 58985 88224 74875 88226
rect 58985 88168 58990 88224
rect 59046 88168 74814 88224
rect 74870 88168 74875 88224
rect 58985 88166 74875 88168
rect 58985 88163 59051 88166
rect 74809 88163 74875 88166
rect 88701 88226 88767 88229
rect 89529 88226 89595 88229
rect 88701 88224 89595 88226
rect 88701 88168 88706 88224
rect 88762 88168 89534 88224
rect 89590 88168 89595 88224
rect 88701 88166 89595 88168
rect 88701 88163 88767 88166
rect 89529 88163 89595 88166
rect 82997 88090 83063 88093
rect 95969 88090 96035 88093
rect 82997 88088 96035 88090
rect 82997 88032 83002 88088
rect 83058 88032 95974 88088
rect 96030 88032 96035 88088
rect 82997 88030 96035 88032
rect 82997 88027 83063 88030
rect 95969 88027 96035 88030
rect 89529 87954 89595 87957
rect 102225 87954 102291 87957
rect 89529 87952 102291 87954
rect 89529 87896 89534 87952
rect 89590 87896 102230 87952
rect 102286 87896 102291 87952
rect 89529 87894 102291 87896
rect 89529 87891 89595 87894
rect 102225 87891 102291 87894
rect 84653 86866 84719 86869
rect 114645 86866 114711 86869
rect 115749 86866 115815 86869
rect 84653 86864 115815 86866
rect 84653 86808 84658 86864
rect 84714 86808 114650 86864
rect 114706 86808 115754 86864
rect 115810 86808 115815 86864
rect 84653 86806 115815 86808
rect 84653 86803 84719 86806
rect 114645 86803 114711 86806
rect 115749 86803 115815 86806
rect 57881 86322 57947 86325
rect 188337 86322 188403 86325
rect 57881 86320 188403 86322
rect 57881 86264 57886 86320
rect 57942 86264 188342 86320
rect 188398 86264 188403 86320
rect 57881 86262 188403 86264
rect 57881 86259 57947 86262
rect 188337 86259 188403 86262
rect 115749 86186 115815 86189
rect 357433 86186 357499 86189
rect 115749 86184 357499 86186
rect 115749 86128 115754 86184
rect 115810 86128 357438 86184
rect 357494 86128 357499 86184
rect 115749 86126 357499 86128
rect 115749 86123 115815 86126
rect 357433 86123 357499 86126
rect 582833 86186 582899 86189
rect 583520 86186 584960 86276
rect 582833 86184 584960 86186
rect 582833 86128 582838 86184
rect 582894 86128 584960 86184
rect 582833 86126 584960 86128
rect 582833 86123 582899 86126
rect 583520 86036 584960 86126
rect 79501 85506 79567 85509
rect 103605 85506 103671 85509
rect 79501 85504 103671 85506
rect 79501 85448 79506 85504
rect 79562 85448 103610 85504
rect 103666 85448 103671 85504
rect 79501 85446 103671 85448
rect 79501 85443 79567 85446
rect 103605 85443 103671 85446
rect 83549 85370 83615 85373
rect 105629 85370 105695 85373
rect 83549 85368 105695 85370
rect 83549 85312 83554 85368
rect 83610 85312 105634 85368
rect 105690 85312 105695 85368
rect 83549 85310 105695 85312
rect 83549 85307 83615 85310
rect 105629 85307 105695 85310
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 69841 84146 69907 84149
rect 274633 84146 274699 84149
rect 69841 84144 274699 84146
rect 69841 84088 69846 84144
rect 69902 84088 274638 84144
rect 274694 84088 274699 84144
rect 69841 84086 274699 84088
rect 69841 84083 69907 84086
rect 274633 84083 274699 84086
rect 274633 83466 274699 83469
rect 320173 83466 320239 83469
rect 274633 83464 320239 83466
rect 274633 83408 274638 83464
rect 274694 83408 320178 83464
rect 320234 83408 320239 83464
rect 274633 83406 320239 83408
rect 274633 83403 274699 83406
rect 320173 83403 320239 83406
rect 87597 76530 87663 76533
rect 211654 76530 211660 76532
rect 87597 76528 211660 76530
rect 87597 76472 87602 76528
rect 87658 76472 211660 76528
rect 87597 76470 211660 76472
rect 87597 76467 87663 76470
rect 211654 76468 211660 76470
rect 211724 76468 211730 76532
rect 77201 73810 77267 73813
rect 208894 73810 208900 73812
rect 77201 73808 208900 73810
rect 77201 73752 77206 73808
rect 77262 73752 208900 73808
rect 77201 73750 208900 73752
rect 77201 73747 77267 73750
rect 208894 73748 208900 73750
rect 208964 73748 208970 73812
rect 582741 72994 582807 72997
rect 583520 72994 584960 73084
rect 582741 72992 584960 72994
rect 582741 72936 582746 72992
rect 582802 72936 584960 72992
rect 582741 72934 584960 72936
rect 582741 72931 582807 72934
rect 583520 72844 584960 72934
rect 83457 72450 83523 72453
rect 229686 72450 229692 72452
rect 83457 72448 229692 72450
rect 83457 72392 83462 72448
rect 83518 72392 229692 72448
rect 83457 72390 229692 72392
rect 83457 72387 83523 72390
rect 229686 72388 229692 72390
rect 229756 72388 229762 72452
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 91001 71090 91067 71093
rect 210366 71090 210372 71092
rect 91001 71088 210372 71090
rect 91001 71032 91006 71088
rect 91062 71032 210372 71088
rect 91001 71030 210372 71032
rect 91001 71027 91067 71030
rect 210366 71028 210372 71030
rect 210436 71028 210442 71092
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 67541 47562 67607 47565
rect 226558 47562 226564 47564
rect 67541 47560 226564 47562
rect 67541 47504 67546 47560
rect 67602 47504 226564 47560
rect 67541 47502 226564 47504
rect 67541 47499 67607 47502
rect 226558 47500 226564 47502
rect 226628 47500 226634 47564
rect 582649 46338 582715 46341
rect 583520 46338 584960 46428
rect 582649 46336 584960 46338
rect 582649 46280 582654 46336
rect 582710 46280 584960 46336
rect 582649 46278 584960 46280
rect 582649 46275 582715 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 6821 39266 6887 39269
rect 196014 39266 196020 39268
rect 6821 39264 196020 39266
rect 6821 39208 6826 39264
rect 6882 39208 196020 39264
rect 6821 39206 196020 39208
rect 6821 39203 6887 39206
rect 196014 39204 196020 39206
rect 196084 39204 196090 39268
rect 45461 36546 45527 36549
rect 223982 36546 223988 36548
rect 45461 36544 223988 36546
rect 45461 36488 45466 36544
rect 45522 36488 223988 36544
rect 45461 36486 223988 36488
rect 45461 36483 45527 36486
rect 223982 36484 223988 36486
rect 224052 36484 224058 36548
rect 42701 35186 42767 35189
rect 222326 35186 222332 35188
rect 42701 35184 222332 35186
rect 42701 35128 42706 35184
rect 42762 35128 222332 35184
rect 42701 35126 222332 35128
rect 42701 35123 42767 35126
rect 222326 35124 222332 35126
rect 222396 35124 222402 35188
rect 23381 33826 23447 33829
rect 219198 33826 219204 33828
rect 23381 33824 219204 33826
rect 23381 33768 23386 33824
rect 23442 33768 219204 33824
rect 23381 33766 219204 33768
rect 23381 33763 23447 33766
rect 219198 33764 219204 33766
rect 219268 33764 219274 33828
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 92381 30970 92447 30973
rect 230422 30970 230428 30972
rect 92381 30968 230428 30970
rect 92381 30912 92386 30968
rect 92442 30912 230428 30968
rect 92381 30910 230428 30912
rect 92381 30907 92447 30910
rect 230422 30908 230428 30910
rect 230492 30908 230498 30972
rect 85481 29610 85547 29613
rect 237782 29610 237788 29612
rect 85481 29608 237788 29610
rect 85481 29552 85486 29608
rect 85542 29552 237788 29608
rect 85481 29550 237788 29552
rect 85481 29547 85547 29550
rect 237782 29548 237788 29550
rect 237852 29548 237858 29612
rect 74441 28250 74507 28253
rect 227662 28250 227668 28252
rect 74441 28248 227668 28250
rect 74441 28192 74446 28248
rect 74502 28192 227668 28248
rect 74441 28190 227668 28192
rect 74441 28187 74507 28190
rect 227662 28188 227668 28190
rect 227732 28188 227738 28252
rect 72509 25530 72575 25533
rect 226374 25530 226380 25532
rect 72509 25528 226380 25530
rect 72509 25472 72514 25528
rect 72570 25472 226380 25528
rect 72509 25470 226380 25472
rect 72509 25467 72575 25470
rect 226374 25468 226380 25470
rect 226444 25468 226450 25532
rect 53741 24170 53807 24173
rect 222694 24170 222700 24172
rect 53741 24168 222700 24170
rect 53741 24112 53746 24168
rect 53802 24112 222700 24168
rect 53741 24110 222700 24112
rect 53741 24107 53807 24110
rect 222694 24108 222700 24110
rect 222764 24108 222770 24172
rect 41321 22674 41387 22677
rect 204294 22674 204300 22676
rect 41321 22672 204300 22674
rect 41321 22616 41326 22672
rect 41382 22616 204300 22672
rect 41321 22614 204300 22616
rect 41321 22611 41387 22614
rect 204294 22612 204300 22614
rect 204364 22612 204370 22676
rect 27521 21314 27587 21317
rect 201534 21314 201540 21316
rect 27521 21312 201540 21314
rect 27521 21256 27526 21312
rect 27582 21256 201540 21312
rect 27521 21254 201540 21256
rect 27521 21251 27587 21254
rect 201534 21252 201540 21254
rect 201604 21252 201610 21316
rect 582557 19818 582623 19821
rect 583520 19818 584960 19908
rect 582557 19816 584960 19818
rect 582557 19760 582562 19816
rect 582618 19760 584960 19816
rect 582557 19758 584960 19760
rect 582557 19755 582623 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 70209 11658 70275 11661
rect 208342 11658 208348 11660
rect 70209 11656 208348 11658
rect 70209 11600 70214 11656
rect 70270 11600 208348 11656
rect 70209 11598 208348 11600
rect 70209 11595 70275 11598
rect 208342 11596 208348 11598
rect 208412 11596 208418 11660
rect 105721 8938 105787 8941
rect 233182 8938 233188 8940
rect 105721 8936 233188 8938
rect 105721 8880 105726 8936
rect 105782 8880 233188 8936
rect 105721 8878 233188 8880
rect 105721 8875 105787 8878
rect 233182 8876 233188 8878
rect 233252 8876 233258 8940
rect 101029 7578 101095 7581
rect 213862 7578 213868 7580
rect 101029 7576 213868 7578
rect 101029 7520 101034 7576
rect 101090 7520 213868 7576
rect 101029 7518 213868 7520
rect 101029 7515 101095 7518
rect 213862 7516 213868 7518
rect 213932 7516 213938 7580
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 130326 4932 130332 4996
rect 130396 4994 130402 4996
rect 136449 4994 136515 4997
rect 130396 4992 136515 4994
rect 130396 4936 136454 4992
rect 136510 4936 136515 4992
rect 130396 4934 136515 4936
rect 130396 4932 130402 4934
rect 136449 4931 136515 4934
rect 77385 4858 77451 4861
rect 215886 4858 215892 4860
rect 77385 4856 215892 4858
rect 77385 4800 77390 4856
rect 77446 4800 215892 4856
rect 77385 4798 215892 4800
rect 77385 4795 77451 4798
rect 215886 4796 215892 4798
rect 215956 4796 215962 4860
rect 16481 4042 16547 4045
rect 18229 4042 18295 4045
rect 16481 4040 18295 4042
rect 16481 3984 16486 4040
rect 16542 3984 18234 4040
rect 18290 3984 18295 4040
rect 16481 3982 18295 3984
rect 16481 3979 16547 3982
rect 18229 3979 18295 3982
rect 238518 3980 238524 4044
rect 238588 4042 238594 4044
rect 239305 4042 239371 4045
rect 238588 4040 239371 4042
rect 238588 3984 239310 4040
rect 239366 3984 239371 4040
rect 238588 3982 239371 3984
rect 238588 3980 238594 3982
rect 239305 3979 239371 3982
rect 348049 4042 348115 4045
rect 356053 4042 356119 4045
rect 348049 4040 356119 4042
rect 348049 3984 348054 4040
rect 348110 3984 356058 4040
rect 356114 3984 356119 4040
rect 348049 3982 356119 3984
rect 348049 3979 348115 3982
rect 356053 3979 356119 3982
rect 231117 3906 231183 3909
rect 244273 3906 244339 3909
rect 231117 3904 244339 3906
rect 231117 3848 231122 3904
rect 231178 3848 244278 3904
rect 244334 3848 244339 3904
rect 231117 3846 244339 3848
rect 231117 3843 231183 3846
rect 244273 3843 244339 3846
rect 98637 3634 98703 3637
rect 99046 3634 99052 3636
rect 98637 3632 99052 3634
rect 98637 3576 98642 3632
rect 98698 3576 99052 3632
rect 98637 3574 99052 3576
rect 98637 3571 98703 3574
rect 99046 3572 99052 3574
rect 99116 3572 99122 3636
rect 116393 3634 116459 3637
rect 117078 3634 117084 3636
rect 116393 3632 117084 3634
rect 116393 3576 116398 3632
rect 116454 3576 117084 3632
rect 116393 3574 117084 3576
rect 116393 3571 116459 3574
rect 117078 3572 117084 3574
rect 117148 3572 117154 3636
rect 244273 3634 244339 3637
rect 245193 3634 245259 3637
rect 244273 3632 245259 3634
rect 244273 3576 244278 3632
rect 244334 3576 245198 3632
rect 245254 3576 245259 3632
rect 244273 3574 245259 3576
rect 244273 3571 244339 3574
rect 245193 3571 245259 3574
rect 85665 3498 85731 3501
rect 105537 3498 105603 3501
rect 85665 3496 105603 3498
rect 85665 3440 85670 3496
rect 85726 3440 105542 3496
rect 105598 3440 105603 3496
rect 85665 3438 105603 3440
rect 85665 3435 85731 3438
rect 105537 3435 105603 3438
rect 110505 3498 110571 3501
rect 111558 3498 111564 3500
rect 110505 3496 111564 3498
rect 110505 3440 110510 3496
rect 110566 3440 111564 3496
rect 110505 3438 111564 3440
rect 110505 3435 110571 3438
rect 111558 3436 111564 3438
rect 111628 3436 111634 3500
rect 112805 3498 112871 3501
rect 126237 3498 126303 3501
rect 112805 3496 126303 3498
rect 112805 3440 112810 3496
rect 112866 3440 126242 3496
rect 126298 3440 126303 3496
rect 112805 3438 126303 3440
rect 112805 3435 112871 3438
rect 126237 3435 126303 3438
rect 240358 3436 240364 3500
rect 240428 3498 240434 3500
rect 240501 3498 240567 3501
rect 240428 3496 240567 3498
rect 240428 3440 240506 3496
rect 240562 3440 240567 3496
rect 240428 3438 240567 3440
rect 240428 3436 240434 3438
rect 240501 3435 240567 3438
rect 244917 3498 244983 3501
rect 254669 3498 254735 3501
rect 244917 3496 254735 3498
rect 244917 3440 244922 3496
rect 244978 3440 254674 3496
rect 254730 3440 254735 3496
rect 244917 3438 254735 3440
rect 244917 3435 244983 3438
rect 254669 3435 254735 3438
rect 8753 3362 8819 3365
rect 17217 3362 17283 3365
rect 8753 3360 17283 3362
rect 8753 3304 8758 3360
rect 8814 3304 17222 3360
rect 17278 3304 17283 3360
rect 8753 3302 17283 3304
rect 8753 3299 8819 3302
rect 17217 3299 17283 3302
rect 31293 3362 31359 3365
rect 54477 3362 54543 3365
rect 31293 3360 54543 3362
rect 31293 3304 31298 3360
rect 31354 3304 54482 3360
rect 54538 3304 54543 3360
rect 31293 3302 54543 3304
rect 31293 3299 31359 3302
rect 54477 3299 54543 3302
rect 63217 3362 63283 3365
rect 88977 3362 89043 3365
rect 63217 3360 89043 3362
rect 63217 3304 63222 3360
rect 63278 3304 88982 3360
rect 89038 3304 89043 3360
rect 63217 3302 89043 3304
rect 63217 3299 63283 3302
rect 88977 3299 89043 3302
rect 109309 3362 109375 3365
rect 152457 3362 152523 3365
rect 109309 3360 152523 3362
rect 109309 3304 109314 3360
rect 109370 3304 152462 3360
rect 152518 3304 152523 3360
rect 109309 3302 152523 3304
rect 109309 3299 109375 3302
rect 152457 3299 152523 3302
rect 242157 3362 242223 3365
rect 290181 3362 290247 3365
rect 242157 3360 290247 3362
rect 242157 3304 242162 3360
rect 242218 3304 290186 3360
rect 290242 3304 290247 3360
rect 242157 3302 290247 3304
rect 242157 3299 242223 3302
rect 290181 3299 290247 3302
rect 324957 3362 325023 3365
rect 332685 3362 332751 3365
rect 324957 3360 332751 3362
rect 324957 3304 324962 3360
rect 325018 3304 332690 3360
rect 332746 3304 332751 3360
rect 324957 3302 332751 3304
rect 324957 3299 325023 3302
rect 332685 3299 332751 3302
rect 335997 3362 336063 3365
rect 350441 3362 350507 3365
rect 335997 3360 350507 3362
rect 335997 3304 336002 3360
rect 336058 3304 350446 3360
rect 350502 3304 350507 3360
rect 335997 3302 350507 3304
rect 335997 3299 336063 3302
rect 350441 3299 350507 3302
<< via3 >>
rect 263364 702612 263428 702676
rect 264100 702476 264164 702540
rect 124260 587964 124324 588028
rect 75868 584836 75932 584900
rect 111748 583748 111812 583812
rect 75684 581028 75748 581092
rect 78444 581028 78508 581092
rect 70900 580816 70964 580820
rect 70900 580760 70950 580816
rect 70950 580760 70964 580816
rect 70900 580756 70964 580760
rect 83964 580756 84028 580820
rect 88380 580756 88444 580820
rect 130332 578308 130396 578372
rect 97212 554100 97276 554164
rect 67772 548252 67836 548316
rect 104940 547844 105004 547908
rect 96660 547028 96724 547092
rect 69428 542132 69492 542196
rect 94084 541588 94148 541652
rect 67772 539820 67836 539884
rect 91508 538188 91572 538252
rect 75868 535528 75932 535532
rect 75868 535472 75918 535528
rect 75918 535472 75932 535528
rect 75868 535468 75932 535472
rect 96660 533292 96724 533356
rect 94084 531932 94148 531996
rect 79916 527716 79980 527780
rect 94452 520916 94516 520980
rect 77156 518060 77220 518124
rect 100708 507860 100772 507924
rect 75684 468420 75748 468484
rect 106412 462980 106476 463044
rect 69612 462844 69676 462908
rect 88748 462844 88812 462908
rect 69612 461484 69676 461548
rect 78444 460124 78508 460188
rect 92612 460124 92676 460188
rect 114508 458764 114572 458828
rect 72556 454684 72620 454748
rect 113220 453188 113284 453252
rect 107700 449108 107764 449172
rect 123340 446388 123404 446452
rect 88380 444892 88444 444956
rect 97212 444212 97276 444276
rect 66116 443532 66180 443596
rect 72740 436188 72804 436252
rect 86172 436188 86236 436252
rect 103284 436188 103348 436252
rect 78260 436052 78324 436116
rect 100524 436052 100588 436116
rect 82124 435916 82188 435980
rect 83964 435916 84028 435980
rect 71636 435372 71700 435436
rect 73476 434828 73540 434892
rect 90956 434828 91020 434892
rect 70164 434692 70228 434756
rect 75684 434692 75748 434756
rect 85436 434692 85500 434756
rect 83412 434556 83476 434620
rect 83596 434420 83660 434484
rect 74580 434284 74644 434348
rect 75868 434284 75932 434348
rect 80284 434344 80348 434348
rect 80284 434288 80298 434344
rect 80298 434288 80348 434344
rect 80284 434284 80348 434288
rect 80652 434284 80716 434348
rect 81940 434344 82004 434348
rect 81940 434288 81954 434344
rect 81954 434288 82004 434344
rect 81940 434284 82004 434288
rect 85804 434344 85868 434348
rect 85804 434288 85854 434344
rect 85854 434288 85868 434344
rect 85804 434284 85868 434288
rect 87092 434344 87156 434348
rect 87092 434288 87142 434344
rect 87142 434288 87156 434344
rect 87092 434284 87156 434288
rect 93900 434284 93964 434348
rect 97212 434344 97276 434348
rect 97212 434288 97226 434344
rect 97226 434288 97276 434344
rect 97212 434284 97276 434288
rect 102180 434284 102244 434348
rect 104204 434344 104268 434348
rect 104204 434288 104218 434344
rect 104218 434288 104268 434344
rect 104204 434284 104268 434288
rect 108252 434344 108316 434348
rect 108252 434288 108266 434344
rect 108266 434288 108316 434344
rect 108252 434284 108316 434288
rect 97396 433876 97460 433940
rect 109172 433876 109236 433940
rect 70900 433800 70964 433804
rect 70900 433744 70914 433800
rect 70914 433744 70964 433800
rect 70900 433740 70964 433744
rect 84700 433740 84764 433804
rect 98132 433740 98196 433804
rect 101996 433740 102060 433804
rect 78444 433664 78508 433668
rect 78444 433608 78458 433664
rect 78458 433608 78508 433664
rect 78444 433604 78508 433608
rect 79732 433604 79796 433668
rect 87276 433664 87340 433668
rect 87276 433608 87326 433664
rect 87326 433608 87340 433664
rect 87276 433604 87340 433608
rect 89668 433604 89732 433668
rect 91324 433604 91388 433668
rect 93716 433604 93780 433668
rect 95188 433664 95252 433668
rect 95188 433608 95202 433664
rect 95202 433608 95252 433664
rect 95188 433604 95252 433608
rect 98500 433604 98564 433668
rect 99972 433604 100036 433668
rect 105124 433664 105188 433668
rect 105124 433608 105174 433664
rect 105174 433608 105188 433664
rect 105124 433604 105188 433608
rect 106780 433604 106844 433668
rect 111196 433604 111260 433668
rect 67404 433256 67468 433260
rect 67404 433200 67454 433256
rect 67454 433200 67468 433256
rect 67404 433196 67468 433200
rect 112116 432788 112180 432852
rect 112116 426532 112180 426596
rect 61884 425172 61948 425236
rect 66852 422180 66916 422244
rect 112300 420276 112364 420340
rect 66852 420140 66916 420204
rect 59124 411300 59188 411364
rect 67404 409728 67468 409732
rect 67404 409672 67454 409728
rect 67454 409672 67468 409728
rect 67404 409668 67468 409672
rect 114508 409668 114572 409732
rect 66116 408852 66180 408916
rect 115060 408580 115124 408644
rect 41276 407008 41340 407012
rect 41276 406952 41290 407008
rect 41290 406952 41340 407008
rect 41276 406948 41340 406952
rect 57836 406948 57900 407012
rect 57836 405724 57900 405788
rect 69428 397700 69492 397764
rect 123340 396612 123404 396676
rect 113220 396340 113284 396404
rect 69612 392124 69676 392188
rect 107700 391852 107764 391916
rect 82124 391096 82188 391100
rect 82124 391040 82138 391096
rect 82138 391040 82188 391096
rect 82124 391036 82188 391040
rect 85436 391096 85500 391100
rect 85436 391040 85486 391096
rect 85486 391040 85500 391096
rect 85436 391036 85500 391040
rect 88748 391036 88812 391100
rect 92612 391036 92676 391100
rect 100708 390960 100772 390964
rect 100708 390904 100722 390960
rect 100722 390904 100772 390960
rect 100708 390900 100772 390904
rect 78444 390628 78508 390692
rect 107700 390688 107764 390692
rect 107700 390632 107750 390688
rect 107750 390632 107764 390688
rect 107700 390628 107764 390632
rect 108252 390628 108316 390692
rect 72556 390356 72620 390420
rect 77156 390416 77220 390420
rect 77156 390360 77206 390416
rect 77206 390360 77220 390416
rect 77156 390356 77220 390360
rect 104940 390356 105004 390420
rect 106412 390356 106476 390420
rect 128676 389268 128740 389332
rect 71820 389056 71884 389060
rect 71820 389000 71870 389056
rect 71870 389000 71884 389056
rect 71820 388996 71884 389000
rect 79916 388996 79980 389060
rect 91508 388996 91572 389060
rect 94452 388996 94516 389060
rect 124260 388996 124324 389060
rect 69612 388860 69676 388924
rect 100524 388452 100588 388516
rect 103284 388452 103348 388516
rect 106412 388316 106476 388380
rect 80652 387908 80716 387972
rect 111012 387772 111076 387836
rect 86172 387636 86236 387700
rect 61700 387500 61764 387564
rect 99972 387092 100036 387156
rect 111748 387092 111812 387156
rect 105124 386956 105188 387020
rect 55076 386472 55140 386476
rect 55076 386416 55126 386472
rect 55126 386416 55140 386472
rect 55076 386412 55140 386416
rect 78260 386276 78324 386340
rect 97396 385596 97460 385660
rect 106780 385596 106844 385660
rect 75868 385052 75932 385116
rect 84700 385052 84764 385116
rect 80284 384372 80348 384436
rect 71820 384236 71884 384300
rect 85804 383692 85868 383756
rect 133828 383692 133892 383756
rect 106044 382332 106108 382396
rect 111196 381516 111260 381580
rect 74580 380836 74644 380900
rect 95188 380156 95252 380220
rect 81940 379476 82004 379540
rect 93900 378660 93964 378724
rect 89668 377300 89732 377364
rect 98132 373220 98196 373284
rect 107700 369004 107764 369068
rect 102180 364924 102244 364988
rect 73476 343708 73540 343772
rect 75684 340852 75748 340916
rect 82860 339492 82924 339556
rect 83596 339552 83660 339556
rect 83596 339496 83610 339552
rect 83610 339496 83660 339552
rect 83596 339492 83660 339496
rect 70164 337996 70228 338060
rect 102732 335412 102796 335476
rect 66116 334052 66180 334116
rect 91324 333236 91388 333300
rect 91508 332692 91572 332756
rect 92980 332692 93044 332756
rect 93716 332692 93780 332756
rect 79180 332556 79244 332620
rect 108252 330380 108316 330444
rect 255452 330380 255516 330444
rect 97948 329836 98012 329900
rect 87092 329020 87156 329084
rect 71452 328476 71516 328540
rect 95004 326980 95068 327044
rect 252508 324940 252572 325004
rect 92980 323580 93044 323644
rect 82860 322900 82924 322964
rect 104204 322084 104268 322148
rect 108988 320996 109052 321060
rect 97212 320860 97276 320924
rect 191052 320180 191116 320244
rect 114508 319500 114572 319564
rect 79180 319364 79244 319428
rect 72740 318820 72804 318884
rect 83412 318684 83476 318748
rect 258396 318004 258460 318068
rect 252692 316236 252756 316300
rect 254532 315284 254596 315348
rect 264100 310796 264164 310860
rect 106780 307804 106844 307868
rect 52316 304948 52380 305012
rect 218652 304948 218716 305012
rect 87276 304132 87340 304196
rect 186820 303860 186884 303924
rect 242020 303860 242084 303924
rect 215892 303724 215956 303788
rect 260236 303724 260300 303788
rect 192708 303588 192772 303652
rect 237788 303588 237852 303652
rect 260052 303588 260116 303652
rect 240364 302228 240428 302292
rect 254164 301548 254228 301612
rect 193444 301412 193508 301476
rect 193260 301140 193324 301204
rect 210372 301140 210436 301204
rect 222700 301140 222764 301204
rect 258580 301140 258644 301204
rect 208900 301004 208964 301068
rect 213684 301004 213748 301068
rect 219388 301004 219452 301068
rect 221228 301004 221292 301068
rect 223804 301004 223868 301068
rect 230428 301004 230492 301068
rect 232084 301004 232148 301068
rect 233188 301004 233252 301068
rect 234844 301004 234908 301068
rect 196020 300928 196084 300932
rect 196020 300872 196070 300928
rect 196070 300872 196084 300928
rect 196020 300868 196084 300872
rect 197492 300868 197556 300932
rect 198780 300928 198844 300932
rect 198780 300872 198830 300928
rect 198830 300872 198844 300928
rect 198780 300868 198844 300872
rect 201540 300868 201604 300932
rect 203012 300928 203076 300932
rect 203012 300872 203062 300928
rect 203062 300872 203076 300928
rect 203012 300868 203076 300872
rect 204300 300868 204364 300932
rect 205588 300868 205652 300932
rect 207060 300928 207124 300932
rect 207060 300872 207110 300928
rect 207110 300872 207124 300928
rect 207060 300868 207124 300872
rect 208348 300868 208412 300932
rect 211660 300868 211724 300932
rect 213868 300868 213932 300932
rect 214420 300868 214484 300932
rect 216076 300868 216140 300932
rect 216812 300868 216876 300932
rect 219572 300928 219636 300932
rect 219572 300872 219586 300928
rect 219586 300872 219636 300928
rect 219572 300868 219636 300872
rect 220860 300868 220924 300932
rect 222332 300868 222396 300932
rect 223988 300928 224052 300932
rect 223988 300872 224038 300928
rect 224038 300872 224052 300928
rect 223988 300868 224052 300872
rect 225092 300868 225156 300932
rect 226380 300928 226444 300932
rect 226380 300872 226394 300928
rect 226394 300872 226444 300928
rect 226380 300868 226444 300872
rect 226564 300868 226628 300932
rect 227668 300868 227732 300932
rect 229692 300928 229756 300932
rect 229692 300872 229742 300928
rect 229742 300872 229756 300928
rect 229692 300868 229756 300872
rect 230980 300928 231044 300932
rect 230980 300872 231030 300928
rect 231030 300872 231044 300928
rect 230980 300868 231044 300872
rect 232268 300928 232332 300932
rect 232268 300872 232318 300928
rect 232318 300872 232332 300928
rect 232268 300868 232332 300872
rect 233372 300928 233436 300932
rect 233372 300872 233386 300928
rect 233386 300872 233436 300928
rect 233372 300868 233436 300872
rect 234660 300868 234724 300932
rect 236500 300868 236564 300932
rect 238156 300868 238220 300932
rect 238708 300868 238772 300932
rect 244412 300868 244476 300932
rect 254532 300188 254596 300252
rect 255452 299780 255516 299844
rect 193444 298828 193508 298892
rect 191052 298692 191116 298756
rect 255268 298420 255332 298484
rect 252876 297876 252940 297940
rect 67772 296924 67836 296988
rect 61884 296788 61948 296852
rect 255268 294476 255332 294540
rect 255452 294340 255516 294404
rect 255820 293796 255884 293860
rect 255452 293116 255516 293180
rect 103836 292708 103900 292772
rect 90956 292572 91020 292636
rect 116532 291756 116596 291820
rect 100156 291348 100220 291412
rect 252876 291348 252940 291412
rect 103836 289852 103900 289916
rect 258580 289036 258644 289100
rect 70164 288356 70228 288420
rect 72924 287676 72988 287740
rect 70164 287132 70228 287196
rect 71636 286996 71700 287060
rect 97948 285364 98012 285428
rect 104940 284412 105004 284476
rect 122604 284276 122668 284340
rect 260236 284820 260300 284884
rect 74212 284200 74276 284204
rect 74212 284144 74262 284200
rect 74262 284144 74276 284200
rect 74212 284140 74276 284144
rect 71636 283732 71700 283796
rect 71084 283460 71148 283524
rect 73476 283520 73540 283524
rect 73476 283464 73526 283520
rect 73526 283464 73540 283520
rect 73476 283460 73540 283464
rect 95188 283460 95252 283524
rect 96660 283460 96724 283524
rect 260052 283460 260116 283524
rect 65932 283188 65996 283252
rect 118004 282916 118068 282980
rect 99972 282644 100036 282708
rect 101996 282644 102060 282708
rect 62988 282100 63052 282164
rect 67956 280468 68020 280532
rect 255820 279380 255884 279444
rect 193260 276660 193324 276724
rect 52316 276116 52380 276180
rect 67772 275844 67836 275908
rect 67772 274756 67836 274820
rect 118740 274680 118804 274684
rect 118740 274624 118790 274680
rect 118790 274624 118804 274680
rect 118740 274620 118804 274624
rect 121684 274620 121748 274684
rect 112300 271960 112364 271964
rect 112300 271904 112314 271960
rect 112314 271904 112364 271960
rect 112300 271900 112364 271904
rect 115980 271900 116044 271964
rect 98500 271084 98564 271148
rect 255820 271084 255884 271148
rect 111748 270404 111812 270468
rect 61884 269180 61948 269244
rect 106780 269240 106844 269244
rect 106780 269184 106830 269240
rect 106830 269184 106844 269240
rect 106780 269180 106844 269184
rect 100156 267276 100220 267340
rect 110644 267276 110708 267340
rect 109540 267004 109604 267068
rect 64644 266460 64708 266524
rect 99236 266324 99300 266388
rect 263364 266460 263428 266524
rect 263732 266460 263796 266524
rect 253980 265916 254044 265980
rect 254164 264964 254228 265028
rect 115060 263664 115124 263668
rect 115060 263608 115074 263664
rect 115074 263608 115124 263664
rect 115060 263604 115124 263608
rect 126836 263604 126900 263668
rect 263548 263060 263612 263124
rect 256740 262244 256804 262308
rect 255820 261836 255884 261900
rect 61884 261428 61948 261492
rect 252876 261700 252940 261764
rect 259684 260884 259748 260948
rect 255268 259932 255332 259996
rect 57652 259388 57716 259452
rect 59124 259388 59188 259452
rect 57652 258164 57716 258228
rect 124444 258028 124508 258092
rect 254532 258164 254596 258228
rect 258396 256804 258460 256868
rect 262260 256668 262324 256732
rect 106044 256320 106108 256324
rect 106044 256264 106094 256320
rect 106094 256264 106108 256320
rect 106044 256260 106108 256264
rect 258396 256048 258460 256052
rect 258396 255992 258410 256048
rect 258410 255992 258460 256048
rect 258396 255988 258460 255992
rect 258396 255308 258460 255372
rect 41276 254492 41340 254556
rect 57836 253948 57900 254012
rect 100708 253268 100772 253332
rect 59124 251228 59188 251292
rect 66116 249868 66180 249932
rect 108252 249052 108316 249116
rect 99236 248236 99300 248300
rect 192340 247556 192404 247620
rect 109540 247012 109604 247076
rect 66668 246196 66732 246260
rect 111012 246196 111076 246260
rect 111196 246060 111260 246124
rect 193444 246196 193508 246260
rect 108252 244836 108316 244900
rect 191052 244836 191116 244900
rect 253612 244700 253676 244764
rect 255268 244700 255332 244764
rect 255268 244428 255332 244492
rect 124260 244352 124324 244356
rect 124260 244296 124310 244352
rect 124310 244296 124324 244352
rect 124260 244292 124324 244296
rect 259500 244292 259564 244356
rect 100892 243476 100956 243540
rect 255820 243068 255884 243132
rect 66116 242932 66180 242996
rect 66668 242932 66732 242996
rect 191236 242932 191300 242996
rect 65932 241708 65996 241772
rect 61700 241572 61764 241636
rect 70164 241768 70228 241772
rect 70164 241712 70178 241768
rect 70178 241712 70228 241768
rect 70164 241708 70228 241712
rect 70900 241708 70964 241772
rect 71452 241708 71516 241772
rect 72924 241708 72988 241772
rect 74212 241768 74276 241772
rect 74212 241712 74262 241768
rect 74262 241712 74276 241768
rect 74212 241708 74276 241712
rect 91508 241768 91572 241772
rect 91508 241712 91558 241768
rect 91558 241712 91572 241768
rect 91508 241708 91572 241712
rect 102732 241708 102796 241772
rect 95004 241632 95068 241636
rect 95004 241576 95018 241632
rect 95018 241576 95068 241632
rect 95004 241572 95068 241576
rect 67772 241436 67836 241500
rect 107700 241436 107764 241500
rect 253980 241436 254044 241500
rect 253612 241164 253676 241228
rect 253612 240756 253676 240820
rect 69796 240076 69860 240140
rect 220860 240136 220924 240140
rect 220860 240080 220874 240136
rect 220874 240080 220924 240136
rect 55076 239940 55140 240004
rect 207060 239940 207124 240004
rect 220860 240076 220924 240080
rect 234660 240136 234724 240140
rect 234660 240080 234710 240136
rect 234710 240080 234724 240136
rect 234660 240076 234724 240080
rect 192708 239804 192772 239868
rect 252508 239532 252572 239596
rect 193812 238444 193876 238508
rect 238892 238308 238956 238372
rect 102732 238036 102796 238100
rect 118740 238036 118804 238100
rect 255268 237900 255332 237964
rect 242020 237356 242084 237420
rect 255268 237356 255332 237420
rect 111196 237220 111260 237284
rect 253612 237220 253676 237284
rect 111564 236676 111628 236740
rect 96660 235452 96724 235516
rect 118740 235452 118804 235516
rect 192340 235724 192404 235788
rect 191236 235180 191300 235244
rect 255820 234636 255884 234700
rect 114508 234500 114572 234564
rect 262260 234500 262324 234564
rect 118004 234364 118068 234428
rect 73108 233820 73172 233884
rect 100892 233820 100956 233884
rect 106780 232732 106844 232796
rect 121684 232732 121748 232796
rect 256740 233140 256804 233204
rect 93900 231236 93964 231300
rect 111748 231236 111812 231300
rect 116532 231780 116596 231844
rect 258396 231780 258460 231844
rect 61884 230420 61948 230484
rect 99972 230284 100036 230348
rect 100708 229740 100772 229804
rect 238708 229120 238772 229124
rect 238708 229064 238722 229120
rect 238722 229064 238772 229120
rect 238708 229060 238772 229064
rect 103836 228788 103900 228852
rect 238708 228848 238772 228852
rect 238708 228792 238722 228848
rect 238722 228792 238772 228848
rect 238708 228788 238772 228792
rect 214420 228244 214484 228308
rect 95188 227020 95252 227084
rect 259684 226884 259748 226948
rect 115980 226068 116044 226132
rect 104940 225932 105004 225996
rect 216812 225524 216876 225588
rect 110644 224164 110708 224228
rect 216076 224164 216140 224228
rect 186820 222804 186884 222868
rect 57652 222184 57716 222188
rect 57652 222128 57666 222184
rect 57666 222128 57716 222184
rect 57652 222124 57716 222128
rect 126836 222048 126900 222052
rect 126836 221992 126886 222048
rect 126886 221992 126900 222048
rect 126836 221988 126900 221992
rect 258396 221988 258460 222052
rect 93716 220628 93780 220692
rect 106412 220628 106476 220692
rect 121684 220220 121748 220284
rect 263732 220628 263796 220692
rect 117084 220084 117148 220148
rect 234844 220084 234908 220148
rect 238892 219404 238956 219468
rect 69980 219268 70044 219332
rect 238892 218996 238956 219060
rect 244412 217228 244476 217292
rect 244412 216684 244476 216748
rect 236500 215868 236564 215932
rect 133828 215188 133892 215252
rect 221228 214508 221292 214572
rect 108252 211924 108316 211988
rect 114508 211788 114572 211852
rect 128676 211848 128740 211852
rect 128676 211792 128690 211848
rect 128690 211792 128740 211848
rect 128676 211788 128740 211792
rect 104020 210292 104084 210356
rect 238708 209808 238772 209812
rect 238708 209752 238722 209808
rect 238722 209752 238772 209808
rect 238708 209748 238772 209752
rect 255820 209612 255884 209676
rect 238892 209476 238956 209540
rect 259500 206756 259564 206820
rect 92980 204172 93044 204236
rect 93716 204172 93780 204236
rect 218652 202812 218716 202876
rect 88196 202132 88260 202196
rect 103836 202132 103900 202196
rect 109540 200636 109604 200700
rect 205588 200636 205652 200700
rect 230980 200636 231044 200700
rect 238892 200092 238956 200156
rect 102732 199956 102796 200020
rect 254532 199956 254596 200020
rect 238892 199820 238956 199884
rect 67956 192476 68020 192540
rect 238708 190496 238772 190500
rect 238708 190440 238722 190496
rect 238722 190440 238772 190496
rect 238708 190436 238772 190440
rect 238708 190164 238772 190228
rect 219572 188260 219636 188324
rect 213684 186900 213748 186964
rect 198780 185540 198844 185604
rect 238708 180840 238772 180844
rect 238708 180784 238722 180840
rect 238722 180784 238772 180840
rect 238708 180780 238772 180784
rect 238708 180508 238772 180572
rect 238708 171184 238772 171188
rect 238708 171128 238722 171184
rect 238722 171128 238772 171184
rect 238708 171124 238772 171128
rect 238708 171048 238772 171052
rect 238708 170992 238722 171048
rect 238722 170992 238772 171048
rect 238708 170988 238772 170992
rect 238892 161468 238956 161532
rect 238708 161196 238772 161260
rect 203012 153716 203076 153780
rect 238708 151872 238772 151876
rect 238708 151816 238722 151872
rect 238722 151816 238772 151872
rect 238708 151812 238772 151816
rect 238708 151540 238772 151604
rect 197492 150996 197556 151060
rect 191052 149636 191116 149700
rect 122604 148276 122668 148340
rect 223804 146916 223868 146980
rect 239260 145556 239324 145620
rect 239260 138620 239324 138684
rect 68876 138076 68940 138140
rect 71084 136852 71148 136916
rect 88196 136716 88260 136780
rect 94084 135220 94148 135284
rect 71636 134736 71700 134740
rect 71636 134680 71686 134736
rect 71686 134680 71700 134736
rect 71636 134676 71700 134680
rect 67772 132772 67836 132836
rect 62988 130596 63052 130660
rect 106780 129916 106844 129980
rect 95188 124128 95252 124132
rect 95188 124072 95238 124128
rect 95238 124072 95252 124128
rect 95188 124068 95252 124072
rect 118740 118900 118804 118964
rect 98500 118628 98564 118692
rect 64644 116044 64708 116108
rect 114508 115092 114572 115156
rect 61884 113052 61948 113116
rect 66852 113052 66916 113116
rect 66852 111556 66916 111620
rect 97212 108292 97276 108356
rect 124444 106252 124508 106316
rect 233372 104076 233436 104140
rect 97212 103396 97276 103460
rect 59124 102172 59188 102236
rect 238524 101356 238588 101420
rect 121684 99996 121748 100060
rect 108252 98500 108316 98564
rect 99052 97140 99116 97204
rect 232084 97140 232148 97204
rect 66116 95236 66180 95300
rect 232268 94420 232332 94484
rect 69980 92652 70044 92716
rect 70900 92652 70964 92716
rect 69612 92516 69676 92580
rect 92980 92380 93044 92444
rect 95188 92380 95252 92444
rect 68876 91020 68940 91084
rect 71636 90884 71700 90948
rect 94084 90748 94148 90812
rect 103836 89660 103900 89724
rect 93900 89524 93964 89588
rect 224908 88980 224972 89044
rect 211660 76468 211724 76532
rect 208900 73748 208964 73812
rect 229692 72388 229756 72452
rect 210372 71028 210436 71092
rect 226564 47500 226628 47564
rect 196020 39204 196084 39268
rect 223988 36484 224052 36548
rect 222332 35124 222396 35188
rect 219204 33764 219268 33828
rect 230428 30908 230492 30972
rect 237788 29548 237852 29612
rect 227668 28188 227732 28252
rect 226380 25468 226444 25532
rect 222700 24108 222764 24172
rect 204300 22612 204364 22676
rect 201540 21252 201604 21316
rect 208348 11596 208412 11660
rect 233188 8876 233252 8940
rect 213868 7516 213932 7580
rect 130332 4932 130396 4996
rect 215892 4796 215956 4860
rect 238524 3980 238588 4044
rect 99052 3572 99116 3636
rect 117084 3572 117148 3636
rect 111564 3436 111628 3500
rect 240364 3436 240428 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41275 407012 41341 407013
rect 41275 406948 41276 407012
rect 41340 406948 41341 407012
rect 41275 406947 41341 406948
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 41278 254557 41338 406947
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41275 254556 41341 254557
rect 41275 254492 41276 254556
rect 41340 254492 41341 254556
rect 41275 254491 41341 254492
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55075 386476 55141 386477
rect 55075 386412 55076 386476
rect 55140 386412 55141 386476
rect 55075 386411 55141 386412
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 52315 305012 52381 305013
rect 52315 304948 52316 305012
rect 52380 304948 52381 305012
rect 52315 304947 52381 304948
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 52318 276181 52378 304947
rect 52315 276180 52381 276181
rect 52315 276116 52316 276180
rect 52380 276116 52381 276180
rect 52315 276115 52381 276116
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 55078 240005 55138 386411
rect 55794 381454 56414 416898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 583166 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 583166 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 75867 584900 75933 584901
rect 75867 584836 75868 584900
rect 75932 584836 75933 584900
rect 75867 584835 75933 584836
rect 75683 581092 75749 581093
rect 75683 581028 75684 581092
rect 75748 581028 75749 581092
rect 75683 581027 75749 581028
rect 70899 580820 70965 580821
rect 70899 580756 70900 580820
rect 70964 580756 70965 580820
rect 70899 580755 70965 580756
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 67771 548316 67837 548317
rect 67771 548252 67772 548316
rect 67836 548252 67837 548316
rect 67771 548251 67837 548252
rect 67774 539885 67834 548251
rect 69427 542196 69493 542197
rect 69427 542132 69428 542196
rect 69492 542132 69493 542196
rect 69427 542131 69493 542132
rect 67771 539884 67837 539885
rect 67771 539820 67772 539884
rect 67836 539820 67837 539884
rect 67771 539819 67837 539820
rect 69430 538230 69490 542131
rect 69430 538170 69674 538230
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 61883 425236 61949 425237
rect 61883 425172 61884 425236
rect 61948 425172 61949 425236
rect 61883 425171 61949 425172
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59123 411364 59189 411365
rect 59123 411300 59124 411364
rect 59188 411300 59189 411364
rect 59123 411299 59189 411300
rect 57835 407012 57901 407013
rect 57835 406948 57836 407012
rect 57900 406948 57901 407012
rect 57835 406947 57901 406948
rect 57838 405789 57898 406947
rect 57835 405788 57901 405789
rect 57835 405724 57836 405788
rect 57900 405724 57901 405788
rect 57835 405723 57901 405724
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55075 240004 55141 240005
rect 55075 239940 55076 240004
rect 55140 239940 55141 240004
rect 55075 239939 55141 239940
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 237454 56414 272898
rect 57651 259452 57717 259453
rect 57651 259388 57652 259452
rect 57716 259388 57717 259452
rect 57651 259387 57717 259388
rect 57654 258229 57714 259387
rect 57651 258228 57717 258229
rect 57651 258164 57652 258228
rect 57716 258164 57717 258228
rect 57651 258163 57717 258164
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 57654 222189 57714 258163
rect 57838 254013 57898 405723
rect 59126 259453 59186 411299
rect 59514 385174 60134 420618
rect 61699 387564 61765 387565
rect 61699 387500 61700 387564
rect 61764 387500 61765 387564
rect 61699 387499 61765 387500
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59123 259452 59189 259453
rect 59123 259388 59124 259452
rect 59188 259388 59189 259452
rect 59123 259387 59189 259388
rect 57835 254012 57901 254013
rect 57835 253948 57836 254012
rect 57900 253948 57901 254012
rect 57835 253947 57901 253948
rect 59123 251292 59189 251293
rect 59123 251228 59124 251292
rect 59188 251228 59189 251292
rect 59123 251227 59189 251228
rect 57651 222188 57717 222189
rect 57651 222124 57652 222188
rect 57716 222124 57717 222188
rect 57651 222123 57717 222124
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 59126 102237 59186 251227
rect 59514 241174 60134 276618
rect 61702 241637 61762 387499
rect 61886 296853 61946 425171
rect 63234 424894 63854 460338
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66115 443596 66181 443597
rect 66115 443532 66116 443596
rect 66180 443532 66181 443596
rect 66115 443531 66181 443532
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66118 408917 66178 443531
rect 66954 436356 67574 464058
rect 69614 462909 69674 538170
rect 69611 462908 69677 462909
rect 69611 462844 69612 462908
rect 69676 462844 69677 462908
rect 69611 462843 69677 462844
rect 69611 461548 69677 461549
rect 69611 461484 69612 461548
rect 69676 461484 69677 461548
rect 69611 461483 69677 461484
rect 67403 433260 67469 433261
rect 67403 433196 67404 433260
rect 67468 433196 67469 433260
rect 67403 433195 67469 433196
rect 66851 422244 66917 422245
rect 66851 422180 66852 422244
rect 66916 422180 66917 422244
rect 66851 422179 66917 422180
rect 66854 420205 66914 422179
rect 66851 420204 66917 420205
rect 66851 420140 66852 420204
rect 66916 420140 66917 420204
rect 66851 420139 66917 420140
rect 67406 409733 67466 433195
rect 67403 409732 67469 409733
rect 67403 409668 67404 409732
rect 67468 409668 67469 409732
rect 67403 409667 67469 409668
rect 66115 408916 66181 408917
rect 66115 408852 66116 408916
rect 66180 408852 66181 408916
rect 66115 408851 66181 408852
rect 69614 402990 69674 461483
rect 70163 434756 70229 434757
rect 70163 434692 70164 434756
rect 70228 434692 70229 434756
rect 70163 434691 70229 434692
rect 69430 402930 69674 402990
rect 69430 397765 69490 402930
rect 69427 397764 69493 397765
rect 69427 397700 69428 397764
rect 69492 397700 69493 397764
rect 69427 397699 69493 397700
rect 69611 392188 69677 392189
rect 69611 392124 69612 392188
rect 69676 392124 69677 392188
rect 69611 392123 69677 392124
rect 69614 388925 69674 392123
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 69611 388924 69677 388925
rect 69611 388860 69612 388924
rect 69676 388860 69677 388924
rect 69611 388859 69677 388860
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 66954 356614 67574 388356
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66115 334116 66181 334117
rect 66115 334052 66116 334116
rect 66180 334052 66181 334116
rect 66115 334051 66181 334052
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 61883 296852 61949 296853
rect 61883 296788 61884 296852
rect 61948 296788 61949 296852
rect 61883 296787 61949 296788
rect 61886 269245 61946 296787
rect 62987 282164 63053 282165
rect 62987 282100 62988 282164
rect 63052 282100 63053 282164
rect 62987 282099 63053 282100
rect 61883 269244 61949 269245
rect 61883 269180 61884 269244
rect 61948 269180 61949 269244
rect 61883 269179 61949 269180
rect 61883 261492 61949 261493
rect 61883 261428 61884 261492
rect 61948 261428 61949 261492
rect 61883 261427 61949 261428
rect 61699 241636 61765 241637
rect 61699 241572 61700 241636
rect 61764 241572 61765 241636
rect 61699 241571 61765 241572
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 61886 230485 61946 261427
rect 61883 230484 61949 230485
rect 61883 230420 61884 230484
rect 61948 230420 61949 230484
rect 61883 230419 61949 230420
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59123 102236 59189 102237
rect 59123 102172 59124 102236
rect 59188 102172 59189 102236
rect 59123 102171 59189 102172
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 97174 60134 132618
rect 61886 113117 61946 230419
rect 62990 130661 63050 282099
rect 63234 280894 63854 316338
rect 65931 283252 65997 283253
rect 65931 283188 65932 283252
rect 65996 283188 65997 283252
rect 65931 283187 65997 283188
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 64643 266524 64709 266525
rect 64643 266460 64644 266524
rect 64708 266460 64709 266524
rect 64643 266459 64709 266460
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 62987 130660 63053 130661
rect 62987 130596 62988 130660
rect 63052 130596 63053 130660
rect 62987 130595 63053 130596
rect 61883 113116 61949 113117
rect 61883 113052 61884 113116
rect 61948 113052 61949 113116
rect 61883 113051 61949 113052
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 100894 63854 136338
rect 64646 116109 64706 266459
rect 65934 241773 65994 283187
rect 66118 249933 66178 334051
rect 66954 320614 67574 356058
rect 70166 338061 70226 434691
rect 70902 433805 70962 580755
rect 73679 543454 73999 543486
rect 73679 543218 73721 543454
rect 73957 543218 73999 543454
rect 73679 543134 73999 543218
rect 73679 542898 73721 543134
rect 73957 542898 73999 543134
rect 73679 542866 73999 542898
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 72555 454748 72621 454749
rect 72555 454684 72556 454748
rect 72620 454684 72621 454748
rect 72555 454683 72621 454684
rect 71635 435436 71701 435437
rect 71635 435372 71636 435436
rect 71700 435372 71701 435436
rect 71635 435371 71701 435372
rect 70899 433804 70965 433805
rect 70899 433740 70900 433804
rect 70964 433740 70965 433804
rect 70899 433739 70965 433740
rect 70163 338060 70229 338061
rect 70163 337996 70164 338060
rect 70228 337996 70229 338060
rect 70163 337995 70229 337996
rect 71451 328540 71517 328541
rect 71451 328476 71452 328540
rect 71516 328476 71517 328540
rect 71451 328475 71517 328476
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 285592 67574 320058
rect 67771 296988 67837 296989
rect 67771 296924 67772 296988
rect 67836 296924 67837 296988
rect 67771 296923 67837 296924
rect 67774 275909 67834 296923
rect 70163 288420 70229 288421
rect 70163 288356 70164 288420
rect 70228 288356 70229 288420
rect 70163 288355 70229 288356
rect 70166 287197 70226 288355
rect 70163 287196 70229 287197
rect 70163 287132 70164 287196
rect 70228 287132 70229 287196
rect 70163 287131 70229 287132
rect 67955 280532 68021 280533
rect 67955 280468 67956 280532
rect 68020 280468 68021 280532
rect 67955 280467 68021 280468
rect 67771 275908 67837 275909
rect 67771 275844 67772 275908
rect 67836 275844 67837 275908
rect 67771 275843 67837 275844
rect 67774 274821 67834 275843
rect 67771 274820 67837 274821
rect 67771 274756 67772 274820
rect 67836 274756 67837 274820
rect 67771 274755 67837 274756
rect 66115 249932 66181 249933
rect 66115 249868 66116 249932
rect 66180 249868 66181 249932
rect 66115 249867 66181 249868
rect 66667 246260 66733 246261
rect 66667 246196 66668 246260
rect 66732 246196 66733 246260
rect 66667 246195 66733 246196
rect 66670 242997 66730 246195
rect 66115 242996 66181 242997
rect 66115 242932 66116 242996
rect 66180 242932 66181 242996
rect 66115 242931 66181 242932
rect 66667 242996 66733 242997
rect 66667 242932 66668 242996
rect 66732 242932 66733 242996
rect 66667 242931 66733 242932
rect 65931 241772 65997 241773
rect 65931 241708 65932 241772
rect 65996 241708 65997 241772
rect 65931 241707 65997 241708
rect 64643 116108 64709 116109
rect 64643 116044 64644 116108
rect 64708 116044 64709 116108
rect 64643 116043 64709 116044
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 66118 95301 66178 242931
rect 67771 241500 67837 241501
rect 67771 241436 67772 241500
rect 67836 241436 67837 241500
rect 67771 241435 67837 241436
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 136782 67574 140058
rect 67774 132837 67834 241435
rect 67958 192541 68018 280467
rect 70166 241773 70226 287131
rect 71083 283524 71149 283525
rect 71083 283460 71084 283524
rect 71148 283460 71149 283524
rect 71083 283459 71149 283460
rect 70163 241772 70229 241773
rect 70163 241770 70164 241772
rect 69614 241710 70164 241770
rect 67955 192540 68021 192541
rect 67955 192476 67956 192540
rect 68020 192476 68021 192540
rect 67955 192475 68021 192476
rect 68875 138140 68941 138141
rect 68875 138076 68876 138140
rect 68940 138076 68941 138140
rect 68875 138075 68941 138076
rect 67771 132836 67837 132837
rect 67771 132772 67772 132836
rect 67836 132772 67837 132836
rect 67771 132771 67837 132772
rect 66851 113116 66917 113117
rect 66851 113052 66852 113116
rect 66916 113052 66917 113116
rect 66851 113051 66917 113052
rect 66854 111621 66914 113051
rect 66851 111620 66917 111621
rect 66851 111556 66852 111620
rect 66916 111556 66917 111620
rect 66851 111555 66917 111556
rect 66115 95300 66181 95301
rect 66115 95236 66116 95300
rect 66180 95236 66181 95300
rect 66115 95235 66181 95236
rect 68878 91085 68938 138075
rect 69614 92581 69674 241710
rect 70163 241708 70164 241710
rect 70228 241708 70229 241772
rect 70163 241707 70229 241708
rect 70899 241772 70965 241773
rect 70899 241708 70900 241772
rect 70964 241708 70965 241772
rect 70899 241707 70965 241708
rect 69795 240140 69861 240141
rect 69795 240076 69796 240140
rect 69860 240076 69861 240140
rect 69795 240075 69861 240076
rect 69798 229110 69858 240075
rect 69798 229050 70042 229110
rect 69982 219333 70042 229050
rect 69979 219332 70045 219333
rect 69979 219268 69980 219332
rect 70044 219268 70045 219332
rect 69979 219267 70045 219268
rect 69982 92717 70042 219267
rect 70902 92717 70962 241707
rect 71086 136917 71146 283459
rect 71454 241773 71514 328475
rect 71638 287061 71698 435371
rect 72558 390421 72618 454683
rect 73794 436356 74414 470898
rect 75686 468485 75746 581027
rect 75870 535533 75930 584835
rect 77514 583166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 583166 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 583166 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 583166 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 583166 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 78443 581092 78509 581093
rect 78443 581028 78444 581092
rect 78508 581028 78509 581092
rect 78443 581027 78509 581028
rect 77644 561454 77964 561486
rect 77644 561218 77686 561454
rect 77922 561218 77964 561454
rect 77644 561134 77964 561218
rect 77644 560898 77686 561134
rect 77922 560898 77964 561134
rect 77644 560866 77964 560898
rect 75867 535532 75933 535533
rect 75867 535468 75868 535532
rect 75932 535468 75933 535532
rect 75867 535467 75933 535468
rect 77155 518124 77221 518125
rect 77155 518060 77156 518124
rect 77220 518060 77221 518124
rect 77155 518059 77221 518060
rect 75683 468484 75749 468485
rect 75683 468420 75684 468484
rect 75748 468420 75749 468484
rect 75683 468419 75749 468420
rect 72739 436252 72805 436253
rect 72739 436188 72740 436252
rect 72804 436188 72805 436252
rect 72739 436187 72805 436188
rect 72555 390420 72621 390421
rect 72555 390356 72556 390420
rect 72620 390356 72621 390420
rect 72555 390355 72621 390356
rect 71819 389060 71885 389061
rect 71819 388996 71820 389060
rect 71884 388996 71885 389060
rect 71819 388995 71885 388996
rect 71822 384301 71882 388995
rect 71819 384300 71885 384301
rect 71819 384236 71820 384300
rect 71884 384236 71885 384300
rect 71819 384235 71885 384236
rect 72742 318885 72802 436187
rect 73475 434892 73541 434893
rect 73475 434828 73476 434892
rect 73540 434828 73541 434892
rect 73475 434827 73541 434828
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 73478 343773 73538 434827
rect 75683 434756 75749 434757
rect 75683 434692 75684 434756
rect 75748 434692 75749 434756
rect 75683 434691 75749 434692
rect 74579 434348 74645 434349
rect 74579 434284 74580 434348
rect 74644 434284 74645 434348
rect 74579 434283 74645 434284
rect 73794 363454 74414 388356
rect 74582 380901 74642 434283
rect 74579 380900 74645 380901
rect 74579 380836 74580 380900
rect 74644 380836 74645 380900
rect 74579 380835 74645 380836
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73475 343772 73541 343773
rect 73475 343708 73476 343772
rect 73540 343708 73541 343772
rect 73475 343707 73541 343708
rect 72739 318884 72805 318885
rect 72739 318820 72740 318884
rect 72804 318820 72805 318884
rect 72739 318819 72805 318820
rect 72923 287740 72989 287741
rect 72923 287676 72924 287740
rect 72988 287676 72989 287740
rect 72923 287675 72989 287676
rect 71635 287060 71701 287061
rect 71635 286996 71636 287060
rect 71700 286996 71701 287060
rect 71635 286995 71701 286996
rect 71638 283797 71698 286995
rect 71635 283796 71701 283797
rect 71635 283732 71636 283796
rect 71700 283732 71701 283796
rect 71635 283731 71701 283732
rect 72926 241773 72986 287675
rect 73478 283525 73538 343707
rect 73794 327454 74414 362898
rect 75686 340917 75746 434691
rect 75867 434348 75933 434349
rect 75867 434284 75868 434348
rect 75932 434284 75933 434348
rect 75867 434283 75933 434284
rect 75870 385117 75930 434283
rect 77158 390421 77218 518059
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 78446 460189 78506 581027
rect 83963 580820 84029 580821
rect 83963 580756 83964 580820
rect 84028 580756 84029 580820
rect 83963 580755 84029 580756
rect 88379 580820 88445 580821
rect 88379 580756 88380 580820
rect 88444 580756 88445 580820
rect 88379 580755 88445 580756
rect 81609 543454 81929 543486
rect 81609 543218 81651 543454
rect 81887 543218 81929 543454
rect 81609 543134 81929 543218
rect 81609 542898 81651 543134
rect 81887 542898 81929 543134
rect 81609 542866 81929 542898
rect 79915 527780 79981 527781
rect 79915 527716 79916 527780
rect 79980 527716 79981 527780
rect 79915 527715 79981 527716
rect 78443 460188 78509 460189
rect 78443 460124 78444 460188
rect 78508 460124 78509 460188
rect 78443 460123 78509 460124
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 436356 78134 438618
rect 78259 436116 78325 436117
rect 78259 436052 78260 436116
rect 78324 436052 78325 436116
rect 78259 436051 78325 436052
rect 77155 390420 77221 390421
rect 77155 390356 77156 390420
rect 77220 390356 77221 390420
rect 77155 390355 77221 390356
rect 75867 385116 75933 385117
rect 75867 385052 75868 385116
rect 75932 385052 75933 385116
rect 75867 385051 75933 385052
rect 77514 367174 78134 388356
rect 78262 386341 78322 436051
rect 78443 433668 78509 433669
rect 78443 433604 78444 433668
rect 78508 433604 78509 433668
rect 78443 433603 78509 433604
rect 79731 433668 79797 433669
rect 79731 433604 79732 433668
rect 79796 433604 79797 433668
rect 79731 433603 79797 433604
rect 78446 390693 78506 433603
rect 78443 390692 78509 390693
rect 78443 390628 78444 390692
rect 78508 390628 78509 390692
rect 78443 390627 78509 390628
rect 78259 386340 78325 386341
rect 78259 386276 78260 386340
rect 78324 386276 78325 386340
rect 78259 386275 78325 386276
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 75683 340916 75749 340917
rect 75683 340852 75684 340916
rect 75748 340852 75749 340916
rect 75683 340851 75749 340852
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 285592 74414 290898
rect 77514 331174 78134 366618
rect 79734 335370 79794 433603
rect 79918 389061 79978 527715
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 436356 81854 442338
rect 83966 435981 84026 580755
rect 85575 561454 85895 561486
rect 85575 561218 85617 561454
rect 85853 561218 85895 561454
rect 85575 561134 85895 561218
rect 85575 560898 85617 561134
rect 85853 560898 85895 561134
rect 85575 560866 85895 560898
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 436356 85574 446058
rect 88382 444957 88442 580755
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 97211 554164 97277 554165
rect 97211 554100 97212 554164
rect 97276 554100 97277 554164
rect 97211 554099 97277 554100
rect 96659 547092 96725 547093
rect 96659 547028 96660 547092
rect 96724 547028 96725 547092
rect 96659 547027 96725 547028
rect 89540 543454 89860 543486
rect 89540 543218 89582 543454
rect 89818 543218 89860 543454
rect 89540 543134 89860 543218
rect 89540 542898 89582 543134
rect 89818 542898 89860 543134
rect 89540 542866 89860 542898
rect 94083 541652 94149 541653
rect 94083 541588 94084 541652
rect 94148 541588 94149 541652
rect 94083 541587 94149 541588
rect 91507 538252 91573 538253
rect 91507 538188 91508 538252
rect 91572 538188 91573 538252
rect 91507 538187 91573 538188
rect 88747 462908 88813 462909
rect 88747 462844 88748 462908
rect 88812 462844 88813 462908
rect 88747 462843 88813 462844
rect 88379 444956 88445 444957
rect 88379 444892 88380 444956
rect 88444 444892 88445 444956
rect 88379 444891 88445 444892
rect 86171 436252 86237 436253
rect 86171 436188 86172 436252
rect 86236 436188 86237 436252
rect 86171 436187 86237 436188
rect 82123 435980 82189 435981
rect 82123 435916 82124 435980
rect 82188 435916 82189 435980
rect 82123 435915 82189 435916
rect 83963 435980 84029 435981
rect 83963 435916 83964 435980
rect 84028 435916 84029 435980
rect 83963 435915 84029 435916
rect 80283 434348 80349 434349
rect 80283 434284 80284 434348
rect 80348 434284 80349 434348
rect 80283 434283 80349 434284
rect 80651 434348 80717 434349
rect 80651 434284 80652 434348
rect 80716 434284 80717 434348
rect 80651 434283 80717 434284
rect 81939 434348 82005 434349
rect 81939 434284 81940 434348
rect 82004 434284 82005 434348
rect 81939 434283 82005 434284
rect 79915 389060 79981 389061
rect 79915 388996 79916 389060
rect 79980 388996 79981 389060
rect 79915 388995 79981 388996
rect 80286 384437 80346 434283
rect 80654 387973 80714 434283
rect 80651 387972 80717 387973
rect 80651 387908 80652 387972
rect 80716 387908 80717 387972
rect 80651 387907 80717 387908
rect 80283 384436 80349 384437
rect 80283 384372 80284 384436
rect 80348 384372 80349 384436
rect 80283 384371 80349 384372
rect 79182 335310 79794 335370
rect 81234 370894 81854 388356
rect 81942 379541 82002 434283
rect 82126 391101 82186 435915
rect 85435 434756 85501 434757
rect 85435 434692 85436 434756
rect 85500 434692 85501 434756
rect 85435 434691 85501 434692
rect 83411 434620 83477 434621
rect 83411 434556 83412 434620
rect 83476 434556 83477 434620
rect 83411 434555 83477 434556
rect 82123 391100 82189 391101
rect 82123 391036 82124 391100
rect 82188 391036 82189 391100
rect 82123 391035 82189 391036
rect 81939 379540 82005 379541
rect 81939 379476 81940 379540
rect 82004 379476 82005 379540
rect 81939 379475 82005 379476
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 79182 332621 79242 335310
rect 81234 334894 81854 370338
rect 82859 339556 82925 339557
rect 82859 339492 82860 339556
rect 82924 339492 82925 339556
rect 82859 339491 82925 339492
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 79179 332620 79245 332621
rect 79179 332556 79180 332620
rect 79244 332556 79245 332620
rect 79179 332555 79245 332556
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 79182 319429 79242 332555
rect 79179 319428 79245 319429
rect 79179 319364 79180 319428
rect 79244 319364 79245 319428
rect 79179 319363 79245 319364
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285592 78134 294618
rect 81234 298894 81854 334338
rect 82862 322965 82922 339491
rect 82859 322964 82925 322965
rect 82859 322900 82860 322964
rect 82924 322900 82925 322964
rect 82859 322899 82925 322900
rect 83414 318749 83474 434555
rect 83595 434484 83661 434485
rect 83595 434420 83596 434484
rect 83660 434420 83661 434484
rect 83595 434419 83661 434420
rect 83598 339557 83658 434419
rect 84699 433804 84765 433805
rect 84699 433740 84700 433804
rect 84764 433740 84765 433804
rect 84699 433739 84765 433740
rect 84702 385117 84762 433739
rect 85438 391101 85498 434691
rect 85803 434348 85869 434349
rect 85803 434284 85804 434348
rect 85868 434284 85869 434348
rect 85803 434283 85869 434284
rect 85435 391100 85501 391101
rect 85435 391036 85436 391100
rect 85500 391036 85501 391100
rect 85435 391035 85501 391036
rect 84699 385116 84765 385117
rect 84699 385052 84700 385116
rect 84764 385052 84765 385116
rect 84699 385051 84765 385052
rect 84954 374614 85574 388356
rect 85806 383757 85866 434283
rect 86174 387701 86234 436187
rect 87091 434348 87157 434349
rect 87091 434284 87092 434348
rect 87156 434284 87157 434348
rect 87091 434283 87157 434284
rect 86171 387700 86237 387701
rect 86171 387636 86172 387700
rect 86236 387636 86237 387700
rect 86171 387635 86237 387636
rect 85803 383756 85869 383757
rect 85803 383692 85804 383756
rect 85868 383692 85869 383756
rect 85803 383691 85869 383692
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 83595 339556 83661 339557
rect 83595 339492 83596 339556
rect 83660 339492 83661 339556
rect 83595 339491 83661 339492
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 83411 318748 83477 318749
rect 83411 318684 83412 318748
rect 83476 318684 83477 318748
rect 83411 318683 83477 318684
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 285592 81854 298338
rect 84954 302614 85574 338058
rect 87094 329085 87154 434283
rect 87275 433668 87341 433669
rect 87275 433604 87276 433668
rect 87340 433604 87341 433668
rect 87275 433603 87341 433604
rect 87091 329084 87157 329085
rect 87091 329020 87092 329084
rect 87156 329020 87157 329084
rect 87091 329019 87157 329020
rect 87278 304197 87338 433603
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 88750 391101 88810 462843
rect 90955 434892 91021 434893
rect 90955 434828 90956 434892
rect 91020 434828 91021 434892
rect 90955 434827 91021 434828
rect 89667 433668 89733 433669
rect 89667 433604 89668 433668
rect 89732 433604 89733 433668
rect 89667 433603 89733 433604
rect 89670 398850 89730 433603
rect 89670 398790 89914 398850
rect 88747 391100 88813 391101
rect 88747 391036 88748 391100
rect 88812 391036 88813 391100
rect 88747 391035 88813 391036
rect 89854 389190 89914 398790
rect 89670 389130 89914 389190
rect 89670 377365 89730 389130
rect 89667 377364 89733 377365
rect 89667 377300 89668 377364
rect 89732 377300 89733 377364
rect 89667 377299 89733 377300
rect 87275 304196 87341 304197
rect 87275 304132 87276 304196
rect 87340 304132 87341 304196
rect 87275 304131 87341 304132
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 285592 85574 302058
rect 90958 292637 91018 434827
rect 91323 433668 91389 433669
rect 91323 433604 91324 433668
rect 91388 433604 91389 433668
rect 91323 433603 91389 433604
rect 91326 333301 91386 433603
rect 91510 389061 91570 538187
rect 91794 525454 92414 537166
rect 94086 531997 94146 541587
rect 94083 531996 94149 531997
rect 94083 531932 94084 531996
rect 94148 531932 94149 531996
rect 94083 531931 94149 531932
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 95514 529174 96134 537166
rect 96662 533357 96722 547027
rect 96659 533356 96725 533357
rect 96659 533292 96660 533356
rect 96724 533292 96725 533356
rect 96659 533291 96725 533292
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 94451 520980 94517 520981
rect 94451 520916 94452 520980
rect 94516 520916 94517 520980
rect 94451 520915 94517 520916
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 92611 460188 92677 460189
rect 92611 460124 92612 460188
rect 92676 460124 92677 460188
rect 92611 460123 92677 460124
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 436356 92414 452898
rect 92614 391101 92674 460123
rect 93899 434348 93965 434349
rect 93899 434284 93900 434348
rect 93964 434284 93965 434348
rect 93899 434283 93965 434284
rect 93715 433668 93781 433669
rect 93715 433604 93716 433668
rect 93780 433604 93781 433668
rect 93715 433603 93781 433604
rect 92611 391100 92677 391101
rect 92611 391036 92612 391100
rect 92676 391036 92677 391100
rect 92611 391035 92677 391036
rect 91507 389060 91573 389061
rect 91507 388996 91508 389060
rect 91572 388996 91573 389060
rect 91507 388995 91573 388996
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91323 333300 91389 333301
rect 91323 333236 91324 333300
rect 91388 333236 91389 333300
rect 91323 333235 91389 333236
rect 91507 332756 91573 332757
rect 91507 332692 91508 332756
rect 91572 332692 91573 332756
rect 91507 332691 91573 332692
rect 90955 292636 91021 292637
rect 90955 292572 90956 292636
rect 91020 292572 91021 292636
rect 90955 292571 91021 292572
rect 74211 284204 74277 284205
rect 74211 284140 74212 284204
rect 74276 284140 74277 284204
rect 74211 284139 74277 284140
rect 73475 283524 73541 283525
rect 73475 283460 73476 283524
rect 73540 283460 73541 283524
rect 73475 283459 73541 283460
rect 73478 282930 73538 283459
rect 73110 282870 73538 282930
rect 71451 241772 71517 241773
rect 71451 241708 71452 241772
rect 71516 241708 71517 241772
rect 71451 241707 71517 241708
rect 72923 241772 72989 241773
rect 72923 241708 72924 241772
rect 72988 241708 72989 241772
rect 72923 241707 72989 241708
rect 73110 233885 73170 282870
rect 74214 241773 74274 284139
rect 78977 273454 79297 273486
rect 78977 273218 79019 273454
rect 79255 273218 79297 273454
rect 78977 273134 79297 273218
rect 78977 272898 79019 273134
rect 79255 272898 79297 273134
rect 78977 272866 79297 272898
rect 88241 273454 88561 273486
rect 88241 273218 88283 273454
rect 88519 273218 88561 273454
rect 88241 273134 88561 273218
rect 88241 272898 88283 273134
rect 88519 272898 88561 273134
rect 88241 272866 88561 272898
rect 74345 255454 74665 255486
rect 74345 255218 74387 255454
rect 74623 255218 74665 255454
rect 74345 255134 74665 255218
rect 74345 254898 74387 255134
rect 74623 254898 74665 255134
rect 74345 254866 74665 254898
rect 83609 255454 83929 255486
rect 83609 255218 83651 255454
rect 83887 255218 83929 255454
rect 83609 255134 83929 255218
rect 83609 254898 83651 255134
rect 83887 254898 83929 255134
rect 83609 254866 83929 254898
rect 91510 241773 91570 332691
rect 91794 309454 92414 344898
rect 93718 332757 93778 433603
rect 93902 378725 93962 434283
rect 94454 389061 94514 520915
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 436356 96134 456618
rect 97214 444277 97274 554099
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 111747 583812 111813 583813
rect 111747 583748 111748 583812
rect 111812 583748 111813 583812
rect 111747 583747 111813 583748
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 104939 547908 105005 547909
rect 104939 547844 104940 547908
rect 105004 547844 105005 547908
rect 104939 547843 105005 547844
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 100707 507924 100773 507925
rect 100707 507860 100708 507924
rect 100772 507860 100773 507924
rect 100707 507859 100773 507860
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 97211 444276 97277 444277
rect 97211 444212 97212 444276
rect 97276 444212 97277 444276
rect 97211 444211 97277 444212
rect 99234 436356 99854 460338
rect 100523 436116 100589 436117
rect 100523 436052 100524 436116
rect 100588 436052 100589 436116
rect 100523 436051 100589 436052
rect 97211 434348 97277 434349
rect 97211 434284 97212 434348
rect 97276 434284 97277 434348
rect 97211 434283 97277 434284
rect 95187 433668 95253 433669
rect 95187 433604 95188 433668
rect 95252 433604 95253 433668
rect 95187 433603 95253 433604
rect 94451 389060 94517 389061
rect 94451 388996 94452 389060
rect 94516 388996 94517 389060
rect 94451 388995 94517 388996
rect 95190 380221 95250 433603
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95187 380220 95253 380221
rect 95187 380156 95188 380220
rect 95252 380156 95253 380220
rect 95187 380155 95253 380156
rect 93899 378724 93965 378725
rect 93899 378660 93900 378724
rect 93964 378660 93965 378724
rect 93899 378659 93965 378660
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 92979 332756 93045 332757
rect 92979 332692 92980 332756
rect 93044 332692 93045 332756
rect 92979 332691 93045 332692
rect 93715 332756 93781 332757
rect 93715 332692 93716 332756
rect 93780 332692 93781 332756
rect 93715 332691 93781 332692
rect 92982 323645 93042 332691
rect 95003 327044 95069 327045
rect 95003 326980 95004 327044
rect 95068 326980 95069 327044
rect 95003 326979 95069 326980
rect 92979 323644 93045 323645
rect 92979 323580 92980 323644
rect 93044 323580 93045 323644
rect 92979 323579 93045 323580
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 285592 92414 308898
rect 92873 255454 93193 255486
rect 92873 255218 92915 255454
rect 93151 255218 93193 255454
rect 92873 255134 93193 255218
rect 92873 254898 92915 255134
rect 93151 254898 93193 255134
rect 92873 254866 93193 254898
rect 74211 241772 74277 241773
rect 74211 241708 74212 241772
rect 74276 241708 74277 241772
rect 74211 241707 74277 241708
rect 91507 241772 91573 241773
rect 91507 241708 91508 241772
rect 91572 241708 91573 241772
rect 91507 241707 91573 241708
rect 95006 241637 95066 326979
rect 95514 313174 96134 348618
rect 97214 320925 97274 434283
rect 97395 433940 97461 433941
rect 97395 433876 97396 433940
rect 97460 433876 97461 433940
rect 97395 433875 97461 433876
rect 97398 385661 97458 433875
rect 98131 433804 98197 433805
rect 98131 433740 98132 433804
rect 98196 433740 98197 433804
rect 98131 433739 98197 433740
rect 97395 385660 97461 385661
rect 97395 385596 97396 385660
rect 97460 385596 97461 385660
rect 97395 385595 97461 385596
rect 98134 373285 98194 433739
rect 98499 433668 98565 433669
rect 98499 433604 98500 433668
rect 98564 433604 98565 433668
rect 98499 433603 98565 433604
rect 99971 433668 100037 433669
rect 99971 433604 99972 433668
rect 100036 433604 100037 433668
rect 99971 433603 100037 433604
rect 98131 373284 98197 373285
rect 98131 373220 98132 373284
rect 98196 373220 98197 373284
rect 98131 373219 98197 373220
rect 98502 335370 98562 433603
rect 97950 335310 98562 335370
rect 99234 352894 99854 388356
rect 99974 387157 100034 433603
rect 100526 388517 100586 436051
rect 100710 390965 100770 507859
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 436356 103574 464058
rect 103283 436252 103349 436253
rect 103283 436188 103284 436252
rect 103348 436188 103349 436252
rect 103283 436187 103349 436188
rect 102179 434348 102245 434349
rect 102179 434284 102180 434348
rect 102244 434284 102245 434348
rect 102179 434283 102245 434284
rect 101995 433804 102061 433805
rect 101995 433740 101996 433804
rect 102060 433740 102061 433804
rect 101995 433739 102061 433740
rect 100707 390964 100773 390965
rect 100707 390900 100708 390964
rect 100772 390900 100773 390964
rect 100707 390899 100773 390900
rect 100523 388516 100589 388517
rect 100523 388452 100524 388516
rect 100588 388452 100589 388516
rect 100523 388451 100589 388452
rect 99971 387156 100037 387157
rect 99971 387092 99972 387156
rect 100036 387092 100037 387156
rect 99971 387091 100037 387092
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 97950 329901 98010 335310
rect 97947 329900 98013 329901
rect 97947 329836 97948 329900
rect 98012 329836 98013 329900
rect 97947 329835 98013 329836
rect 97211 320924 97277 320925
rect 97211 320860 97212 320924
rect 97276 320860 97277 320924
rect 97211 320859 97277 320860
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 285592 96134 312618
rect 97950 285429 98010 329835
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 285592 99854 316338
rect 100155 291412 100221 291413
rect 100155 291348 100156 291412
rect 100220 291348 100221 291412
rect 100155 291347 100221 291348
rect 97947 285428 98013 285429
rect 97947 285364 97948 285428
rect 98012 285364 98013 285428
rect 97947 285363 98013 285364
rect 95187 283524 95253 283525
rect 95187 283460 95188 283524
rect 95252 283460 95253 283524
rect 95187 283459 95253 283460
rect 96659 283524 96725 283525
rect 96659 283460 96660 283524
rect 96724 283460 96725 283524
rect 96659 283459 96725 283460
rect 95003 241636 95069 241637
rect 95003 241572 95004 241636
rect 95068 241572 95069 241636
rect 95003 241571 95069 241572
rect 73107 233884 73173 233885
rect 73107 233820 73108 233884
rect 73172 233820 73173 233884
rect 73107 233819 73173 233820
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 71083 136916 71149 136917
rect 71083 136852 71084 136916
rect 71148 136852 71149 136916
rect 71083 136851 71149 136852
rect 73794 136782 74414 146898
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 136782 78134 150618
rect 81234 226894 81854 239592
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 136782 81854 154338
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 88195 202196 88261 202197
rect 88195 202132 88196 202196
rect 88260 202132 88261 202196
rect 88195 202131 88261 202132
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 136782 85574 158058
rect 88198 136781 88258 202131
rect 91794 201454 92414 236898
rect 93899 231300 93965 231301
rect 93899 231236 93900 231300
rect 93964 231236 93965 231300
rect 93899 231235 93965 231236
rect 93715 220692 93781 220693
rect 93715 220628 93716 220692
rect 93780 220628 93781 220692
rect 93715 220627 93781 220628
rect 93718 204237 93778 220627
rect 92979 204236 93045 204237
rect 92979 204172 92980 204236
rect 93044 204172 93045 204236
rect 92979 204171 93045 204172
rect 93715 204236 93781 204237
rect 93715 204172 93716 204236
rect 93780 204172 93781 204236
rect 93715 204171 93781 204172
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 136782 92414 164898
rect 88195 136780 88261 136781
rect 88195 136716 88196 136780
rect 88260 136716 88261 136780
rect 88195 136715 88261 136716
rect 71635 134740 71701 134741
rect 71635 134676 71636 134740
rect 71700 134676 71701 134740
rect 71635 134675 71701 134676
rect 69979 92716 70045 92717
rect 69979 92652 69980 92716
rect 70044 92652 70045 92716
rect 69979 92651 70045 92652
rect 70899 92716 70965 92717
rect 70899 92652 70900 92716
rect 70964 92652 70965 92716
rect 70899 92651 70965 92652
rect 69611 92580 69677 92581
rect 69611 92516 69612 92580
rect 69676 92516 69677 92580
rect 69611 92515 69677 92516
rect 68875 91084 68941 91085
rect 68875 91020 68876 91084
rect 68940 91020 68941 91084
rect 68875 91019 68941 91020
rect 71638 90949 71698 134675
rect 77644 129454 77964 129486
rect 77644 129218 77686 129454
rect 77922 129218 77964 129454
rect 77644 129134 77964 129218
rect 77644 128898 77686 129134
rect 77922 128898 77964 129134
rect 77644 128866 77964 128898
rect 85575 129454 85895 129486
rect 85575 129218 85617 129454
rect 85853 129218 85895 129454
rect 85575 129134 85895 129218
rect 85575 128898 85617 129134
rect 85853 128898 85895 129134
rect 85575 128866 85895 128898
rect 73679 111454 73999 111486
rect 73679 111218 73721 111454
rect 73957 111218 73999 111454
rect 73679 111134 73999 111218
rect 73679 110898 73721 111134
rect 73957 110898 73999 111134
rect 73679 110866 73999 110898
rect 81609 111454 81929 111486
rect 81609 111218 81651 111454
rect 81887 111218 81929 111454
rect 81609 111134 81929 111218
rect 81609 110898 81651 111134
rect 81887 110898 81929 111134
rect 81609 110866 81929 110898
rect 89540 111454 89860 111486
rect 89540 111218 89582 111454
rect 89818 111218 89860 111454
rect 89540 111134 89860 111218
rect 89540 110898 89582 111134
rect 89818 110898 89860 111134
rect 89540 110866 89860 110898
rect 92982 92445 93042 204171
rect 92979 92444 93045 92445
rect 92979 92380 92980 92444
rect 93044 92380 93045 92444
rect 92979 92379 93045 92380
rect 71635 90948 71701 90949
rect 71635 90884 71636 90948
rect 71700 90884 71701 90948
rect 71635 90883 71701 90884
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 90782
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 90782
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 90782
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 90782
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 90782
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 90782
rect 93902 89589 93962 231235
rect 95190 227085 95250 283459
rect 95187 227084 95253 227085
rect 95187 227020 95188 227084
rect 95252 227020 95253 227084
rect 95187 227019 95253 227020
rect 95514 205174 96134 239592
rect 96662 235517 96722 283459
rect 97950 282930 98010 285363
rect 97950 282870 98562 282930
rect 98502 271149 98562 282870
rect 99971 282708 100037 282709
rect 99971 282644 99972 282708
rect 100036 282644 100037 282708
rect 99971 282643 100037 282644
rect 98499 271148 98565 271149
rect 98499 271084 98500 271148
rect 98564 271084 98565 271148
rect 98499 271083 98565 271084
rect 99235 266388 99301 266389
rect 99235 266324 99236 266388
rect 99300 266324 99301 266388
rect 99235 266323 99301 266324
rect 99238 248430 99298 266323
rect 98502 248370 99298 248430
rect 96659 235516 96725 235517
rect 96659 235452 96660 235516
rect 96724 235452 96725 235516
rect 96659 235451 96725 235452
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 136782 96134 168618
rect 94083 135284 94149 135285
rect 94083 135220 94084 135284
rect 94148 135220 94149 135284
rect 94083 135219 94149 135220
rect 94086 90813 94146 135219
rect 95187 124132 95253 124133
rect 95187 124068 95188 124132
rect 95252 124068 95253 124132
rect 95187 124067 95253 124068
rect 95190 92445 95250 124067
rect 98502 118693 98562 248370
rect 99238 248301 99298 248370
rect 99235 248300 99301 248301
rect 99235 248236 99236 248300
rect 99300 248236 99301 248300
rect 99235 248235 99301 248236
rect 99234 208894 99854 239592
rect 99974 230349 100034 282643
rect 100158 267341 100218 291347
rect 101998 282709 102058 433739
rect 102182 364989 102242 434283
rect 103286 388517 103346 436187
rect 104203 434348 104269 434349
rect 104203 434284 104204 434348
rect 104268 434284 104269 434348
rect 104203 434283 104269 434284
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 103283 388516 103349 388517
rect 103283 388452 103284 388516
rect 103348 388452 103349 388516
rect 103283 388451 103349 388452
rect 102179 364988 102245 364989
rect 102179 364924 102180 364988
rect 102244 364924 102245 364988
rect 102179 364923 102245 364924
rect 102954 356614 103574 388356
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102731 335476 102797 335477
rect 102731 335412 102732 335476
rect 102796 335412 102797 335476
rect 102731 335411 102797 335412
rect 101995 282708 102061 282709
rect 101995 282644 101996 282708
rect 102060 282644 102061 282708
rect 101995 282643 102061 282644
rect 100155 267340 100221 267341
rect 100155 267276 100156 267340
rect 100220 267276 100221 267340
rect 100155 267275 100221 267276
rect 100707 253332 100773 253333
rect 100707 253268 100708 253332
rect 100772 253268 100773 253332
rect 100707 253267 100773 253268
rect 99971 230348 100037 230349
rect 99971 230284 99972 230348
rect 100036 230284 100037 230348
rect 99971 230283 100037 230284
rect 100710 229805 100770 253267
rect 100891 243540 100957 243541
rect 100891 243476 100892 243540
rect 100956 243476 100957 243540
rect 100891 243475 100957 243476
rect 100894 233885 100954 243475
rect 102734 241773 102794 335411
rect 102954 320614 103574 356058
rect 104206 322149 104266 434283
rect 104942 390421 105002 547843
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 106411 463044 106477 463045
rect 106411 462980 106412 463044
rect 106476 462980 106477 463044
rect 106411 462979 106477 462980
rect 105123 433668 105189 433669
rect 105123 433604 105124 433668
rect 105188 433604 105189 433668
rect 105123 433603 105189 433604
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 105126 387021 105186 433603
rect 106414 390421 106474 462979
rect 107699 449172 107765 449173
rect 107699 449108 107700 449172
rect 107764 449108 107765 449172
rect 107699 449107 107765 449108
rect 106779 433668 106845 433669
rect 106779 433604 106780 433668
rect 106844 433604 106845 433668
rect 106779 433603 106845 433604
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 106411 388380 106477 388381
rect 106411 388316 106412 388380
rect 106476 388316 106477 388380
rect 106411 388315 106477 388316
rect 105123 387020 105189 387021
rect 105123 386956 105124 387020
rect 105188 386956 105189 387020
rect 105123 386955 105189 386956
rect 106043 382396 106109 382397
rect 106043 382332 106044 382396
rect 106108 382332 106109 382396
rect 106043 382331 106109 382332
rect 104203 322148 104269 322149
rect 104203 322084 104204 322148
rect 104268 322084 104269 322148
rect 104203 322083 104269 322084
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 103835 292772 103901 292773
rect 103835 292770 103836 292772
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102731 241772 102797 241773
rect 102731 241708 102732 241772
rect 102796 241708 102797 241772
rect 102731 241707 102797 241708
rect 102731 238100 102797 238101
rect 102731 238036 102732 238100
rect 102796 238036 102797 238100
rect 102731 238035 102797 238036
rect 100891 233884 100957 233885
rect 100891 233820 100892 233884
rect 100956 233820 100957 233884
rect 100891 233819 100957 233820
rect 100707 229804 100773 229805
rect 100707 229740 100708 229804
rect 100772 229740 100773 229804
rect 100707 229739 100773 229740
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 102734 200021 102794 238035
rect 102954 212614 103574 248058
rect 103654 292710 103836 292770
rect 103654 230890 103714 292710
rect 103835 292708 103836 292710
rect 103900 292708 103901 292772
rect 103835 292707 103901 292708
rect 103835 289916 103901 289917
rect 103835 289852 103836 289916
rect 103900 289852 103901 289916
rect 103835 289851 103901 289852
rect 103838 234630 103898 289851
rect 104939 284476 105005 284477
rect 104939 284412 104940 284476
rect 105004 284412 105005 284476
rect 104939 284411 105005 284412
rect 103838 234570 104266 234630
rect 103654 230830 103898 230890
rect 103838 228853 103898 230830
rect 103835 228852 103901 228853
rect 103835 228788 103836 228852
rect 103900 228788 103901 228852
rect 103835 228787 103901 228788
rect 104206 224970 104266 234570
rect 104942 225997 105002 284411
rect 106046 256325 106106 382331
rect 106043 256324 106109 256325
rect 106043 256260 106044 256324
rect 106108 256260 106109 256324
rect 106043 256259 106109 256260
rect 104939 225996 105005 225997
rect 104939 225932 104940 225996
rect 105004 225932 105005 225996
rect 104939 225931 105005 225932
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102731 200020 102797 200021
rect 102731 199956 102732 200020
rect 102796 199956 102797 200020
rect 102731 199955 102797 199956
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 98499 118692 98565 118693
rect 98499 118628 98500 118692
rect 98564 118628 98565 118692
rect 98499 118627 98565 118628
rect 97211 108356 97277 108357
rect 97211 108292 97212 108356
rect 97276 108292 97277 108356
rect 97211 108291 97277 108292
rect 97214 103461 97274 108291
rect 97211 103460 97277 103461
rect 97211 103396 97212 103460
rect 97276 103396 97277 103460
rect 97211 103395 97277 103396
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99051 97204 99117 97205
rect 99051 97140 99052 97204
rect 99116 97140 99117 97204
rect 99051 97139 99117 97140
rect 95187 92444 95253 92445
rect 95187 92380 95188 92444
rect 95252 92380 95253 92444
rect 95187 92379 95253 92380
rect 94083 90812 94149 90813
rect 94083 90748 94084 90812
rect 94148 90748 94149 90812
rect 94083 90747 94149 90748
rect 93899 89588 93965 89589
rect 93899 89524 93900 89588
rect 93964 89524 93965 89588
rect 93899 89523 93965 89524
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 90782
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 99054 3637 99114 97139
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99051 3636 99117 3637
rect 99051 3572 99052 3636
rect 99116 3572 99117 3636
rect 99051 3571 99117 3572
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 176614 103574 212058
rect 103838 224910 104266 224970
rect 103838 202197 103898 224910
rect 106414 220693 106474 388315
rect 106782 385661 106842 433603
rect 107702 391917 107762 449107
rect 109794 436356 110414 470898
rect 111750 441630 111810 583747
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113219 453252 113285 453253
rect 113219 453188 113220 453252
rect 113284 453188 113285 453252
rect 113219 453187 113285 453188
rect 111750 441570 112178 441630
rect 108251 434348 108317 434349
rect 108251 434284 108252 434348
rect 108316 434284 108317 434348
rect 108251 434283 108317 434284
rect 107699 391916 107765 391917
rect 107699 391852 107700 391916
rect 107764 391852 107765 391916
rect 107699 391851 107765 391852
rect 107702 390693 107762 391851
rect 108254 390693 108314 434283
rect 109171 433940 109237 433941
rect 109171 433876 109172 433940
rect 109236 433876 109237 433940
rect 109171 433875 109237 433876
rect 109174 427830 109234 433875
rect 111195 433668 111261 433669
rect 111195 433604 111196 433668
rect 111260 433604 111261 433668
rect 111195 433603 111261 433604
rect 108990 427770 109234 427830
rect 107699 390692 107765 390693
rect 107699 390628 107700 390692
rect 107764 390628 107765 390692
rect 107699 390627 107765 390628
rect 108251 390692 108317 390693
rect 108251 390628 108252 390692
rect 108316 390628 108317 390692
rect 108251 390627 108317 390628
rect 106779 385660 106845 385661
rect 106779 385596 106780 385660
rect 106844 385596 106845 385660
rect 106779 385595 106845 385596
rect 107699 369068 107765 369069
rect 107699 369004 107700 369068
rect 107764 369004 107765 369068
rect 107699 369003 107765 369004
rect 106779 307868 106845 307869
rect 106779 307804 106780 307868
rect 106844 307804 106845 307868
rect 106779 307803 106845 307804
rect 106782 269245 106842 307803
rect 106779 269244 106845 269245
rect 106779 269180 106780 269244
rect 106844 269180 106845 269244
rect 106779 269179 106845 269180
rect 107702 241501 107762 369003
rect 108251 330444 108317 330445
rect 108251 330380 108252 330444
rect 108316 330380 108317 330444
rect 108251 330379 108317 330380
rect 108254 249117 108314 330379
rect 108990 321061 109050 427770
rect 109794 363454 110414 388356
rect 111011 387836 111077 387837
rect 111011 387772 111012 387836
rect 111076 387772 111077 387836
rect 111011 387771 111077 387772
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 108987 321060 109053 321061
rect 108987 320996 108988 321060
rect 109052 320996 109053 321060
rect 108987 320995 109053 320996
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109539 267068 109605 267069
rect 109539 267004 109540 267068
rect 109604 267004 109605 267068
rect 109539 267003 109605 267004
rect 108251 249116 108317 249117
rect 108251 249052 108252 249116
rect 108316 249052 108317 249116
rect 108251 249051 108317 249052
rect 108254 244901 108314 249051
rect 109542 247077 109602 267003
rect 109794 255454 110414 290898
rect 110643 267340 110709 267341
rect 110643 267276 110644 267340
rect 110708 267276 110709 267340
rect 110643 267275 110709 267276
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109539 247076 109605 247077
rect 109539 247012 109540 247076
rect 109604 247012 109605 247076
rect 109539 247011 109605 247012
rect 108251 244900 108317 244901
rect 108251 244836 108252 244900
rect 108316 244836 108317 244900
rect 108251 244835 108317 244836
rect 107699 241500 107765 241501
rect 107699 241436 107700 241500
rect 107764 241436 107765 241500
rect 107699 241435 107765 241436
rect 106779 232796 106845 232797
rect 106779 232732 106780 232796
rect 106844 232732 106845 232796
rect 106779 232731 106845 232732
rect 106411 220692 106477 220693
rect 106411 220628 106412 220692
rect 106476 220628 106477 220692
rect 106411 220627 106477 220628
rect 104019 210356 104085 210357
rect 104019 210292 104020 210356
rect 104084 210292 104085 210356
rect 104019 210291 104085 210292
rect 103835 202196 103901 202197
rect 103835 202132 103836 202196
rect 103900 202132 103901 202196
rect 103835 202131 103901 202132
rect 104022 200130 104082 210291
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 103654 200070 104082 200130
rect 103654 113190 103714 200070
rect 106782 129981 106842 232731
rect 108251 211988 108317 211989
rect 108251 211924 108252 211988
rect 108316 211924 108317 211988
rect 108251 211923 108317 211924
rect 106779 129980 106845 129981
rect 106779 129916 106780 129980
rect 106844 129916 106845 129980
rect 106779 129915 106845 129916
rect 103654 113130 103898 113190
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 103838 89725 103898 113130
rect 108254 98565 108314 211923
rect 109542 200701 109602 247011
rect 109794 219454 110414 254898
rect 110646 224229 110706 267275
rect 111014 246261 111074 387771
rect 111198 381581 111258 433603
rect 112118 432853 112178 441570
rect 112115 432852 112181 432853
rect 112115 432788 112116 432852
rect 112180 432788 112181 432852
rect 112115 432787 112181 432788
rect 112115 426596 112181 426597
rect 112115 426532 112116 426596
rect 112180 426532 112181 426596
rect 112115 426531 112181 426532
rect 112118 412650 112178 426531
rect 112299 420340 112365 420341
rect 112299 420276 112300 420340
rect 112364 420276 112365 420340
rect 112299 420275 112365 420276
rect 111750 412590 112178 412650
rect 111750 387157 111810 412590
rect 111747 387156 111813 387157
rect 111747 387092 111748 387156
rect 111812 387092 111813 387156
rect 111747 387091 111813 387092
rect 111195 381580 111261 381581
rect 111195 381516 111196 381580
rect 111260 381516 111261 381580
rect 111195 381515 111261 381516
rect 112302 271965 112362 420275
rect 113222 396405 113282 453187
rect 113514 439174 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 114507 458828 114573 458829
rect 114507 458764 114508 458828
rect 114572 458764 114573 458828
rect 114507 458763 114573 458764
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 436356 114134 438618
rect 114510 409733 114570 458763
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 114507 409732 114573 409733
rect 114507 409668 114508 409732
rect 114572 409668 114573 409732
rect 114507 409667 114573 409668
rect 115059 408644 115125 408645
rect 115059 408580 115060 408644
rect 115124 408580 115125 408644
rect 115059 408579 115125 408580
rect 113219 396404 113285 396405
rect 113219 396340 113220 396404
rect 113284 396340 113285 396404
rect 113219 396339 113285 396340
rect 113514 367174 114134 388356
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 114507 319564 114573 319565
rect 114507 319500 114508 319564
rect 114572 319500 114573 319564
rect 114507 319499 114573 319500
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 112299 271964 112365 271965
rect 112299 271900 112300 271964
rect 112364 271900 112365 271964
rect 112299 271899 112365 271900
rect 111747 270468 111813 270469
rect 111747 270404 111748 270468
rect 111812 270404 111813 270468
rect 111747 270403 111813 270404
rect 111011 246260 111077 246261
rect 111011 246196 111012 246260
rect 111076 246196 111077 246260
rect 111011 246195 111077 246196
rect 111195 246124 111261 246125
rect 111195 246060 111196 246124
rect 111260 246060 111261 246124
rect 111195 246059 111261 246060
rect 111198 237285 111258 246059
rect 111195 237284 111261 237285
rect 111195 237220 111196 237284
rect 111260 237220 111261 237284
rect 111195 237219 111261 237220
rect 111563 236740 111629 236741
rect 111563 236676 111564 236740
rect 111628 236676 111629 236740
rect 111563 236675 111629 236676
rect 110643 224228 110709 224229
rect 110643 224164 110644 224228
rect 110708 224164 110709 224228
rect 110643 224163 110709 224164
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109539 200700 109605 200701
rect 109539 200636 109540 200700
rect 109604 200636 109605 200700
rect 109539 200635 109605 200636
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 108251 98564 108317 98565
rect 108251 98500 108252 98564
rect 108316 98500 108317 98564
rect 108251 98499 108317 98500
rect 103835 89724 103901 89725
rect 103835 89660 103836 89724
rect 103900 89660 103901 89724
rect 103835 89659 103901 89660
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 111566 3501 111626 236675
rect 111750 231301 111810 270403
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 111747 231300 111813 231301
rect 111747 231236 111748 231300
rect 111812 231236 111813 231300
rect 111747 231235 111813 231236
rect 113514 223174 114134 258618
rect 114510 234565 114570 319499
rect 115062 263669 115122 408579
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 116531 291820 116597 291821
rect 116531 291756 116532 291820
rect 116596 291756 116597 291820
rect 116531 291755 116597 291756
rect 115979 271964 116045 271965
rect 115979 271900 115980 271964
rect 116044 271900 116045 271964
rect 115979 271899 116045 271900
rect 115059 263668 115125 263669
rect 115059 263604 115060 263668
rect 115124 263604 115125 263668
rect 115059 263603 115125 263604
rect 114507 234564 114573 234565
rect 114507 234500 114508 234564
rect 114572 234500 114573 234564
rect 114507 234499 114573 234500
rect 115982 226133 116042 271899
rect 116534 231845 116594 291755
rect 117234 262894 117854 298338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 124259 588028 124325 588029
rect 124259 587964 124260 588028
rect 124324 587964 124325 588028
rect 124259 587963 124325 587964
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 123339 446452 123405 446453
rect 123339 446388 123340 446452
rect 123404 446388 123405 446452
rect 123339 446387 123405 446388
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 123342 396677 123402 446387
rect 123339 396676 123405 396677
rect 123339 396612 123340 396676
rect 123404 396612 123405 396676
rect 123339 396611 123405 396612
rect 124262 389061 124322 587963
rect 127794 561454 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 130331 578372 130397 578373
rect 130331 578308 130332 578372
rect 130396 578308 130397 578372
rect 130331 578307 130397 578308
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 124259 389060 124325 389061
rect 124259 388996 124260 389060
rect 124324 388996 124325 389060
rect 124259 388995 124325 388996
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 118003 282980 118069 282981
rect 118003 282916 118004 282980
rect 118068 282916 118069 282980
rect 118003 282915 118069 282916
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 116531 231844 116597 231845
rect 116531 231780 116532 231844
rect 116596 231780 116597 231844
rect 116531 231779 116597 231780
rect 117234 226894 117854 262338
rect 118006 234429 118066 282915
rect 118739 274684 118805 274685
rect 118739 274620 118740 274684
rect 118804 274620 118805 274684
rect 118739 274619 118805 274620
rect 118742 238101 118802 274619
rect 120954 266614 121574 302058
rect 122603 284340 122669 284341
rect 122603 284276 122604 284340
rect 122668 284276 122669 284340
rect 122603 284275 122669 284276
rect 121683 274684 121749 274685
rect 121683 274620 121684 274684
rect 121748 274620 121749 274684
rect 121683 274619 121749 274620
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 118739 238100 118805 238101
rect 118739 238036 118740 238100
rect 118804 238036 118805 238100
rect 118739 238035 118805 238036
rect 118739 235516 118805 235517
rect 118739 235452 118740 235516
rect 118804 235452 118805 235516
rect 118739 235451 118805 235452
rect 118003 234428 118069 234429
rect 118003 234364 118004 234428
rect 118068 234364 118069 234428
rect 118003 234363 118069 234364
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 115979 226132 116045 226133
rect 115979 226068 115980 226132
rect 116044 226068 116045 226132
rect 115979 226067 116045 226068
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 117083 220148 117149 220149
rect 117083 220084 117084 220148
rect 117148 220084 117149 220148
rect 117083 220083 117149 220084
rect 114507 211852 114573 211853
rect 114507 211788 114508 211852
rect 114572 211788 114573 211852
rect 114507 211787 114573 211788
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 114510 115157 114570 211787
rect 114507 115156 114573 115157
rect 114507 115092 114508 115156
rect 114572 115092 114573 115156
rect 114507 115091 114573 115092
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 111563 3500 111629 3501
rect 111563 3436 111564 3500
rect 111628 3436 111629 3500
rect 111563 3435 111629 3436
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 -2266 114134 6618
rect 117086 3637 117146 220083
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 118742 118965 118802 235451
rect 120954 230614 121574 266058
rect 121686 232797 121746 274619
rect 121683 232796 121749 232797
rect 121683 232732 121684 232796
rect 121748 232732 121749 232796
rect 121683 232731 121749 232732
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 121683 220284 121749 220285
rect 121683 220220 121684 220284
rect 121748 220220 121749 220284
rect 121683 220219 121749 220220
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 118739 118964 118805 118965
rect 118739 118900 118740 118964
rect 118804 118900 118805 118964
rect 118739 118899 118805 118900
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117083 3636 117149 3637
rect 117083 3572 117084 3636
rect 117148 3572 117149 3636
rect 117083 3571 117149 3572
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 122058
rect 121686 100061 121746 220219
rect 122606 148341 122666 284275
rect 124262 244357 124322 388995
rect 127794 381454 128414 416898
rect 128675 389332 128741 389333
rect 128675 389330 128676 389332
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 126835 263668 126901 263669
rect 126835 263604 126836 263668
rect 126900 263604 126901 263668
rect 126835 263603 126901 263604
rect 124443 258092 124509 258093
rect 124443 258028 124444 258092
rect 124508 258028 124509 258092
rect 124443 258027 124509 258028
rect 124259 244356 124325 244357
rect 124259 244292 124260 244356
rect 124324 244292 124325 244356
rect 124259 244291 124325 244292
rect 122603 148340 122669 148341
rect 122603 148276 122604 148340
rect 122668 148276 122669 148340
rect 122603 148275 122669 148276
rect 124446 106317 124506 258027
rect 126838 222053 126898 263603
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 126835 222052 126901 222053
rect 126835 221988 126836 222052
rect 126900 221988 126901 222052
rect 126835 221987 126901 221988
rect 127794 201454 128414 236898
rect 128494 389270 128676 389330
rect 128494 229110 128554 389270
rect 128675 389268 128676 389270
rect 128740 389268 128741 389332
rect 128675 389267 128741 389268
rect 128494 229050 128738 229110
rect 128678 211853 128738 229050
rect 128675 211852 128741 211853
rect 128675 211788 128676 211852
rect 128740 211788 128741 211852
rect 128675 211787 128741 211788
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 124443 106316 124509 106317
rect 124443 106252 124444 106316
rect 124508 106252 124509 106316
rect 124443 106251 124509 106252
rect 121683 100060 121749 100061
rect 121683 99996 121684 100060
rect 121748 99996 121749 100060
rect 121683 99995 121749 99996
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 130334 4997 130394 578307
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 133827 383756 133893 383757
rect 133827 383692 133828 383756
rect 133892 383692 133893 383756
rect 133827 383691 133893 383692
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 133830 215253 133890 383691
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 133827 215252 133893 215253
rect 133827 215188 133828 215252
rect 133892 215188 133893 215252
rect 133827 215187 133893 215188
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 130331 4996 130397 4997
rect 130331 4932 130332 4996
rect 130396 4932 130397 4996
rect 130331 4931 130397 4932
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 186819 303924 186885 303925
rect 186819 303860 186820 303924
rect 186884 303860 186885 303924
rect 186819 303859 186885 303860
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 186822 222869 186882 303859
rect 189234 298894 189854 334338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 191051 320244 191117 320245
rect 191051 320180 191052 320244
rect 191116 320180 191117 320244
rect 191051 320179 191117 320180
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 191054 298757 191114 320179
rect 192707 303652 192773 303653
rect 192707 303588 192708 303652
rect 192772 303588 192773 303652
rect 192954 303592 193574 338058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 303592 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 303592 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 303592 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 303592 211574 320058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 215891 303788 215957 303789
rect 215891 303724 215892 303788
rect 215956 303724 215957 303788
rect 215891 303723 215957 303724
rect 192707 303587 192773 303588
rect 191051 298756 191117 298757
rect 191051 298692 191052 298756
rect 191116 298692 191117 298756
rect 191051 298691 191117 298692
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 192339 247620 192405 247621
rect 192339 247556 192340 247620
rect 192404 247556 192405 247620
rect 192339 247555 192405 247556
rect 191051 244900 191117 244901
rect 191051 244836 191052 244900
rect 191116 244836 191117 244900
rect 191051 244835 191117 244836
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 186819 222868 186885 222869
rect 186819 222804 186820 222868
rect 186884 222804 186885 222868
rect 186819 222803 186885 222804
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 191054 149701 191114 244835
rect 191235 242996 191301 242997
rect 191235 242932 191236 242996
rect 191300 242932 191301 242996
rect 191235 242931 191301 242932
rect 191238 235245 191298 242931
rect 192342 235789 192402 247555
rect 192710 239869 192770 303587
rect 193443 301476 193509 301477
rect 193443 301412 193444 301476
rect 193508 301412 193509 301476
rect 193443 301411 193509 301412
rect 193259 301204 193325 301205
rect 193259 301140 193260 301204
rect 193324 301140 193325 301204
rect 193259 301139 193325 301140
rect 193262 276725 193322 301139
rect 193446 298893 193506 301411
rect 210371 301204 210437 301205
rect 210371 301140 210372 301204
rect 210436 301140 210437 301204
rect 210371 301139 210437 301140
rect 208899 301068 208965 301069
rect 208899 301004 208900 301068
rect 208964 301004 208965 301068
rect 208899 301003 208965 301004
rect 196019 300932 196085 300933
rect 196019 300868 196020 300932
rect 196084 300868 196085 300932
rect 196019 300867 196085 300868
rect 197491 300932 197557 300933
rect 197491 300868 197492 300932
rect 197556 300868 197557 300932
rect 197491 300867 197557 300868
rect 198779 300932 198845 300933
rect 198779 300868 198780 300932
rect 198844 300868 198845 300932
rect 198779 300867 198845 300868
rect 201539 300932 201605 300933
rect 201539 300868 201540 300932
rect 201604 300868 201605 300932
rect 201539 300867 201605 300868
rect 203011 300932 203077 300933
rect 203011 300868 203012 300932
rect 203076 300868 203077 300932
rect 203011 300867 203077 300868
rect 204299 300932 204365 300933
rect 204299 300868 204300 300932
rect 204364 300868 204365 300932
rect 204299 300867 204365 300868
rect 205587 300932 205653 300933
rect 205587 300868 205588 300932
rect 205652 300868 205653 300932
rect 205587 300867 205653 300868
rect 207059 300932 207125 300933
rect 207059 300868 207060 300932
rect 207124 300868 207125 300932
rect 207059 300867 207125 300868
rect 208347 300932 208413 300933
rect 208347 300868 208348 300932
rect 208412 300868 208413 300932
rect 208347 300867 208413 300868
rect 193443 298892 193509 298893
rect 193443 298828 193444 298892
rect 193508 298828 193509 298892
rect 193443 298827 193509 298828
rect 193259 276724 193325 276725
rect 193259 276660 193260 276724
rect 193324 276660 193325 276724
rect 193259 276659 193325 276660
rect 193443 246260 193509 246261
rect 193443 246196 193444 246260
rect 193508 246196 193509 246260
rect 193443 246195 193509 246196
rect 193446 245850 193506 246195
rect 193446 245790 193874 245850
rect 192707 239868 192773 239869
rect 192707 239804 192708 239868
rect 192772 239804 192773 239868
rect 192707 239803 192773 239804
rect 192339 235788 192405 235789
rect 192339 235724 192340 235788
rect 192404 235724 192405 235788
rect 192339 235723 192405 235724
rect 191235 235244 191301 235245
rect 191235 235180 191236 235244
rect 191300 235180 191301 235244
rect 191235 235179 191301 235180
rect 192954 230614 193574 239592
rect 193814 238509 193874 245790
rect 193811 238508 193877 238509
rect 193811 238444 193812 238508
rect 193876 238444 193877 238508
rect 193811 238443 193877 238444
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 191051 149700 191117 149701
rect 191051 149636 191052 149700
rect 191116 149636 191117 149700
rect 191051 149635 191117 149636
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 196022 39269 196082 300867
rect 197494 151061 197554 300867
rect 197776 291454 198096 291486
rect 197776 291218 197818 291454
rect 198054 291218 198096 291454
rect 197776 291134 198096 291218
rect 197776 290898 197818 291134
rect 198054 290898 198096 291134
rect 197776 290866 198096 290898
rect 197776 255454 198096 255486
rect 197776 255218 197818 255454
rect 198054 255218 198096 255454
rect 197776 255134 198096 255218
rect 197776 254898 197818 255134
rect 198054 254898 198096 255134
rect 197776 254866 198096 254898
rect 198782 185605 198842 300867
rect 199794 237454 200414 239592
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 198779 185604 198845 185605
rect 198779 185540 198780 185604
rect 198844 185540 198845 185604
rect 198779 185539 198845 185540
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 197491 151060 197557 151061
rect 197491 150996 197492 151060
rect 197556 150996 197557 151060
rect 197491 150995 197557 150996
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 196019 39268 196085 39269
rect 196019 39204 196020 39268
rect 196084 39204 196085 39268
rect 196019 39203 196085 39204
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 201542 21317 201602 300867
rect 203014 153781 203074 300867
rect 203514 205174 204134 239592
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203011 153780 203077 153781
rect 203011 153716 203012 153780
rect 203076 153716 203077 153780
rect 203011 153715 203077 153716
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 201539 21316 201605 21317
rect 201539 21252 201540 21316
rect 201604 21252 201605 21316
rect 201539 21251 201605 21252
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 24618
rect 204302 22677 204362 300867
rect 205590 200701 205650 300867
rect 207062 240005 207122 300867
rect 207059 240004 207125 240005
rect 207059 239940 207060 240004
rect 207124 239940 207125 240004
rect 207059 239939 207125 239940
rect 207234 208894 207854 239592
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 205587 200700 205653 200701
rect 205587 200636 205588 200700
rect 205652 200636 205653 200700
rect 205587 200635 205653 200636
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 204299 22676 204365 22677
rect 204299 22612 204300 22676
rect 204364 22612 204365 22676
rect 204299 22611 204365 22612
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28338
rect 208350 11661 208410 300867
rect 208902 73813 208962 301003
rect 208899 73812 208965 73813
rect 208899 73748 208900 73812
rect 208964 73748 208965 73812
rect 208899 73747 208965 73748
rect 210374 71093 210434 301139
rect 213683 301068 213749 301069
rect 213683 301004 213684 301068
rect 213748 301004 213749 301068
rect 213683 301003 213749 301004
rect 211659 300932 211725 300933
rect 211659 300868 211660 300932
rect 211724 300868 211725 300932
rect 211659 300867 211725 300868
rect 210954 212614 211574 239592
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210371 71092 210437 71093
rect 210371 71028 210372 71092
rect 210436 71028 210437 71092
rect 210371 71027 210437 71028
rect 210954 68614 211574 104058
rect 211662 76533 211722 300867
rect 213136 273454 213456 273486
rect 213136 273218 213178 273454
rect 213414 273218 213456 273454
rect 213136 273134 213456 273218
rect 213136 272898 213178 273134
rect 213414 272898 213456 273134
rect 213136 272866 213456 272898
rect 213686 186965 213746 301003
rect 213867 300932 213933 300933
rect 213867 300868 213868 300932
rect 213932 300868 213933 300932
rect 213867 300867 213933 300868
rect 214419 300932 214485 300933
rect 214419 300868 214420 300932
rect 214484 300868 214485 300932
rect 214419 300867 214485 300868
rect 213683 186964 213749 186965
rect 213683 186900 213684 186964
rect 213748 186900 213749 186964
rect 213683 186899 213749 186900
rect 211659 76532 211725 76533
rect 211659 76468 211660 76532
rect 211724 76468 211725 76532
rect 211659 76467 211725 76468
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 208347 11660 208413 11661
rect 208347 11596 208348 11660
rect 208412 11596 208413 11660
rect 208347 11595 208413 11596
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 213870 7581 213930 300867
rect 214422 228309 214482 300867
rect 214419 228308 214485 228309
rect 214419 228244 214420 228308
rect 214484 228244 214485 228308
rect 214419 228243 214485 228244
rect 213867 7580 213933 7581
rect 213867 7516 213868 7580
rect 213932 7516 213933 7580
rect 213867 7515 213933 7516
rect 215894 4861 215954 303723
rect 217794 303592 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 218651 305012 218717 305013
rect 218651 304948 218652 305012
rect 218716 304948 218717 305012
rect 218651 304947 218717 304948
rect 216075 300932 216141 300933
rect 216075 300868 216076 300932
rect 216140 300868 216141 300932
rect 216075 300867 216141 300868
rect 216811 300932 216877 300933
rect 216811 300868 216812 300932
rect 216876 300868 216877 300932
rect 216811 300867 216877 300868
rect 216078 224229 216138 300867
rect 216814 225589 216874 300867
rect 216811 225588 216877 225589
rect 216811 225524 216812 225588
rect 216876 225524 216877 225588
rect 216811 225523 216877 225524
rect 216075 224228 216141 224229
rect 216075 224164 216076 224228
rect 216140 224164 216141 224228
rect 216075 224163 216141 224164
rect 217794 219454 218414 239592
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 218654 202877 218714 304947
rect 221514 303592 222134 330618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 303592 225854 334338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 303592 229574 338058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 303592 236414 308898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 237787 303652 237853 303653
rect 237787 303588 237788 303652
rect 237852 303588 237853 303652
rect 239514 303592 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 242019 303924 242085 303925
rect 242019 303860 242020 303924
rect 242084 303860 242085 303924
rect 242019 303859 242085 303860
rect 237787 303587 237853 303588
rect 222699 301204 222765 301205
rect 222699 301140 222700 301204
rect 222764 301140 222765 301204
rect 222699 301139 222765 301140
rect 219387 301068 219453 301069
rect 219387 301004 219388 301068
rect 219452 301004 219453 301068
rect 219387 301003 219453 301004
rect 221227 301068 221293 301069
rect 221227 301004 221228 301068
rect 221292 301004 221293 301068
rect 221227 301003 221293 301004
rect 219390 300930 219450 301003
rect 219206 300870 219450 300930
rect 219571 300932 219637 300933
rect 218651 202876 218717 202877
rect 218651 202812 218652 202876
rect 218716 202812 218717 202876
rect 218651 202811 218717 202812
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 215891 4860 215957 4861
rect 215891 4796 215892 4860
rect 215956 4796 215957 4860
rect 215891 4795 215957 4796
rect 217794 3454 218414 38898
rect 219206 33829 219266 300870
rect 219571 300868 219572 300932
rect 219636 300868 219637 300932
rect 219571 300867 219637 300868
rect 220859 300932 220925 300933
rect 220859 300868 220860 300932
rect 220924 300868 220925 300932
rect 220859 300867 220925 300868
rect 219574 188325 219634 300867
rect 220862 240141 220922 300867
rect 220859 240140 220925 240141
rect 220859 240076 220860 240140
rect 220924 240076 220925 240140
rect 220859 240075 220925 240076
rect 221230 214573 221290 301003
rect 222331 300932 222397 300933
rect 222331 300868 222332 300932
rect 222396 300868 222397 300932
rect 222331 300867 222397 300868
rect 221514 223174 222134 239592
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221227 214572 221293 214573
rect 221227 214508 221228 214572
rect 221292 214508 221293 214572
rect 221227 214507 221293 214508
rect 219571 188324 219637 188325
rect 219571 188260 219572 188324
rect 219636 188260 219637 188324
rect 219571 188259 219637 188260
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 219203 33828 219269 33829
rect 219203 33764 219204 33828
rect 219268 33764 219269 33828
rect 219203 33763 219269 33764
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 42618
rect 222334 35189 222394 300867
rect 222331 35188 222397 35189
rect 222331 35124 222332 35188
rect 222396 35124 222397 35188
rect 222331 35123 222397 35124
rect 222702 24173 222762 301139
rect 223803 301068 223869 301069
rect 223803 301004 223804 301068
rect 223868 301004 223869 301068
rect 223803 301003 223869 301004
rect 230427 301068 230493 301069
rect 230427 301004 230428 301068
rect 230492 301004 230493 301068
rect 230427 301003 230493 301004
rect 232083 301068 232149 301069
rect 232083 301004 232084 301068
rect 232148 301004 232149 301068
rect 232083 301003 232149 301004
rect 233187 301068 233253 301069
rect 233187 301004 233188 301068
rect 233252 301004 233253 301068
rect 233187 301003 233253 301004
rect 234843 301068 234909 301069
rect 234843 301004 234844 301068
rect 234908 301004 234909 301068
rect 234843 301003 234909 301004
rect 223806 146981 223866 301003
rect 223987 300932 224053 300933
rect 223987 300868 223988 300932
rect 224052 300868 224053 300932
rect 223987 300867 224053 300868
rect 225091 300932 225157 300933
rect 225091 300868 225092 300932
rect 225156 300868 225157 300932
rect 225091 300867 225157 300868
rect 226379 300932 226445 300933
rect 226379 300868 226380 300932
rect 226444 300868 226445 300932
rect 226379 300867 226445 300868
rect 226563 300932 226629 300933
rect 226563 300868 226564 300932
rect 226628 300868 226629 300932
rect 226563 300867 226629 300868
rect 227667 300932 227733 300933
rect 227667 300868 227668 300932
rect 227732 300868 227733 300932
rect 227667 300867 227733 300868
rect 229691 300932 229757 300933
rect 229691 300868 229692 300932
rect 229756 300868 229757 300932
rect 229691 300867 229757 300868
rect 223803 146980 223869 146981
rect 223803 146916 223804 146980
rect 223868 146916 223869 146980
rect 223803 146915 223869 146916
rect 223990 36549 224050 300867
rect 225094 93870 225154 300867
rect 224910 93810 225154 93870
rect 225234 226894 225854 239592
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 224910 89045 224970 93810
rect 224907 89044 224973 89045
rect 224907 88980 224908 89044
rect 224972 88980 224973 89044
rect 224907 88979 224973 88980
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 223987 36548 224053 36549
rect 223987 36484 223988 36548
rect 224052 36484 224053 36548
rect 223987 36483 224053 36484
rect 222699 24172 222765 24173
rect 222699 24108 222700 24172
rect 222764 24108 222765 24172
rect 222699 24107 222765 24108
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 46338
rect 226382 25533 226442 300867
rect 226566 47565 226626 300867
rect 226563 47564 226629 47565
rect 226563 47500 226564 47564
rect 226628 47500 226629 47564
rect 226563 47499 226629 47500
rect 227670 28253 227730 300867
rect 228496 291454 228816 291486
rect 228496 291218 228538 291454
rect 228774 291218 228816 291454
rect 228496 291134 228816 291218
rect 228496 290898 228538 291134
rect 228774 290898 228816 291134
rect 228496 290866 228816 290898
rect 228496 255454 228816 255486
rect 228496 255218 228538 255454
rect 228774 255218 228816 255454
rect 228496 255134 228816 255218
rect 228496 254898 228538 255134
rect 228774 254898 228816 255134
rect 228496 254866 228816 254898
rect 228954 230614 229574 239592
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 229694 72453 229754 300867
rect 229691 72452 229757 72453
rect 229691 72388 229692 72452
rect 229756 72388 229757 72452
rect 229691 72387 229757 72388
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 227667 28252 227733 28253
rect 227667 28188 227668 28252
rect 227732 28188 227733 28252
rect 227667 28187 227733 28188
rect 226379 25532 226445 25533
rect 226379 25468 226380 25532
rect 226444 25468 226445 25532
rect 226379 25467 226445 25468
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 50058
rect 230430 30973 230490 301003
rect 230979 300932 231045 300933
rect 230979 300868 230980 300932
rect 231044 300868 231045 300932
rect 230979 300867 231045 300868
rect 230982 200701 231042 300867
rect 230979 200700 231045 200701
rect 230979 200636 230980 200700
rect 231044 200636 231045 200700
rect 230979 200635 231045 200636
rect 232086 97205 232146 301003
rect 232267 300932 232333 300933
rect 232267 300868 232268 300932
rect 232332 300868 232333 300932
rect 232267 300867 232333 300868
rect 232083 97204 232149 97205
rect 232083 97140 232084 97204
rect 232148 97140 232149 97204
rect 232083 97139 232149 97140
rect 232270 94485 232330 300867
rect 232267 94484 232333 94485
rect 232267 94420 232268 94484
rect 232332 94420 232333 94484
rect 232267 94419 232333 94420
rect 230427 30972 230493 30973
rect 230427 30908 230428 30972
rect 230492 30908 230493 30972
rect 230427 30907 230493 30908
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 233190 8941 233250 301003
rect 233371 300932 233437 300933
rect 233371 300868 233372 300932
rect 233436 300868 233437 300932
rect 233371 300867 233437 300868
rect 234659 300932 234725 300933
rect 234659 300868 234660 300932
rect 234724 300868 234725 300932
rect 234659 300867 234725 300868
rect 233374 104141 233434 300867
rect 234662 240141 234722 300867
rect 234659 240140 234725 240141
rect 234659 240076 234660 240140
rect 234724 240076 234725 240140
rect 234659 240075 234725 240076
rect 234846 220149 234906 301003
rect 236499 300932 236565 300933
rect 236499 300868 236500 300932
rect 236564 300868 236565 300932
rect 236499 300867 236565 300868
rect 235794 237454 236414 239592
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 234843 220148 234909 220149
rect 234843 220084 234844 220148
rect 234908 220084 234909 220148
rect 234843 220083 234909 220084
rect 235794 201454 236414 236898
rect 236502 215933 236562 300867
rect 236499 215932 236565 215933
rect 236499 215868 236500 215932
rect 236564 215868 236565 215932
rect 236499 215867 236565 215868
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 233371 104140 233437 104141
rect 233371 104076 233372 104140
rect 233436 104076 233437 104140
rect 233371 104075 233437 104076
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 237790 29613 237850 303587
rect 240363 302292 240429 302293
rect 240363 302228 240364 302292
rect 240428 302228 240429 302292
rect 240363 302227 240429 302228
rect 238155 300932 238221 300933
rect 238155 300868 238156 300932
rect 238220 300868 238221 300932
rect 238707 300932 238773 300933
rect 238707 300930 238708 300932
rect 238155 300867 238221 300868
rect 238526 300870 238708 300930
rect 238158 239050 238218 300867
rect 238526 296730 238586 300870
rect 238707 300868 238708 300870
rect 238772 300868 238773 300932
rect 238707 300867 238773 300868
rect 238526 296670 238954 296730
rect 238894 295490 238954 296670
rect 238526 295430 238954 295490
rect 238526 288010 238586 295430
rect 238526 287950 238954 288010
rect 238894 287070 238954 287950
rect 238526 287010 238954 287070
rect 238526 277410 238586 287010
rect 238526 277350 238954 277410
rect 238894 276450 238954 277350
rect 238526 276390 238954 276450
rect 238526 268970 238586 276390
rect 238526 268910 238954 268970
rect 238894 267750 238954 268910
rect 238526 267690 238954 267750
rect 238526 258090 238586 267690
rect 238526 258030 238954 258090
rect 238894 256730 238954 258030
rect 238526 256670 238954 256730
rect 238526 249250 238586 256670
rect 238526 249190 238954 249250
rect 238894 248430 238954 249190
rect 238526 248370 238954 248430
rect 238526 239730 238586 248370
rect 238526 239670 238954 239730
rect 238158 238990 238586 239050
rect 238526 101421 238586 238990
rect 238894 238373 238954 239670
rect 238891 238372 238957 238373
rect 238891 238308 238892 238372
rect 238956 238308 238957 238372
rect 238891 238307 238957 238308
rect 238707 229124 238773 229125
rect 238707 229060 238708 229124
rect 238772 229060 238773 229124
rect 238707 229059 238773 229060
rect 238710 228853 238770 229059
rect 238707 228852 238773 228853
rect 238707 228788 238708 228852
rect 238772 228788 238773 228852
rect 238707 228787 238773 228788
rect 238891 219468 238957 219469
rect 238891 219404 238892 219468
rect 238956 219404 238957 219468
rect 238891 219403 238957 219404
rect 238894 219061 238954 219403
rect 238891 219060 238957 219061
rect 238891 218996 238892 219060
rect 238956 218996 238957 219060
rect 238891 218995 238957 218996
rect 238707 209812 238773 209813
rect 238707 209748 238708 209812
rect 238772 209790 238773 209812
rect 238772 209748 238954 209790
rect 238707 209747 238954 209748
rect 238710 209730 238954 209747
rect 238894 209541 238954 209730
rect 238891 209540 238957 209541
rect 238891 209476 238892 209540
rect 238956 209476 238957 209540
rect 238891 209475 238957 209476
rect 239514 205174 240134 239592
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 238891 200156 238957 200157
rect 238891 200092 238892 200156
rect 238956 200092 238957 200156
rect 238891 200091 238957 200092
rect 238894 199885 238954 200091
rect 238891 199884 238957 199885
rect 238891 199820 238892 199884
rect 238956 199820 238957 199884
rect 238891 199819 238957 199820
rect 238707 190500 238773 190501
rect 238707 190436 238708 190500
rect 238772 190436 238773 190500
rect 238707 190435 238773 190436
rect 238710 190229 238770 190435
rect 238707 190228 238773 190229
rect 238707 190164 238708 190228
rect 238772 190164 238773 190228
rect 238707 190163 238773 190164
rect 238707 180844 238773 180845
rect 238707 180780 238708 180844
rect 238772 180780 238773 180844
rect 238707 180779 238773 180780
rect 238710 180573 238770 180779
rect 238707 180572 238773 180573
rect 238707 180508 238708 180572
rect 238772 180508 238773 180572
rect 238707 180507 238773 180508
rect 238707 171188 238773 171189
rect 238707 171124 238708 171188
rect 238772 171124 238773 171188
rect 238707 171123 238773 171124
rect 238710 171053 238770 171123
rect 238707 171052 238773 171053
rect 238707 170988 238708 171052
rect 238772 170988 238773 171052
rect 238707 170987 238773 170988
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238891 161532 238957 161533
rect 238891 161490 238892 161532
rect 238710 161468 238892 161490
rect 238956 161468 238957 161532
rect 238710 161467 238957 161468
rect 238710 161430 238954 161467
rect 238710 161261 238770 161430
rect 238707 161260 238773 161261
rect 238707 161196 238708 161260
rect 238772 161196 238773 161260
rect 238707 161195 238773 161196
rect 238707 151876 238773 151877
rect 238707 151812 238708 151876
rect 238772 151812 238773 151876
rect 238707 151811 238773 151812
rect 238710 151605 238770 151811
rect 238707 151604 238773 151605
rect 238707 151540 238708 151604
rect 238772 151540 238773 151604
rect 238707 151539 238773 151540
rect 239259 145620 239325 145621
rect 239259 145556 239260 145620
rect 239324 145556 239325 145620
rect 239259 145555 239325 145556
rect 239262 138685 239322 145555
rect 239259 138684 239325 138685
rect 239259 138620 239260 138684
rect 239324 138620 239325 138684
rect 239259 138619 239325 138620
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 238523 101420 238589 101421
rect 238523 101356 238524 101420
rect 238588 101356 238589 101420
rect 238523 101355 238589 101356
rect 237787 29612 237853 29613
rect 237787 29548 237788 29612
rect 237852 29548 237853 29612
rect 237787 29547 237853 29548
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 233187 8940 233253 8941
rect 233187 8876 233188 8940
rect 233252 8876 233253 8940
rect 233187 8875 233253 8876
rect 235794 -1306 236414 20898
rect 238526 4045 238586 101355
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 238523 4044 238589 4045
rect 238523 3980 238524 4044
rect 238588 3980 238589 4044
rect 238523 3979 238589 3980
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 24618
rect 240366 3501 240426 302227
rect 242022 237421 242082 303859
rect 243234 303592 243854 316338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 255451 330444 255517 330445
rect 255451 330380 255452 330444
rect 255516 330380 255517 330444
rect 255451 330379 255517 330380
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 252507 325004 252573 325005
rect 252507 324940 252508 325004
rect 252572 324940 252573 325004
rect 252507 324939 252573 324940
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 303592 247574 320058
rect 244411 300932 244477 300933
rect 244411 300868 244412 300932
rect 244476 300868 244477 300932
rect 244411 300867 244477 300868
rect 243856 273454 244176 273486
rect 243856 273218 243898 273454
rect 244134 273218 244176 273454
rect 243856 273134 244176 273218
rect 243856 272898 243898 273134
rect 244134 272898 244176 273134
rect 243856 272866 244176 272898
rect 242019 237420 242085 237421
rect 242019 237356 242020 237420
rect 242084 237356 242085 237420
rect 242019 237355 242085 237356
rect 243234 208894 243854 239592
rect 244414 217293 244474 300867
rect 252510 296730 252570 324939
rect 252691 316300 252757 316301
rect 252691 316236 252692 316300
rect 252756 316236 252757 316300
rect 252691 316235 252757 316236
rect 252694 306390 252754 316235
rect 252694 306330 252938 306390
rect 252878 297941 252938 306330
rect 253794 303592 254414 326898
rect 254531 315348 254597 315349
rect 254531 315284 254532 315348
rect 254596 315284 254597 315348
rect 254531 315283 254597 315284
rect 254163 301612 254229 301613
rect 254163 301548 254164 301612
rect 254228 301548 254229 301612
rect 254163 301547 254229 301548
rect 252875 297940 252941 297941
rect 252875 297876 252876 297940
rect 252940 297876 252941 297940
rect 252875 297875 252941 297876
rect 252510 296670 252938 296730
rect 252878 291413 252938 296670
rect 252875 291412 252941 291413
rect 252875 291348 252876 291412
rect 252940 291348 252941 291412
rect 252875 291347 252941 291348
rect 253979 265980 254045 265981
rect 253979 265916 253980 265980
rect 254044 265916 254045 265980
rect 253979 265915 254045 265916
rect 252875 261764 252941 261765
rect 252875 261700 252876 261764
rect 252940 261700 252941 261764
rect 252875 261699 252941 261700
rect 252878 258090 252938 261699
rect 252510 258030 252938 258090
rect 252510 239597 252570 258030
rect 253611 244764 253677 244765
rect 253611 244700 253612 244764
rect 253676 244700 253677 244764
rect 253611 244699 253677 244700
rect 253614 241229 253674 244699
rect 253982 241501 254042 265915
rect 254166 265029 254226 301547
rect 254534 300253 254594 315283
rect 254531 300252 254597 300253
rect 254531 300188 254532 300252
rect 254596 300188 254597 300252
rect 254531 300187 254597 300188
rect 255454 299845 255514 330379
rect 255451 299844 255517 299845
rect 255451 299780 255452 299844
rect 255516 299780 255517 299844
rect 255451 299779 255517 299780
rect 255267 298484 255333 298485
rect 255267 298420 255268 298484
rect 255332 298420 255333 298484
rect 255267 298419 255333 298420
rect 255270 294541 255330 298419
rect 257514 295174 258134 330618
rect 261234 694894 261854 708122
rect 263363 702676 263429 702677
rect 263363 702612 263364 702676
rect 263428 702612 263429 702676
rect 263363 702611 263429 702612
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 258395 318068 258461 318069
rect 258395 318004 258396 318068
rect 258460 318004 258461 318068
rect 258395 318003 258461 318004
rect 258398 296730 258458 318003
rect 260235 303788 260301 303789
rect 260235 303724 260236 303788
rect 260300 303724 260301 303788
rect 260235 303723 260301 303724
rect 260051 303652 260117 303653
rect 260051 303588 260052 303652
rect 260116 303588 260117 303652
rect 260051 303587 260117 303588
rect 258579 301204 258645 301205
rect 258579 301140 258580 301204
rect 258644 301140 258645 301204
rect 258579 301139 258645 301140
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 255267 294540 255333 294541
rect 255267 294476 255268 294540
rect 255332 294476 255333 294540
rect 255267 294475 255333 294476
rect 255451 294404 255517 294405
rect 255451 294340 255452 294404
rect 255516 294340 255517 294404
rect 255451 294339 255517 294340
rect 255454 293181 255514 294339
rect 255819 293860 255885 293861
rect 255819 293796 255820 293860
rect 255884 293796 255885 293860
rect 255819 293795 255885 293796
rect 255451 293180 255517 293181
rect 255451 293116 255452 293180
rect 255516 293116 255517 293180
rect 255451 293115 255517 293116
rect 255822 279445 255882 293795
rect 255819 279444 255885 279445
rect 255819 279380 255820 279444
rect 255884 279380 255885 279444
rect 255819 279379 255885 279380
rect 255819 271148 255885 271149
rect 255819 271084 255820 271148
rect 255884 271084 255885 271148
rect 255819 271083 255885 271084
rect 254163 265028 254229 265029
rect 254163 264964 254164 265028
rect 254228 264964 254229 265028
rect 254163 264963 254229 264964
rect 255822 261901 255882 271083
rect 256739 262308 256805 262309
rect 256739 262244 256740 262308
rect 256804 262244 256805 262308
rect 256739 262243 256805 262244
rect 255819 261900 255885 261901
rect 255819 261836 255820 261900
rect 255884 261836 255885 261900
rect 255819 261835 255885 261836
rect 255267 259996 255333 259997
rect 255267 259932 255268 259996
rect 255332 259932 255333 259996
rect 255267 259931 255333 259932
rect 254531 258228 254597 258229
rect 254531 258164 254532 258228
rect 254596 258164 254597 258228
rect 254531 258163 254597 258164
rect 253979 241500 254045 241501
rect 253979 241436 253980 241500
rect 254044 241436 254045 241500
rect 253979 241435 254045 241436
rect 253611 241228 253677 241229
rect 253611 241164 253612 241228
rect 253676 241164 253677 241228
rect 253611 241163 253677 241164
rect 253611 240820 253677 240821
rect 253611 240756 253612 240820
rect 253676 240756 253677 240820
rect 253611 240755 253677 240756
rect 252507 239596 252573 239597
rect 244411 217292 244477 217293
rect 244411 217228 244412 217292
rect 244476 217228 244477 217292
rect 244411 217227 244477 217228
rect 244414 216749 244474 217227
rect 244411 216748 244477 216749
rect 244411 216684 244412 216748
rect 244476 216684 244477 216748
rect 244411 216683 244477 216684
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 240363 3500 240429 3501
rect 240363 3436 240364 3500
rect 240428 3436 240429 3500
rect 240363 3435 240429 3436
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 212614 247574 239592
rect 252507 239532 252508 239596
rect 252572 239532 252573 239596
rect 252507 239531 252573 239532
rect 253614 237285 253674 240755
rect 253611 237284 253677 237285
rect 253611 237220 253612 237284
rect 253676 237220 253677 237284
rect 253611 237219 253677 237220
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 219454 254414 239592
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 254534 200021 254594 258163
rect 255270 244765 255330 259931
rect 255267 244764 255333 244765
rect 255267 244700 255268 244764
rect 255332 244700 255333 244764
rect 255267 244699 255333 244700
rect 255267 244492 255333 244493
rect 255267 244428 255268 244492
rect 255332 244428 255333 244492
rect 255267 244427 255333 244428
rect 255270 237965 255330 244427
rect 255819 243132 255885 243133
rect 255819 243068 255820 243132
rect 255884 243068 255885 243132
rect 255819 243067 255885 243068
rect 255267 237964 255333 237965
rect 255267 237900 255268 237964
rect 255332 237900 255333 237964
rect 255267 237899 255333 237900
rect 255270 237421 255330 237899
rect 255267 237420 255333 237421
rect 255267 237356 255268 237420
rect 255332 237356 255333 237420
rect 255267 237355 255333 237356
rect 255822 234701 255882 243067
rect 255819 234700 255885 234701
rect 255819 234636 255820 234700
rect 255884 234636 255885 234700
rect 255819 234635 255885 234636
rect 255822 209677 255882 234635
rect 256742 233205 256802 262243
rect 257514 259174 258134 294618
rect 258214 296670 258458 296730
rect 258214 267750 258274 296670
rect 258582 289101 258642 301139
rect 258579 289100 258645 289101
rect 258579 289036 258580 289100
rect 258644 289036 258645 289100
rect 258579 289035 258645 289036
rect 260054 283525 260114 303587
rect 260238 284885 260298 303723
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 260235 284884 260301 284885
rect 260235 284820 260236 284884
rect 260300 284820 260301 284884
rect 260235 284819 260301 284820
rect 260051 283524 260117 283525
rect 260051 283460 260052 283524
rect 260116 283460 260117 283524
rect 260051 283459 260117 283460
rect 258214 267690 258458 267750
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 256739 233204 256805 233205
rect 256739 233140 256740 233204
rect 256804 233140 256805 233204
rect 256739 233139 256805 233140
rect 257514 223174 258134 258618
rect 258398 256869 258458 267690
rect 261234 262894 261854 298338
rect 263366 266525 263426 702611
rect 264099 702540 264165 702541
rect 264099 702476 264100 702540
rect 264164 702476 264165 702540
rect 264099 702475 264165 702476
rect 264102 310861 264162 702475
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264099 310860 264165 310861
rect 264099 310796 264100 310860
rect 264164 310796 264165 310860
rect 264099 310795 264165 310796
rect 264102 296730 264162 310795
rect 263550 296670 264162 296730
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 263363 266524 263429 266525
rect 263363 266460 263364 266524
rect 263428 266460 263429 266524
rect 263363 266459 263429 266460
rect 263550 263125 263610 296670
rect 264954 266614 265574 302058
rect 263731 266524 263797 266525
rect 263731 266460 263732 266524
rect 263796 266460 263797 266524
rect 263731 266459 263797 266460
rect 263547 263124 263613 263125
rect 263547 263060 263548 263124
rect 263612 263060 263613 263124
rect 263547 263059 263613 263060
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 259683 260948 259749 260949
rect 259683 260884 259684 260948
rect 259748 260884 259749 260948
rect 259683 260883 259749 260884
rect 258395 256868 258461 256869
rect 258395 256804 258396 256868
rect 258460 256804 258461 256868
rect 258395 256803 258461 256804
rect 258395 256052 258461 256053
rect 258395 256050 258396 256052
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 255819 209676 255885 209677
rect 255819 209612 255820 209676
rect 255884 209612 255885 209676
rect 255819 209611 255885 209612
rect 254531 200020 254597 200021
rect 254531 199956 254532 200020
rect 254596 199956 254597 200020
rect 254531 199955 254597 199956
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 187174 258134 222618
rect 258214 255990 258396 256050
rect 258214 222050 258274 255990
rect 258395 255988 258396 255990
rect 258460 255988 258461 256052
rect 258395 255987 258461 255988
rect 258395 255372 258461 255373
rect 258395 255308 258396 255372
rect 258460 255308 258461 255372
rect 258395 255307 258461 255308
rect 258398 231845 258458 255307
rect 259499 244356 259565 244357
rect 259499 244292 259500 244356
rect 259564 244292 259565 244356
rect 259499 244291 259565 244292
rect 258395 231844 258461 231845
rect 258395 231780 258396 231844
rect 258460 231780 258461 231844
rect 258395 231779 258461 231780
rect 258395 222052 258461 222053
rect 258395 222050 258396 222052
rect 258214 221990 258396 222050
rect 258395 221988 258396 221990
rect 258460 221988 258461 222052
rect 258395 221987 258461 221988
rect 259502 206821 259562 244291
rect 259686 226949 259746 260883
rect 259683 226948 259749 226949
rect 259683 226884 259684 226948
rect 259748 226884 259749 226948
rect 259683 226883 259749 226884
rect 261234 226894 261854 262338
rect 262259 256732 262325 256733
rect 262259 256668 262260 256732
rect 262324 256668 262325 256732
rect 262259 256667 262325 256668
rect 262262 234565 262322 256667
rect 262259 234564 262325 234565
rect 262259 234500 262260 234564
rect 262324 234500 262325 234564
rect 262259 234499 262325 234500
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 259499 206820 259565 206821
rect 259499 206756 259500 206820
rect 259564 206756 259565 206820
rect 259499 206755 259565 206756
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 190894 261854 226338
rect 263734 220693 263794 266459
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 263731 220692 263797 220693
rect 263731 220628 263732 220692
rect 263796 220628 263797 220692
rect 263731 220627 263797 220628
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 73721 543218 73957 543454
rect 73721 542898 73957 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 77686 561218 77922 561454
rect 77686 560898 77922 561134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81651 543218 81887 543454
rect 81651 542898 81887 543134
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 85617 561218 85853 561454
rect 85617 560898 85853 561134
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 89582 543218 89818 543454
rect 89582 542898 89818 543134
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 79019 273218 79255 273454
rect 79019 272898 79255 273134
rect 88283 273218 88519 273454
rect 88283 272898 88519 273134
rect 74387 255218 74623 255454
rect 74387 254898 74623 255134
rect 83651 255218 83887 255454
rect 83651 254898 83887 255134
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 92915 255218 93151 255454
rect 92915 254898 93151 255134
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 77686 129218 77922 129454
rect 77686 128898 77922 129134
rect 85617 129218 85853 129454
rect 85617 128898 85853 129134
rect 73721 111218 73957 111454
rect 73721 110898 73957 111134
rect 81651 111218 81887 111454
rect 81651 110898 81887 111134
rect 89582 111218 89818 111454
rect 89582 110898 89818 111134
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 197818 291218 198054 291454
rect 197818 290898 198054 291134
rect 197818 255218 198054 255454
rect 197818 254898 198054 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 213178 273218 213414 273454
rect 213178 272898 213414 273134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 228538 291218 228774 291454
rect 228538 290898 228774 291134
rect 228538 255218 228774 255454
rect 228538 254898 228774 255134
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 243898 273218 244134 273454
rect 243898 272898 244134 273134
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 77686 561454
rect 77922 561218 85617 561454
rect 85853 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 77686 561134
rect 77922 560898 85617 561134
rect 85853 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73721 543454
rect 73957 543218 81651 543454
rect 81887 543218 89582 543454
rect 89818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73721 543134
rect 73957 542898 81651 543134
rect 81887 542898 89582 543134
rect 89818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 197818 291454
rect 198054 291218 228538 291454
rect 228774 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 197818 291134
rect 198054 290898 228538 291134
rect 228774 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 79019 273454
rect 79255 273218 88283 273454
rect 88519 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 213178 273454
rect 213414 273218 243898 273454
rect 244134 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 79019 273134
rect 79255 272898 88283 273134
rect 88519 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 213178 273134
rect 213414 272898 243898 273134
rect 244134 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74387 255454
rect 74623 255218 83651 255454
rect 83887 255218 92915 255454
rect 93151 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 197818 255454
rect 198054 255218 228538 255454
rect 228774 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74387 255134
rect 74623 254898 83651 255134
rect 83887 254898 92915 255134
rect 93151 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 197818 255134
rect 198054 254898 228538 255134
rect 228774 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 77686 129454
rect 77922 129218 85617 129454
rect 85853 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 77686 129134
rect 77922 128898 85617 129134
rect 85853 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73721 111454
rect 73957 111218 81651 111454
rect 81887 111218 89582 111454
rect 89818 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73721 111134
rect 73957 110898 81651 111134
rect 81887 110898 89582 111134
rect 89818 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use zube_wrapped_project  zube_wrapped_project_5
timestamp 1635173914
transform 1 0 193568 0 1 241592
box 0 0 60000 60000
use wrapped_vga_clock  wrapped_vga_clock_2
timestamp 1635173914
transform 1 0 68770 0 1 390356
box 0 0 44000 44000
use wrapped_tpm2137  wrapped_tpm2137_3
timestamp 1635173914
transform 1 0 68770 0 1 539166
box 0 0 26000 42000
use wrapped_rgb_mixer  wrapped_rgb_mixer_0
timestamp 1635173914
transform 1 0 68770 0 1 92782
box 0 0 26000 42000
use wrapped_frequency_counter  wrapped_frequency_counter_1
timestamp 1635173914
transform 1 0 68770 0 1 241592
box 0 0 30000 42000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 90782 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 136782 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 436356 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 583166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 436356 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 303592 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 303592 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 90782 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 136782 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 436356 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 583166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 436356 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 303592 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 90782 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 136782 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 436356 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 583166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 303592 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 90782 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 136782 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 436356 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 583166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 303592 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 303592 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 436356 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 303592 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 303592 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 90782 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 136782 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 436356 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 583166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 436356 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 303592 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 303592 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 90782 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 136782 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 436356 92414 537166 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 583166 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 303592 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 303592 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 90782 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 136782 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 436356 96134 537166 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 583166 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 303592 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 303592 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
